module real_jpeg_17449_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_572;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_0),
.A2(n_80),
.B1(n_84),
.B2(n_87),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_0),
.A2(n_87),
.B1(n_196),
.B2(n_202),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_0),
.A2(n_87),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_1),
.A2(n_41),
.B1(n_177),
.B2(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_3),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_3),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_3),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_4),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_4),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_4),
.A2(n_166),
.B1(n_214),
.B2(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_4),
.A2(n_214),
.B1(n_409),
.B2(n_412),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_4),
.A2(n_214),
.B1(n_504),
.B2(n_507),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_5),
.A2(n_119),
.B1(n_123),
.B2(n_125),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_5),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_5),
.A2(n_125),
.B1(n_220),
.B2(n_223),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_5),
.A2(n_125),
.B1(n_312),
.B2(n_317),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_5),
.A2(n_125),
.B1(n_373),
.B2(n_375),
.Y(n_372)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_6),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_7),
.Y(n_151)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_7),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_7),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_8),
.A2(n_68),
.B1(n_72),
.B2(n_77),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_8),
.A2(n_77),
.B1(n_165),
.B2(n_170),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_8),
.A2(n_77),
.B1(n_289),
.B2(n_292),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_9),
.B(n_279),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_9),
.A2(n_278),
.B(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_9),
.Y(n_378)
);

OAI32xp33_ASAP7_75t_L g419 ( 
.A1(n_9),
.A2(n_411),
.A3(n_420),
.B1(n_424),
.B2(n_426),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_9),
.A2(n_378),
.B1(n_466),
.B2(n_470),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_9),
.B(n_161),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_9),
.A2(n_26),
.B1(n_543),
.B2(n_551),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_10),
.A2(n_116),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_10),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_10),
.A2(n_302),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_10),
.A2(n_302),
.B1(n_454),
.B2(n_457),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_SL g518 ( 
.A1(n_10),
.A2(n_302),
.B1(n_519),
.B2(n_522),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_11),
.A2(n_297),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_11),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_11),
.A2(n_300),
.B1(n_364),
.B2(n_368),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_11),
.A2(n_80),
.B1(n_300),
.B2(n_499),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_11),
.A2(n_300),
.B1(n_544),
.B2(n_547),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_12),
.A2(n_155),
.B1(n_158),
.B2(n_160),
.Y(n_154)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_12),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_12),
.A2(n_80),
.B1(n_160),
.B2(n_188),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_12),
.A2(n_116),
.B1(n_160),
.B2(n_234),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_12),
.A2(n_160),
.B1(n_284),
.B2(n_287),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_13),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_13),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_13),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_14),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_14),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_15),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_15),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_15),
.A2(n_114),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_15),
.A2(n_114),
.B1(n_350),
.B2(n_352),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_15),
.A2(n_114),
.B1(n_430),
.B2(n_434),
.Y(n_429)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_16),
.Y(n_201)
);

BUFx4f_ASAP7_75t_L g205 ( 
.A(n_16),
.Y(n_205)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_17),
.Y(n_113)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_17),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g280 ( 
.A(n_17),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_249),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_248),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_227),
.Y(n_20)
);

NAND2x1_ASAP7_75t_SL g248 ( 
.A(n_21),
.B(n_227),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_127),
.C(n_184),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_23),
.B(n_128),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_88),
.B1(n_89),
.B2(n_126),
.Y(n_23)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_24),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_42),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_25),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_25),
.A2(n_42),
.B1(n_90),
.B2(n_386),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_35),
.B(n_38),
.Y(n_25)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_26),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_26),
.A2(n_35),
.B1(n_282),
.B2(n_288),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_26),
.A2(n_195),
.B1(n_288),
.B2(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_26),
.A2(n_207),
.B1(n_503),
.B2(n_508),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_26),
.A2(n_518),
.B1(n_543),
.B2(n_555),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_27),
.A2(n_193),
.B1(n_283),
.B2(n_372),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_27),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_29),
.Y(n_323)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_29),
.Y(n_557)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_30),
.Y(n_208)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_33),
.Y(n_521)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_34),
.Y(n_286)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_34),
.Y(n_293)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_34),
.Y(n_376)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_34),
.Y(n_491)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_37),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_38),
.Y(n_209)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_40),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_42),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_67),
.B1(n_78),
.B2(n_79),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_43),
.A2(n_78),
.B1(n_349),
.B2(n_353),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_43),
.A2(n_78),
.B1(n_349),
.B2(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_44),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_44),
.B(n_187),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g244 ( 
.A1(n_44),
.A2(n_175),
.B(n_176),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_44),
.A2(n_175),
.B1(n_187),
.B2(n_311),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_44),
.A2(n_175),
.B1(n_408),
.B2(n_453),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_44),
.A2(n_175),
.B1(n_494),
.B2(n_498),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_44),
.A2(n_175),
.B1(n_453),
.B2(n_498),
.Y(n_512)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_55),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_50),
.Y(n_436)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_51),
.Y(n_537)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_52),
.Y(n_481)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_52),
.Y(n_546)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_59),
.B1(n_62),
.B2(n_66),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_57),
.Y(n_148)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_58),
.Y(n_456)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_64),
.Y(n_483)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_67),
.Y(n_191)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_70),
.Y(n_189)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_71),
.Y(n_351)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_76),
.Y(n_182)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_78),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_78),
.B(n_378),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_79),
.Y(n_174)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_90),
.A2(n_92),
.B(n_126),
.Y(n_228)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_110),
.B1(n_117),
.B2(n_118),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_93),
.A2(n_110),
.B1(n_117),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_93),
.A2(n_117),
.B1(n_118),
.B2(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_93),
.A2(n_117),
.B1(n_296),
.B2(n_301),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_93),
.A2(n_117),
.B1(n_211),
.B2(n_301),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_93),
.A2(n_117),
.B1(n_296),
.B2(n_345),
.Y(n_344)
);

AO21x2_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_98),
.B(n_103),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_94),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_95),
.Y(n_213)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_95),
.Y(n_235)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

AO22x2_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_103)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_105),
.Y(n_243)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_106),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_107),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_107),
.Y(n_277)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_108),
.Y(n_369)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_117),
.B(n_378),
.Y(n_377)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_119),
.Y(n_303)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_121),
.Y(n_216)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_121),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_173),
.B(n_183),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_129),
.B(n_173),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_153),
.B1(n_161),
.B2(n_163),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g218 ( 
.A(n_130),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_130),
.A2(n_161),
.B1(n_257),
.B2(n_262),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_138),
.B(n_144),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_137),
.Y(n_423)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_138),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_142),
.Y(n_342)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_143),
.Y(n_367)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_143),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_147),
.B1(n_149),
.B2(n_152),
.Y(n_144)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_151),
.Y(n_411)
);

BUFx12f_ASAP7_75t_L g497 ( 
.A(n_151),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22x1_ASAP7_75t_SL g217 ( 
.A1(n_154),
.A2(n_162),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_157),
.Y(n_263)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_159),
.Y(n_240)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22x1_ASAP7_75t_L g237 ( 
.A1(n_162),
.A2(n_164),
.B1(n_218),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_162),
.A2(n_218),
.B1(n_219),
.B2(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_162),
.A2(n_218),
.B1(n_336),
.B2(n_343),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_162),
.A2(n_218),
.B1(n_336),
.B2(n_363),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_162),
.A2(n_218),
.B1(n_363),
.B2(n_465),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_169),
.Y(n_472)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_175),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_182),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_183),
.A2(n_230),
.B1(n_246),
.B2(n_247),
.Y(n_229)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_184),
.B(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_210),
.C(n_217),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_185),
.B(n_388),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_190),
.B(n_192),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_186),
.B(n_190),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_192),
.B(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_206),
.B2(n_209),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_193),
.A2(n_372),
.B1(n_429),
.B2(n_437),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_193),
.A2(n_517),
.B1(n_526),
.B2(n_527),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_200),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_201),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_204),
.Y(n_550)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_205),
.Y(n_506)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_210),
.B(n_217),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_213),
.Y(n_299)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_223),
.Y(n_337)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_236),
.B2(n_245),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_235),
.Y(n_347)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_244),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_397),
.B(n_570),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_379),
.C(n_392),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_328),
.B(n_354),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_254),
.B(n_328),
.C(n_572),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_304),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_255),
.B(n_305),
.C(n_307),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_265),
.C(n_294),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_256),
.A2(n_294),
.B1(n_295),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_256),
.Y(n_331)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_257),
.Y(n_343)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_265),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_281),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_266),
.B(n_281),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_273),
.B(n_278),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_286),
.Y(n_525)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_291),
.Y(n_374)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_291),
.Y(n_507)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_324),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_308),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_320),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_309),
.A2(n_310),
.B1(n_320),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_314),
.Y(n_425)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_316),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_316),
.Y(n_500)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_320),
.Y(n_333)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_382),
.C(n_383),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.C(n_334),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_329),
.B(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_334),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_344),
.C(n_348),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_348),
.Y(n_359)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_344),
.B(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_355),
.B(n_357),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.C(n_361),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_361),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_370),
.C(n_377),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_362),
.B(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_365),
.Y(n_364)
);

INVx6_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx6_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_370),
.A2(n_371),
.B1(n_377),
.B2(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_378),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_378),
.B(n_485),
.Y(n_484)
);

OAI21xp33_ASAP7_75t_SL g494 ( 
.A1(n_378),
.A2(n_484),
.B(n_495),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_378),
.B(n_539),
.Y(n_538)
);

A2O1A1O1Ixp25_ASAP7_75t_L g570 ( 
.A1(n_379),
.A2(n_392),
.B(n_571),
.C(n_573),
.D(n_574),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_391),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_380),
.B(n_391),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_381),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_387),
.B1(n_389),
.B2(n_390),
.Y(n_384)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_385),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_390),
.C(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_387),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_395),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_393),
.B(n_395),
.Y(n_574)
);

AOI21x1_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_443),
.B(n_569),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_401),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_399),
.B(n_401),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_406),
.C(n_417),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_402),
.A2(n_403),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_406),
.A2(n_417),
.B1(n_418),
.B2(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_406),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_415),
.Y(n_479)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_427),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_419),
.A2(n_427),
.B1(n_428),
.B2(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_429),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx5_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_442),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_473),
.B(n_568),
.Y(n_443)
);

NOR2xp67_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_449),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_445),
.B(n_449),
.Y(n_568)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.C(n_463),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_450),
.B(n_565),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_452),
.A2(n_463),
.B1(n_464),
.B2(n_566),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_452),
.Y(n_566)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_461),
.Y(n_485)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_467),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_469),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx8_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

AOI21x1_ASAP7_75t_SL g473 ( 
.A1(n_474),
.A2(n_562),
.B(n_567),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_475),
.A2(n_514),
.B(n_561),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_501),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_476),
.B(n_501),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_492),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_477),
.A2(n_492),
.B1(n_493),
.B2(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_477),
.Y(n_529)
);

OAI32xp33_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_480),
.A3(n_482),
.B1(n_484),
.B2(n_486),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_482),
.Y(n_487)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_509),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_502),
.B(n_511),
.C(n_513),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_503),
.Y(n_527)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_511),
.B1(n_512),
.B2(n_513),
.Y(n_509)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_510),
.Y(n_513)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_515),
.A2(n_530),
.B(n_560),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_528),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_516),
.B(n_528),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_531),
.A2(n_553),
.B(n_559),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_542),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_538),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_558),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_554),
.B(n_558),
.Y(n_559)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_564),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_SL g567 ( 
.A(n_563),
.B(n_564),
.Y(n_567)
);


endmodule