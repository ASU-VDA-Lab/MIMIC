module real_aes_2169_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_0), .A2(n_219), .B1(n_554), .B2(n_556), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_1), .A2(n_187), .B1(n_429), .B2(n_430), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_2), .A2(n_83), .B1(n_394), .B2(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_3), .A2(n_184), .B1(n_435), .B2(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_4), .A2(n_117), .B1(n_277), .B2(n_310), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_5), .A2(n_76), .B1(n_344), .B2(n_599), .Y(n_598) );
OA22x2_ASAP7_75t_L g240 ( .A1(n_6), .A2(n_241), .B1(n_242), .B2(n_243), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_6), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_7), .A2(n_54), .B1(n_246), .B2(n_262), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_8), .A2(n_101), .B1(n_413), .B2(n_414), .Y(n_412) );
AO22x2_ASAP7_75t_L g248 ( .A1(n_9), .A2(n_166), .B1(n_249), .B2(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g576 ( .A(n_9), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_10), .A2(n_142), .B1(n_292), .B2(n_293), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_11), .A2(n_141), .B1(n_394), .B2(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_12), .A2(n_64), .B1(n_386), .B2(n_440), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_13), .Y(n_639) );
XOR2x2_ASAP7_75t_L g517 ( .A(n_14), .B(n_518), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_15), .A2(n_81), .B1(n_302), .B2(n_303), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_16), .A2(n_95), .B1(n_296), .B2(n_507), .Y(n_506) );
AO22x2_ASAP7_75t_L g252 ( .A1(n_17), .A2(n_53), .B1(n_249), .B2(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_17), .B(n_575), .Y(n_574) );
OA22x2_ASAP7_75t_L g423 ( .A1(n_18), .A2(n_424), .B1(n_441), .B2(n_442), .Y(n_423) );
INVx1_ASAP7_75t_L g441 ( .A(n_18), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_19), .A2(n_48), .B1(n_369), .B2(n_371), .Y(n_368) );
AOI22xp5_ASAP7_75t_SL g356 ( .A1(n_20), .A2(n_199), .B1(n_357), .B2(n_359), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_21), .A2(n_221), .B1(n_409), .B2(n_411), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_22), .A2(n_130), .B1(n_409), .B2(n_411), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_23), .A2(n_110), .B1(n_246), .B2(n_262), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_24), .B(n_463), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_25), .A2(n_125), .B1(n_341), .B2(n_482), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_26), .A2(n_161), .B1(n_348), .B2(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_27), .A2(n_195), .B1(n_350), .B2(n_386), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_28), .A2(n_154), .B1(n_296), .B2(n_339), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_29), .A2(n_214), .B1(n_369), .B2(n_533), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_30), .A2(n_94), .B1(n_352), .B2(n_440), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_31), .B(n_584), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_32), .Y(n_649) );
OA22x2_ASAP7_75t_L g611 ( .A1(n_33), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_33), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_34), .A2(n_153), .B1(n_404), .B2(n_405), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_35), .B(n_355), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_36), .A2(n_67), .B1(n_296), .B2(n_299), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_37), .A2(n_176), .B1(n_369), .B2(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_38), .A2(n_40), .B1(n_363), .B2(n_394), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_39), .A2(n_177), .B1(n_594), .B2(n_595), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_41), .A2(n_146), .B1(n_299), .B2(n_383), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_42), .A2(n_149), .B1(n_523), .B2(n_524), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_43), .A2(n_133), .B1(n_277), .B2(n_310), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_44), .A2(n_215), .B1(n_624), .B2(n_626), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_45), .A2(n_213), .B1(n_369), .B2(n_417), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_46), .A2(n_182), .B1(n_413), .B2(n_414), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_47), .A2(n_174), .B1(n_586), .B2(n_588), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_49), .A2(n_55), .B1(n_527), .B2(n_528), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_50), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_51), .Y(n_632) );
AOI222xp33_ASAP7_75t_L g419 ( .A1(n_52), .A2(n_57), .B1(n_209), .B2(n_270), .C1(n_392), .C2(n_420), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_56), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_58), .A2(n_169), .B1(n_277), .B2(n_310), .Y(n_309) );
AOI222xp33_ASAP7_75t_L g391 ( .A1(n_59), .A2(n_128), .B1(n_189), .B2(n_363), .C1(n_392), .C2(n_394), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_60), .A2(n_118), .B1(n_359), .B2(n_429), .Y(n_534) );
INVx3_ASAP7_75t_L g249 ( .A(n_61), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_62), .A2(n_127), .B1(n_246), .B2(n_262), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_63), .B(n_314), .Y(n_313) );
XNOR2x2_ASAP7_75t_L g305 ( .A(n_65), .B(n_306), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_66), .A2(n_204), .B1(n_341), .B2(n_344), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_68), .A2(n_192), .B1(n_267), .B2(n_312), .Y(n_311) );
OA22x2_ASAP7_75t_L g399 ( .A1(n_69), .A2(n_400), .B1(n_401), .B2(n_421), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_69), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_70), .A2(n_85), .B1(n_300), .B2(n_348), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_71), .A2(n_103), .B1(n_333), .B2(n_381), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_72), .B(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_73), .A2(n_102), .B1(n_274), .B2(n_277), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_74), .A2(n_126), .B1(n_348), .B2(n_351), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_75), .A2(n_96), .B1(n_333), .B2(n_335), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_77), .A2(n_98), .B1(n_429), .B2(n_430), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_78), .Y(n_633) );
INVx1_ASAP7_75t_SL g257 ( .A(n_79), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_79), .B(n_100), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_80), .Y(n_618) );
INVx2_ASAP7_75t_L g232 ( .A(n_82), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_84), .A2(n_137), .B1(n_293), .B2(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_86), .A2(n_208), .B1(n_288), .B2(n_289), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_87), .B(n_355), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_88), .A2(n_180), .B1(n_267), .B2(n_270), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_89), .A2(n_121), .B1(n_369), .B2(n_417), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_90), .A2(n_113), .B1(n_591), .B2(n_620), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_91), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_92), .A2(n_135), .B1(n_299), .B2(n_435), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_93), .A2(n_193), .B1(n_300), .B2(n_341), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_97), .A2(n_191), .B1(n_296), .B2(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_99), .A2(n_138), .B1(n_337), .B2(n_437), .Y(n_436) );
AO22x2_ASAP7_75t_L g260 ( .A1(n_100), .A2(n_170), .B1(n_249), .B2(n_261), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_104), .Y(n_469) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_105), .A2(n_210), .B1(n_394), .B2(n_536), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_106), .A2(n_159), .B1(n_363), .B2(n_394), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_107), .A2(n_163), .B1(n_292), .B2(n_293), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_108), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_109), .A2(n_150), .B1(n_482), .B2(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_111), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_112), .A2(n_131), .B1(n_296), .B2(n_386), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_114), .A2(n_148), .B1(n_386), .B2(n_440), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_115), .A2(n_190), .B1(n_369), .B2(n_427), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_116), .A2(n_212), .B1(n_333), .B2(n_381), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_119), .A2(n_157), .B1(n_484), .B2(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_120), .A2(n_216), .B1(n_590), .B2(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g258 ( .A(n_122), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_123), .B(n_280), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_124), .A2(n_151), .B1(n_357), .B2(n_477), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_129), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_132), .A2(n_143), .B1(n_320), .B2(n_321), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_134), .A2(n_140), .B1(n_288), .B2(n_289), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_136), .A2(n_200), .B1(n_601), .B2(n_602), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_139), .A2(n_156), .B1(n_405), .B2(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_144), .A2(n_218), .B1(n_292), .B2(n_293), .Y(n_316) );
AOI22xp33_ASAP7_75t_SL g487 ( .A1(n_145), .A2(n_172), .B1(n_296), .B2(n_488), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_147), .A2(n_171), .B1(n_333), .B2(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_152), .B(n_280), .Y(n_279) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_155), .A2(n_160), .B1(n_357), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_158), .A2(n_217), .B1(n_551), .B2(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_162), .B(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_SL g499 ( .A1(n_164), .A2(n_173), .B1(n_437), .B2(n_500), .Y(n_499) );
XNOR2x1_ASAP7_75t_L g545 ( .A(n_165), .B(n_546), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_167), .A2(n_181), .B1(n_274), .B2(n_277), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_168), .A2(n_220), .B1(n_531), .B2(n_533), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_175), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_178), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_179), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g572 ( .A(n_179), .Y(n_572) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_183), .A2(n_223), .B(n_233), .C(n_578), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_185), .A2(n_206), .B1(n_302), .B2(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g229 ( .A(n_186), .Y(n_229) );
AND2x2_ASAP7_75t_R g608 ( .A(n_186), .B(n_572), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_188), .A2(n_207), .B1(n_430), .B2(n_628), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_194), .A2(n_202), .B1(n_417), .B2(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_196), .A2(n_205), .B1(n_363), .B2(n_365), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_197), .B(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_198), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_201), .A2(n_580), .B1(n_581), .B2(n_606), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_201), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_203), .B(n_394), .Y(n_465) );
AO22x1_ASAP7_75t_L g471 ( .A1(n_211), .A2(n_472), .B1(n_489), .B2(n_490), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_211), .Y(n_489) );
CKINVDCx6p67_ASAP7_75t_R g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
BUFx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_SL g226 ( .A(n_227), .B(n_230), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g661 ( .A(n_228), .B(n_230), .Y(n_661) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_229), .B(n_572), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_444), .B1(n_567), .B2(n_568), .C(n_569), .Y(n_233) );
INVx1_ASAP7_75t_L g567 ( .A(n_234), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B1(n_323), .B2(n_324), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B1(n_304), .B2(n_322), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2x1_ASAP7_75t_L g243 ( .A(n_244), .B(n_285), .Y(n_243) );
NAND4xp25_ASAP7_75t_L g244 ( .A(n_245), .B(n_266), .C(n_273), .D(n_279), .Y(n_244) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_254), .Y(n_246) );
AND2x2_ASAP7_75t_L g288 ( .A(n_247), .B(n_275), .Y(n_288) );
AND2x6_ASAP7_75t_L g293 ( .A(n_247), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g334 ( .A(n_247), .B(n_275), .Y(n_334) );
AND2x4_ASAP7_75t_L g346 ( .A(n_247), .B(n_294), .Y(n_346) );
AND2x2_ASAP7_75t_L g370 ( .A(n_247), .B(n_254), .Y(n_370) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_251), .Y(n_247) );
INVx2_ASAP7_75t_L g269 ( .A(n_248), .Y(n_269) );
AND2x2_ASAP7_75t_L g272 ( .A(n_248), .B(n_252), .Y(n_272) );
INVx1_ASAP7_75t_L g250 ( .A(n_249), .Y(n_250) );
INVx2_ASAP7_75t_L g253 ( .A(n_249), .Y(n_253) );
OAI22x1_ASAP7_75t_L g255 ( .A1(n_249), .A2(n_256), .B1(n_257), .B2(n_258), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_249), .Y(n_256) );
INVx1_ASAP7_75t_L g261 ( .A(n_249), .Y(n_261) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_251), .Y(n_264) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g268 ( .A(n_252), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g284 ( .A(n_252), .Y(n_284) );
AND2x4_ASAP7_75t_L g267 ( .A(n_254), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g302 ( .A(n_254), .B(n_283), .Y(n_302) );
AND2x4_ASAP7_75t_L g350 ( .A(n_254), .B(n_283), .Y(n_350) );
AND2x2_ASAP7_75t_L g364 ( .A(n_254), .B(n_268), .Y(n_364) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_259), .Y(n_254) );
AND2x2_ASAP7_75t_L g265 ( .A(n_255), .B(n_260), .Y(n_265) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_255), .Y(n_271) );
INVx2_ASAP7_75t_L g276 ( .A(n_255), .Y(n_276) );
AND2x4_ASAP7_75t_L g294 ( .A(n_259), .B(n_276), .Y(n_294) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g275 ( .A(n_260), .B(n_276), .Y(n_275) );
BUFx2_ASAP7_75t_L g290 ( .A(n_260), .Y(n_290) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
AND2x4_ASAP7_75t_L g373 ( .A(n_263), .B(n_265), .Y(n_373) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g277 ( .A(n_265), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g282 ( .A(n_265), .B(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g361 ( .A(n_265), .B(n_278), .Y(n_361) );
AND2x4_ASAP7_75t_L g393 ( .A(n_265), .B(n_283), .Y(n_393) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_267), .Y(n_420) );
AND2x2_ASAP7_75t_L g274 ( .A(n_268), .B(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g300 ( .A(n_268), .B(n_294), .Y(n_300) );
AND2x2_ASAP7_75t_L g310 ( .A(n_268), .B(n_275), .Y(n_310) );
AND2x2_ASAP7_75t_L g321 ( .A(n_268), .B(n_294), .Y(n_321) );
AND2x4_ASAP7_75t_L g358 ( .A(n_268), .B(n_275), .Y(n_358) );
INVxp67_ASAP7_75t_L g278 ( .A(n_269), .Y(n_278) );
AND2x4_ASAP7_75t_L g283 ( .A(n_269), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_SL g270 ( .A(n_271), .B(n_272), .Y(n_270) );
AND2x2_ASAP7_75t_SL g312 ( .A(n_271), .B(n_272), .Y(n_312) );
AND2x2_ASAP7_75t_L g367 ( .A(n_271), .B(n_272), .Y(n_367) );
AND2x4_ASAP7_75t_L g289 ( .A(n_272), .B(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g303 ( .A(n_272), .B(n_294), .Y(n_303) );
AND2x4_ASAP7_75t_L g337 ( .A(n_272), .B(n_290), .Y(n_337) );
AND2x4_ASAP7_75t_L g352 ( .A(n_272), .B(n_294), .Y(n_352) );
AND2x6_ASAP7_75t_L g292 ( .A(n_275), .B(n_283), .Y(n_292) );
AND2x2_ASAP7_75t_L g343 ( .A(n_275), .B(n_283), .Y(n_343) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_280), .Y(n_565) );
INVx3_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
INVx4_ASAP7_75t_SL g314 ( .A(n_281), .Y(n_314) );
INVx4_ASAP7_75t_SL g355 ( .A(n_281), .Y(n_355) );
INVx3_ASAP7_75t_L g538 ( .A(n_281), .Y(n_538) );
INVx6_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g298 ( .A(n_283), .B(n_294), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_295), .C(n_301), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_291), .Y(n_286) );
INVx1_ASAP7_75t_L g503 ( .A(n_292), .Y(n_503) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx4_ASAP7_75t_L g320 ( .A(n_297), .Y(n_320) );
INVx3_ASAP7_75t_SL g383 ( .A(n_297), .Y(n_383) );
INVx2_ASAP7_75t_L g435 ( .A(n_297), .Y(n_435) );
INVx2_ASAP7_75t_SL g527 ( .A(n_297), .Y(n_527) );
INVx2_ASAP7_75t_SL g558 ( .A(n_297), .Y(n_558) );
INVx8_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g634 ( .A(n_299), .Y(n_634) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_300), .Y(n_339) );
BUFx3_ASAP7_75t_L g405 ( .A(n_300), .Y(n_405) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_300), .Y(n_488) );
INVx2_ASAP7_75t_L g508 ( .A(n_300), .Y(n_508) );
INVx1_ASAP7_75t_SL g322 ( .A(n_304), .Y(n_322) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_315), .Y(n_306) );
NAND4xp25_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .C(n_311), .D(n_313), .Y(n_307) );
BUFx2_ASAP7_75t_L g584 ( .A(n_314), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .C(n_318), .D(n_319), .Y(n_315) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI22xp5_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_326), .B1(n_396), .B2(n_443), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI22xp33_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_328), .B1(n_375), .B2(n_376), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
XNOR2x1_ASAP7_75t_L g329 ( .A(n_330), .B(n_374), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_353), .Y(n_330) );
NAND4xp25_ASAP7_75t_L g331 ( .A(n_332), .B(n_338), .C(n_340), .D(n_347), .Y(n_331) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g410 ( .A(n_334), .Y(n_410) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g411 ( .A(n_336), .Y(n_411) );
INVx2_ASAP7_75t_L g602 ( .A(n_336), .Y(n_602) );
OAI22xp33_ASAP7_75t_SL g650 ( .A1(n_336), .A2(n_651), .B1(n_654), .B2(n_655), .Y(n_650) );
INVx5_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
BUFx3_ASAP7_75t_L g381 ( .A(n_337), .Y(n_381) );
BUFx2_ASAP7_75t_L g500 ( .A(n_337), .Y(n_500) );
BUFx2_ASAP7_75t_L g556 ( .A(n_337), .Y(n_556) );
BUFx2_ASAP7_75t_L g645 ( .A(n_341), .Y(n_645) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_SL g551 ( .A(n_342), .Y(n_551) );
INVx3_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g413 ( .A(n_343), .Y(n_413) );
BUFx2_ASAP7_75t_L g521 ( .A(n_343), .Y(n_521) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g414 ( .A(n_345), .Y(n_414) );
INVx2_ASAP7_75t_SL g457 ( .A(n_345), .Y(n_457) );
INVx2_ASAP7_75t_L g482 ( .A(n_345), .Y(n_482) );
INVx1_ASAP7_75t_SL g552 ( .A(n_345), .Y(n_552) );
INVx2_ASAP7_75t_L g648 ( .A(n_345), .Y(n_648) );
INVx8_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g523 ( .A(n_349), .Y(n_523) );
INVx2_ASAP7_75t_L g549 ( .A(n_349), .Y(n_549) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_349), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_631) );
INVx6_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx3_ASAP7_75t_L g404 ( .A(n_350), .Y(n_404) );
BUFx3_ASAP7_75t_L g440 ( .A(n_350), .Y(n_440) );
BUFx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g386 ( .A(n_352), .Y(n_386) );
INVx2_ASAP7_75t_L g485 ( .A(n_352), .Y(n_485) );
BUFx2_ASAP7_75t_SL g641 ( .A(n_352), .Y(n_641) );
NAND4xp25_ASAP7_75t_SL g353 ( .A(n_354), .B(n_356), .C(n_362), .D(n_368), .Y(n_353) );
BUFx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx3_ASAP7_75t_L g429 ( .A(n_358), .Y(n_429) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_358), .Y(n_629) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g430 ( .A(n_360), .Y(n_430) );
INVx2_ASAP7_75t_L g477 ( .A(n_360), .Y(n_477) );
INVx2_ASAP7_75t_SL g562 ( .A(n_360), .Y(n_562) );
INVx2_ASAP7_75t_L g588 ( .A(n_360), .Y(n_588) );
INVx6_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_363), .Y(n_590) );
BUFx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g464 ( .A(n_364), .Y(n_464) );
BUFx5_ASAP7_75t_L g536 ( .A(n_364), .Y(n_536) );
BUFx3_ASAP7_75t_L g621 ( .A(n_364), .Y(n_621) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx3_ASAP7_75t_L g592 ( .A(n_366), .Y(n_592) );
INVx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx12f_ASAP7_75t_L g394 ( .A(n_367), .Y(n_394) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_370), .Y(n_515) );
INVx3_ASAP7_75t_L g532 ( .A(n_370), .Y(n_532) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx6f_ASAP7_75t_SL g417 ( .A(n_373), .Y(n_417) );
BUFx3_ASAP7_75t_L g427 ( .A(n_373), .Y(n_427) );
BUFx4f_ASAP7_75t_L g533 ( .A(n_373), .Y(n_533) );
INVx2_ASAP7_75t_L g596 ( .A(n_373), .Y(n_596) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
XOR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_395), .Y(n_377) );
NAND4xp75_ASAP7_75t_L g378 ( .A(n_379), .B(n_384), .C(n_388), .D(n_391), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_386), .Y(n_604) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
BUFx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_SL g461 ( .A(n_393), .Y(n_461) );
INVx1_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AO22x1_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_422), .B2(n_423), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g421 ( .A(n_401), .Y(n_421) );
NAND4xp75_ASAP7_75t_L g401 ( .A(n_402), .B(n_407), .C(n_415), .D(n_419), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_406), .Y(n_402) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_412), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g437 ( .A(n_410), .Y(n_437) );
INVx2_ASAP7_75t_L g555 ( .A(n_410), .Y(n_555) );
BUFx3_ASAP7_75t_L g599 ( .A(n_413), .Y(n_599) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g442 ( .A(n_424), .Y(n_442) );
NOR2x1_ASAP7_75t_L g424 ( .A(n_425), .B(n_433), .Y(n_424) );
NAND4xp25_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .C(n_431), .D(n_432), .Y(n_425) );
BUFx6f_ASAP7_75t_SL g626 ( .A(n_427), .Y(n_626) );
INVx1_ASAP7_75t_L g587 ( .A(n_429), .Y(n_587) );
NAND4xp25_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .C(n_438), .D(n_439), .Y(n_433) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_437), .Y(n_601) );
INVx1_ASAP7_75t_L g568 ( .A(n_444), .Y(n_568) );
XOR2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_492), .Y(n_444) );
OAI22xp33_ASAP7_75t_R g445 ( .A1(n_446), .A2(n_447), .B1(n_470), .B2(n_491), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
XOR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_469), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_458), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_452), .B(n_453), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_466), .Y(n_458) );
OAI211xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B(n_462), .C(n_465), .Y(n_459) );
OAI21xp5_ASAP7_75t_SL g510 ( .A1(n_461), .A2(n_511), .B(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g475 ( .A(n_464), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g491 ( .A(n_470), .Y(n_491) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_SL g490 ( .A(n_472), .Y(n_490) );
NOR2x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_480), .Y(n_472) );
NAND4xp25_ASAP7_75t_L g473 ( .A(n_474), .B(n_476), .C(n_478), .D(n_479), .Y(n_473) );
NAND4xp25_ASAP7_75t_L g480 ( .A(n_481), .B(n_483), .C(n_486), .D(n_487), .Y(n_480) );
INVx2_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g524 ( .A(n_485), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_541), .B1(n_542), .B2(n_566), .Y(n_492) );
INVx2_ASAP7_75t_L g566 ( .A(n_493), .Y(n_566) );
OA22x2_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_517), .B1(n_539), .B2(n_540), .Y(n_493) );
INVxp67_ASAP7_75t_SL g540 ( .A(n_494), .Y(n_540) );
XNOR2x1_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
NAND2x1p5_ASAP7_75t_L g496 ( .A(n_497), .B(n_509), .Y(n_496) );
NOR2x1_ASAP7_75t_L g497 ( .A(n_498), .B(n_504), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g528 ( .A(n_508), .Y(n_528) );
NOR2x1_ASAP7_75t_L g509 ( .A(n_510), .B(n_513), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .Y(n_513) );
BUFx6f_ASAP7_75t_SL g594 ( .A(n_515), .Y(n_594) );
INVx1_ASAP7_75t_L g539 ( .A(n_517), .Y(n_539) );
NOR2xp67_ASAP7_75t_L g518 ( .A(n_519), .B(n_529), .Y(n_518) );
NAND4xp25_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .C(n_525), .D(n_526), .Y(n_519) );
BUFx2_ASAP7_75t_L g638 ( .A(n_527), .Y(n_638) );
NAND4xp25_ASAP7_75t_L g529 ( .A(n_530), .B(n_534), .C(n_535), .D(n_537), .Y(n_529) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g625 ( .A(n_532), .Y(n_625) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_559), .Y(n_546) );
NAND4xp25_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .C(n_553), .D(n_557), .Y(n_547) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g653 ( .A(n_555), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .C(n_563), .D(n_564), .Y(n_559) );
INVx3_ASAP7_75t_L g617 ( .A(n_565), .Y(n_617) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_571), .B(n_574), .Y(n_658) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
OAI222xp33_ASAP7_75t_R g578 ( .A1(n_579), .A2(n_607), .B1(n_609), .B2(n_612), .C1(n_656), .C2(n_659), .Y(n_578) );
INVx2_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_597), .Y(n_581) );
NAND4xp25_ASAP7_75t_SL g582 ( .A(n_583), .B(n_585), .C(n_589), .D(n_593), .Y(n_582) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND4xp25_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .C(n_603), .D(n_605), .Y(n_597) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND3x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_630), .C(n_642), .Y(n_614) );
NOR2xp67_ASAP7_75t_SL g615 ( .A(n_616), .B(n_622), .Y(n_615) );
OAI21xp5_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_618), .B(n_619), .Y(n_616) );
BUFx6f_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_623), .B(n_627), .Y(n_622) );
BUFx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_635), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_639), .B2(n_640), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_650), .Y(n_642) );
OAI22xp33_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_646), .B1(n_647), .B2(n_649), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_657), .Y(n_656) );
CKINVDCx6p67_ASAP7_75t_R g657 ( .A(n_658), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_660), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_661), .Y(n_660) );
endmodule