module fake_netlist_6_4582_n_1277 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1277);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1277;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1249;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1272;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_236;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_172),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_155),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_46),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_98),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_52),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_40),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_76),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_88),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_46),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_97),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_2),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_86),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_16),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_77),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_103),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_130),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_57),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_162),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_4),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_116),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_179),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_138),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_100),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_173),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_121),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_134),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_133),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_122),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_73),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_1),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_17),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_72),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_3),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_63),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_148),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_8),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_66),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_37),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_9),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_79),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_3),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_91),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_143),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_36),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_168),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_78),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_21),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_59),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_27),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_56),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_152),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_114),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_60),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_175),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_81),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_39),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_80),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_90),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_144),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_33),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_101),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_2),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_94),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_123),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_21),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_70),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_108),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_99),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_151),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_37),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_164),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_45),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_62),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_132),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_48),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_135),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_31),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_38),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_1),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_32),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_92),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_0),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_171),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_18),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_112),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_5),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_154),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_10),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_174),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_83),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_85),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_156),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_107),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_82),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_27),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_18),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_50),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_0),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_28),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_54),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_180),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_140),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_40),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_65),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_16),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_75),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_74),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_128),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_166),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_51),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_87),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_30),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_96),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_42),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_221),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_194),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_295),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_4),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_221),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_197),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_253),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_191),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_220),
.Y(n_314)
);

AND2x6_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_58),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_210),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_258),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_226),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_211),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_212),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_213),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_229),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_214),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_247),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_196),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_296),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_215),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_187),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_271),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_258),
.Y(n_331)
);

INVxp33_ASAP7_75t_SL g332 ( 
.A(n_187),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_189),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_189),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_190),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_201),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_196),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_201),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_190),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_288),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_288),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_200),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_202),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_208),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_209),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_218),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_222),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_217),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_237),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_219),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_R g355 ( 
.A(n_206),
.B(n_61),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_239),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_249),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_290),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_301),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_301),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_305),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_228),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_250),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_252),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_251),
.B(n_5),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_262),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_205),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_264),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_207),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_272),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_199),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_223),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_291),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_199),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_224),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_L g376 ( 
.A(n_251),
.B(n_6),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_231),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_216),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_234),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_225),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_238),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_240),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_216),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_241),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_230),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_232),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_256),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_232),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_236),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_258),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_233),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_236),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_242),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_244),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_245),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_261),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_308),
.A2(n_280),
.B1(n_287),
.B2(n_286),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_293),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

INVx6_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_313),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_311),
.B(n_185),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_315),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_315),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_314),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_315),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g407 ( 
.A1(n_371),
.A2(n_297),
.B(n_293),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_322),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_317),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_307),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_373),
.B(n_185),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_324),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_315),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_316),
.B(n_319),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_392),
.B(n_297),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

OA21x2_ASAP7_75t_L g418 ( 
.A1(n_374),
.A2(n_383),
.B(n_378),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_320),
.B(n_246),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_344),
.B(n_283),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_315),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_386),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_321),
.B(n_323),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_328),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_328),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_330),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_388),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_369),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_325),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_325),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_331),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_345),
.B(n_283),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_377),
.B(n_186),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_307),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_346),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_347),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_331),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_340),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_327),
.B(n_274),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_348),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_352),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_356),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_390),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_333),
.A2(n_255),
.B1(n_302),
.B2(n_227),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_390),
.Y(n_447)
);

AND2x6_ASAP7_75t_L g448 ( 
.A(n_357),
.B(n_283),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_332),
.B(n_334),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_351),
.B(n_248),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_364),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_366),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_368),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_349),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_370),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_337),
.B(n_289),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_354),
.B(n_254),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_341),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_396),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_312),
.B(n_235),
.Y(n_461)
);

OAI21xp33_ASAP7_75t_L g462 ( 
.A1(n_309),
.A2(n_289),
.B(n_266),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_306),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_310),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_318),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_365),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_411),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_438),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_438),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_399),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_445),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_445),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_403),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_399),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_440),
.B(n_375),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_447),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_432),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_398),
.B(n_376),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_447),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_419),
.B(n_380),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_439),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_432),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_432),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_409),
.B(n_258),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_409),
.B(n_418),
.Y(n_486)
);

BUFx4f_ASAP7_75t_L g487 ( 
.A(n_403),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_447),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_409),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_465),
.B(n_385),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_409),
.B(n_258),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_410),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_462),
.A2(n_339),
.B1(n_292),
.B2(n_285),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_418),
.Y(n_494)
);

NAND3xp33_ASAP7_75t_L g495 ( 
.A(n_462),
.B(n_336),
.C(n_382),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_SL g496 ( 
.A(n_412),
.B(n_367),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_447),
.Y(n_497)
);

NAND2xp33_ASAP7_75t_SL g498 ( 
.A(n_428),
.B(n_367),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_447),
.Y(n_499)
);

AO22x2_ASAP7_75t_L g500 ( 
.A1(n_397),
.A2(n_282),
.B1(n_353),
.B2(n_338),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_455),
.B(n_391),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_418),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_447),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_418),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_435),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_407),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_398),
.B(n_258),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_398),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_457),
.B(n_465),
.Y(n_509)
);

BUFx6f_ASAP7_75t_SL g510 ( 
.A(n_403),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_398),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_465),
.Y(n_512)
);

OAI22xp33_ASAP7_75t_L g513 ( 
.A1(n_446),
.A2(n_263),
.B1(n_269),
.B2(n_268),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_457),
.B(n_393),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_407),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_459),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_459),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_416),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_403),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_463),
.Y(n_521)
);

BUFx10_ASAP7_75t_L g522 ( 
.A(n_400),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_463),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_451),
.B(n_394),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_463),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_416),
.B(n_258),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g527 ( 
.A(n_407),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_416),
.B(n_258),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_463),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_415),
.B(n_283),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_416),
.B(n_395),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_466),
.B(n_273),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_420),
.B(n_285),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_464),
.B(n_285),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_463),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_422),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_511),
.B(n_458),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_505),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_467),
.Y(n_540)
);

A2O1A1Ixp33_ASAP7_75t_L g541 ( 
.A1(n_511),
.A2(n_508),
.B(n_519),
.C(n_475),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_470),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_511),
.B(n_423),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_467),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_470),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_508),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_508),
.B(n_453),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_L g548 ( 
.A(n_531),
.B(n_403),
.Y(n_548)
);

NOR3xp33_ASAP7_75t_L g549 ( 
.A(n_513),
.B(n_402),
.C(n_449),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_519),
.B(n_453),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_519),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_531),
.A2(n_243),
.B1(n_434),
.B2(n_400),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_512),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_512),
.B(n_355),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_481),
.B(n_453),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_514),
.B(n_403),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_479),
.B(n_453),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_516),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_501),
.B(n_372),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_L g560 ( 
.A(n_506),
.B(n_404),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_495),
.B(n_514),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_506),
.B(n_404),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_514),
.B(n_404),
.Y(n_563)
);

O2A1O1Ixp33_ASAP7_75t_L g564 ( 
.A1(n_494),
.A2(n_442),
.B(n_436),
.C(n_437),
.Y(n_564)
);

BUFx5_ASAP7_75t_L g565 ( 
.A(n_522),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_495),
.B(n_372),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_470),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_509),
.B(n_464),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_473),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_479),
.B(n_527),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_479),
.A2(n_387),
.B1(n_396),
.B2(n_384),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_SL g572 ( 
.A(n_501),
.B(n_379),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_494),
.A2(n_404),
.B1(n_421),
.B2(n_414),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_473),
.Y(n_574)
);

O2A1O1Ixp33_ASAP7_75t_L g575 ( 
.A1(n_502),
.A2(n_441),
.B(n_436),
.C(n_437),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_516),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_527),
.B(n_453),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_490),
.B(n_379),
.Y(n_578)
);

OAI22xp33_ASAP7_75t_L g579 ( 
.A1(n_513),
.A2(n_446),
.B1(n_466),
.B2(n_361),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_509),
.A2(n_381),
.B1(n_387),
.B2(n_384),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_517),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_482),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_482),
.B(n_460),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_509),
.B(n_456),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_506),
.B(n_456),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_493),
.B(n_404),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_532),
.B(n_493),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_515),
.B(n_404),
.Y(n_588)
);

A2O1A1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_502),
.A2(n_433),
.B(n_420),
.C(n_454),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_L g590 ( 
.A1(n_532),
.A2(n_358),
.B1(n_360),
.B2(n_359),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_524),
.A2(n_400),
.B1(n_381),
.B2(n_192),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_487),
.B(n_406),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_477),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_515),
.B(n_518),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_504),
.B(n_333),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_517),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_496),
.A2(n_359),
.B1(n_361),
.B2(n_360),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_515),
.B(n_456),
.Y(n_598)
);

INVx8_ASAP7_75t_L g599 ( 
.A(n_530),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_518),
.B(n_456),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_518),
.B(n_456),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_504),
.B(n_486),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_477),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_537),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_537),
.Y(n_605)
);

OR2x2_ASAP7_75t_SL g606 ( 
.A(n_500),
.B(n_461),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_533),
.B(n_430),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_487),
.B(n_406),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_486),
.B(n_456),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_487),
.B(n_406),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_507),
.B(n_338),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_537),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_487),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_530),
.A2(n_400),
.B1(n_188),
.B2(n_192),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_497),
.B(n_499),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_477),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_497),
.B(n_463),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_535),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_533),
.B(n_430),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_507),
.B(n_342),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_500),
.A2(n_343),
.B1(n_342),
.B2(n_358),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_535),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_497),
.B(n_420),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_SL g624 ( 
.A(n_510),
.B(n_343),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_526),
.B(n_441),
.Y(n_625)
);

O2A1O1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_526),
.A2(n_450),
.B(n_452),
.C(n_444),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_499),
.B(n_420),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_492),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_478),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_498),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_528),
.B(n_442),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_528),
.B(n_443),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_499),
.B(n_433),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_473),
.B(n_406),
.Y(n_634)
);

AOI21x1_ASAP7_75t_L g635 ( 
.A1(n_592),
.A2(n_610),
.B(n_608),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_560),
.A2(n_520),
.B(n_530),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_553),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_602),
.A2(n_520),
.B(n_503),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_613),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_562),
.A2(n_520),
.B(n_530),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_588),
.A2(n_520),
.B(n_530),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_553),
.Y(n_642)
);

O2A1O1Ixp33_ASAP7_75t_L g643 ( 
.A1(n_561),
.A2(n_534),
.B(n_452),
.C(n_443),
.Y(n_643)
);

AO21x1_ASAP7_75t_L g644 ( 
.A1(n_561),
.A2(n_534),
.B(n_491),
.Y(n_644)
);

AOI33xp33_ASAP7_75t_L g645 ( 
.A1(n_590),
.A2(n_401),
.A3(n_429),
.B1(n_426),
.B2(n_417),
.B3(n_413),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_587),
.B(n_503),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_613),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_609),
.A2(n_530),
.B(n_503),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_555),
.A2(n_510),
.B(n_522),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_546),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_540),
.B(n_424),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_543),
.B(n_476),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_568),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_613),
.B(n_406),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_546),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_625),
.B(n_476),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_544),
.B(n_425),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_611),
.B(n_461),
.C(n_425),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_568),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_611),
.A2(n_500),
.B1(n_535),
.B2(n_529),
.Y(n_660)
);

A2O1A1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_625),
.A2(n_485),
.B(n_491),
.C(n_489),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_577),
.A2(n_510),
.B(n_522),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_618),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_L g664 ( 
.A(n_565),
.B(n_414),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_631),
.B(n_476),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_613),
.B(n_414),
.Y(n_666)
);

O2A1O1Ixp33_ASAP7_75t_L g667 ( 
.A1(n_595),
.A2(n_450),
.B(n_454),
.C(n_444),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_604),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_607),
.B(n_500),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_586),
.A2(n_489),
.B(n_480),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_619),
.B(n_500),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_546),
.B(n_522),
.Y(n_672)
);

AO21x1_ASAP7_75t_L g673 ( 
.A1(n_549),
.A2(n_485),
.B(n_521),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_631),
.B(n_476),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_585),
.A2(n_510),
.B(n_488),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_632),
.B(n_480),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_632),
.B(n_480),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_538),
.B(n_480),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_628),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_598),
.A2(n_488),
.B(n_521),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_594),
.B(n_488),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_620),
.B(n_488),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_620),
.B(n_570),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_600),
.A2(n_525),
.B(n_523),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_601),
.A2(n_525),
.B(n_523),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_L g686 ( 
.A1(n_541),
.A2(n_474),
.B(n_478),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_R g687 ( 
.A(n_624),
.B(n_312),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_582),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_584),
.B(n_468),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_546),
.Y(n_690)
);

A2O1A1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_549),
.A2(n_468),
.B(n_469),
.C(n_471),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_551),
.B(n_414),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_595),
.B(n_326),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_566),
.B(n_326),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_573),
.B(n_469),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_604),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_573),
.B(n_414),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_548),
.A2(n_574),
.B(n_569),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_569),
.A2(n_536),
.B(n_529),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_574),
.A2(n_536),
.B(n_421),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_551),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_551),
.B(n_414),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_622),
.B(n_471),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_551),
.B(n_421),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_558),
.B(n_472),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_576),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_557),
.A2(n_421),
.B(n_472),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_566),
.A2(n_474),
.B(n_433),
.C(n_484),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g709 ( 
.A1(n_589),
.A2(n_483),
.B(n_478),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_579),
.B(n_401),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_552),
.B(n_421),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_539),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_SL g713 ( 
.A(n_559),
.B(n_186),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_581),
.B(n_484),
.Y(n_714)
);

O2A1O1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_564),
.A2(n_426),
.B(n_408),
.C(n_413),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_556),
.B(n_405),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_579),
.B(n_405),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_563),
.A2(n_188),
.B1(n_193),
.B2(n_195),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_547),
.A2(n_483),
.B(n_427),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_596),
.B(n_422),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_575),
.B(n_427),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_550),
.A2(n_292),
.B(n_285),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_634),
.A2(n_292),
.B(n_285),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_542),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_554),
.B(n_257),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_605),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_623),
.A2(n_292),
.B(n_408),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_545),
.Y(n_728)
);

OR2x6_ASAP7_75t_L g729 ( 
.A(n_599),
.B(n_630),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_626),
.B(n_259),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_612),
.A2(n_292),
.B1(n_429),
.B2(n_417),
.Y(n_731)
);

INVxp67_ASAP7_75t_SL g732 ( 
.A(n_639),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_693),
.B(n_642),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_668),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_637),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_639),
.Y(n_736)
);

CKINVDCx8_ASAP7_75t_R g737 ( 
.A(n_712),
.Y(n_737)
);

INVx3_ASAP7_75t_SL g738 ( 
.A(n_679),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_693),
.B(n_580),
.Y(n_739)
);

CKINVDCx14_ASAP7_75t_R g740 ( 
.A(n_687),
.Y(n_740)
);

OAI22x1_ASAP7_75t_L g741 ( 
.A1(n_694),
.A2(n_621),
.B1(n_597),
.B2(n_658),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_642),
.B(n_578),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_706),
.Y(n_743)
);

NOR2xp67_ASAP7_75t_L g744 ( 
.A(n_725),
.B(n_591),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_663),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_637),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_683),
.A2(n_578),
.B(n_590),
.C(n_614),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_653),
.B(n_583),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_659),
.B(n_571),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_687),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_639),
.B(n_572),
.Y(n_751)
);

O2A1O1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_667),
.A2(n_633),
.B(n_627),
.C(n_615),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_664),
.A2(n_565),
.B(n_599),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_696),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_724),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_690),
.Y(n_756)
);

CKINVDCx14_ASAP7_75t_R g757 ( 
.A(n_651),
.Y(n_757)
);

AO32x1_ASAP7_75t_L g758 ( 
.A1(n_669),
.A2(n_629),
.A3(n_567),
.B1(n_616),
.B2(n_593),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_638),
.A2(n_565),
.B(n_617),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_661),
.A2(n_603),
.B(n_448),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_R g761 ( 
.A(n_688),
.B(n_599),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_636),
.A2(n_565),
.B(n_431),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_640),
.A2(n_565),
.B(n_431),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_694),
.B(n_606),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_646),
.B(n_565),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_657),
.Y(n_766)
);

O2A1O1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_710),
.A2(n_275),
.B(n_277),
.C(n_279),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_680),
.A2(n_111),
.B(n_184),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_690),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_639),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_724),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_671),
.B(n_193),
.Y(n_772)
);

INVx3_ASAP7_75t_SL g773 ( 
.A(n_729),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_713),
.A2(n_278),
.B1(n_260),
.B2(n_265),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_689),
.B(n_195),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_729),
.B(n_64),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_R g777 ( 
.A(n_655),
.B(n_198),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_682),
.B(n_198),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_729),
.B(n_650),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_728),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_690),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_641),
.A2(n_284),
.B(n_267),
.Y(n_782)
);

OAI21x1_ASAP7_75t_L g783 ( 
.A1(n_684),
.A2(n_102),
.B(n_183),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_650),
.B(n_655),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_726),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_710),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_690),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_656),
.B(n_203),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_665),
.B(n_203),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_705),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_701),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_647),
.B(n_204),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_698),
.A2(n_281),
.B(n_304),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_701),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_717),
.B(n_204),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_701),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_717),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_674),
.B(n_298),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_676),
.B(n_298),
.Y(n_799)
);

INVx5_ASAP7_75t_L g800 ( 
.A(n_647),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_677),
.A2(n_304),
.B(n_300),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_660),
.A2(n_300),
.B1(n_299),
.B2(n_448),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_SL g803 ( 
.A(n_647),
.B(n_299),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_648),
.A2(n_448),
.B(n_89),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_643),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_762),
.A2(n_686),
.B(n_675),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_762),
.A2(n_685),
.B(n_709),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_790),
.B(n_645),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_766),
.B(n_720),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_738),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_739),
.A2(n_716),
.B1(n_673),
.B2(n_718),
.Y(n_811)
);

NOR2x1_ASAP7_75t_L g812 ( 
.A(n_794),
.B(n_701),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_764),
.A2(n_716),
.B1(n_711),
.B2(n_730),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_795),
.A2(n_741),
.B1(n_786),
.B2(n_742),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_759),
.A2(n_649),
.B(n_662),
.Y(n_815)
);

BUFx12f_ASAP7_75t_L g816 ( 
.A(n_746),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_735),
.B(n_721),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_747),
.A2(n_715),
.B(n_691),
.C(n_695),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_733),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_775),
.B(n_652),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_743),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_784),
.Y(n_822)
);

AO31x2_ASAP7_75t_L g823 ( 
.A1(n_759),
.A2(n_644),
.A3(n_708),
.B(n_727),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_737),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_745),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_744),
.A2(n_678),
.B(n_707),
.Y(n_826)
);

AO31x2_ASAP7_75t_L g827 ( 
.A1(n_804),
.A2(n_722),
.A3(n_719),
.B(n_723),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_749),
.A2(n_703),
.B1(n_714),
.B2(n_731),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_757),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_775),
.B(n_681),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_765),
.A2(n_753),
.B(n_763),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_772),
.B(n_670),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_750),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_778),
.B(n_692),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_785),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_765),
.A2(n_697),
.B(n_647),
.Y(n_836)
);

AO22x2_ASAP7_75t_L g837 ( 
.A1(n_751),
.A2(n_697),
.B1(n_654),
.B2(n_666),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_748),
.A2(n_672),
.B1(n_654),
.B2(n_666),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_767),
.A2(n_699),
.B(n_700),
.C(n_731),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_752),
.A2(n_702),
.B(n_704),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_800),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_788),
.A2(n_448),
.B1(n_12),
.B2(n_13),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_777),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_797),
.A2(n_635),
.B(n_12),
.C(n_13),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_SL g845 ( 
.A1(n_805),
.A2(n_11),
.B(n_14),
.C(n_15),
.Y(n_845)
);

AO31x2_ASAP7_75t_L g846 ( 
.A1(n_804),
.A2(n_11),
.A3(n_14),
.B(n_15),
.Y(n_846)
);

AOI221x1_ASAP7_75t_L g847 ( 
.A1(n_782),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.C(n_22),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_761),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_788),
.B(n_19),
.Y(n_849)
);

NAND2x1p5_ASAP7_75t_L g850 ( 
.A(n_800),
.B(n_67),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_773),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_789),
.B(n_20),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_789),
.B(n_22),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_781),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_760),
.A2(n_113),
.B(n_181),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_SL g856 ( 
.A1(n_774),
.A2(n_23),
.B(n_24),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_SL g857 ( 
.A(n_778),
.B(n_23),
.C(n_24),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_780),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_801),
.A2(n_448),
.B(n_115),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_801),
.A2(n_448),
.B(n_109),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_776),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_760),
.A2(n_117),
.B(n_177),
.Y(n_862)
);

AOI211x1_ASAP7_75t_L g863 ( 
.A1(n_798),
.A2(n_25),
.B(n_26),
.C(n_28),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_SL g864 ( 
.A1(n_776),
.A2(n_106),
.B(n_176),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_802),
.A2(n_25),
.B(n_26),
.C(n_29),
.Y(n_865)
);

INVx3_ASAP7_75t_SL g866 ( 
.A(n_779),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_800),
.A2(n_799),
.B(n_798),
.Y(n_867)
);

NAND3xp33_ASAP7_75t_L g868 ( 
.A(n_799),
.B(n_29),
.C(n_30),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_821),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_837),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_814),
.A2(n_740),
.B1(n_779),
.B2(n_792),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_809),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_814),
.A2(n_771),
.B1(n_755),
.B2(n_800),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_837),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_854),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_837),
.Y(n_876)
);

BUFx12f_ASAP7_75t_L g877 ( 
.A(n_816),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_825),
.Y(n_878)
);

INVx6_ASAP7_75t_L g879 ( 
.A(n_851),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_846),
.Y(n_880)
);

CKINVDCx11_ASAP7_75t_R g881 ( 
.A(n_810),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_841),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_857),
.A2(n_793),
.B1(n_803),
.B2(n_782),
.Y(n_883)
);

INVx6_ASAP7_75t_L g884 ( 
.A(n_824),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_819),
.B(n_734),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_846),
.Y(n_886)
);

INVx4_ASAP7_75t_SL g887 ( 
.A(n_846),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_835),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_857),
.A2(n_793),
.B1(n_754),
.B2(n_784),
.Y(n_889)
);

BUFx12f_ASAP7_75t_L g890 ( 
.A(n_829),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_819),
.B(n_732),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_858),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_861),
.A2(n_736),
.B1(n_770),
.B2(n_787),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_822),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_811),
.A2(n_736),
.B1(n_770),
.B2(n_791),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_807),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_832),
.B(n_756),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_822),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_846),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_808),
.A2(n_796),
.B1(n_769),
.B2(n_756),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_841),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_823),
.Y(n_902)
);

CKINVDCx14_ASAP7_75t_R g903 ( 
.A(n_833),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_843),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_806),
.B(n_768),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_868),
.A2(n_783),
.B1(n_796),
.B2(n_769),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_849),
.A2(n_796),
.B1(n_769),
.B2(n_756),
.Y(n_907)
);

INVx6_ASAP7_75t_L g908 ( 
.A(n_834),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_823),
.Y(n_909)
);

BUFx12f_ASAP7_75t_L g910 ( 
.A(n_850),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_852),
.A2(n_448),
.B1(n_758),
.B2(n_33),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_866),
.Y(n_912)
);

CKINVDCx11_ASAP7_75t_R g913 ( 
.A(n_866),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_817),
.Y(n_914)
);

CKINVDCx6p67_ASAP7_75t_R g915 ( 
.A(n_848),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_850),
.Y(n_916)
);

BUFx10_ASAP7_75t_L g917 ( 
.A(n_864),
.Y(n_917)
);

INVx5_ASAP7_75t_L g918 ( 
.A(n_818),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_SL g919 ( 
.A1(n_853),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_818),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_842),
.A2(n_813),
.B1(n_820),
.B2(n_830),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_812),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_838),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_828),
.A2(n_758),
.B1(n_35),
.B2(n_36),
.Y(n_924)
);

INVx5_ASAP7_75t_L g925 ( 
.A(n_855),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_856),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_823),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_867),
.Y(n_928)
);

CKINVDCx6p67_ASAP7_75t_R g929 ( 
.A(n_847),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_827),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_SL g931 ( 
.A1(n_926),
.A2(n_842),
.B(n_865),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_880),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_896),
.Y(n_933)
);

NOR2x1_ASAP7_75t_SL g934 ( 
.A(n_918),
.B(n_826),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_880),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_882),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_886),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_896),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_918),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_886),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_928),
.Y(n_941)
);

OR2x6_ASAP7_75t_L g942 ( 
.A(n_905),
.B(n_815),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_928),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_899),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_905),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_899),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_927),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_927),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_887),
.Y(n_949)
);

CKINVDCx16_ASAP7_75t_R g950 ( 
.A(n_890),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_L g951 ( 
.A1(n_926),
.A2(n_859),
.B1(n_860),
.B2(n_862),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_870),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_870),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_902),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_923),
.B(n_865),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_902),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_874),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_930),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_918),
.Y(n_959)
);

AO21x2_ASAP7_75t_L g960 ( 
.A1(n_874),
.A2(n_831),
.B(n_844),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_908),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_876),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_905),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_909),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_918),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_909),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_876),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_930),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_887),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_887),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_931),
.A2(n_918),
.B(n_844),
.C(n_923),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_955),
.A2(n_918),
.B1(n_929),
.B2(n_920),
.Y(n_972)
);

OA21x2_ASAP7_75t_L g973 ( 
.A1(n_935),
.A2(n_906),
.B(n_883),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_931),
.A2(n_921),
.B(n_925),
.C(n_919),
.Y(n_974)
);

AOI221xp5_ASAP7_75t_L g975 ( 
.A1(n_955),
.A2(n_845),
.B1(n_863),
.B2(n_872),
.C(n_924),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_941),
.B(n_872),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_SL g977 ( 
.A1(n_941),
.A2(n_914),
.B(n_871),
.C(n_922),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_951),
.A2(n_925),
.B(n_840),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_961),
.Y(n_979)
);

AOI221xp5_ASAP7_75t_L g980 ( 
.A1(n_951),
.A2(n_845),
.B1(n_885),
.B2(n_911),
.C(n_875),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_961),
.B(n_882),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_961),
.B(n_897),
.Y(n_982)
);

OAI21x1_ASAP7_75t_SL g983 ( 
.A1(n_934),
.A2(n_869),
.B(n_873),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_SL g984 ( 
.A1(n_939),
.A2(n_965),
.B(n_959),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_943),
.B(n_875),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_943),
.B(n_908),
.Y(n_986)
);

AO32x2_ASAP7_75t_L g987 ( 
.A1(n_933),
.A2(n_900),
.A3(n_929),
.B1(n_887),
.B2(n_895),
.Y(n_987)
);

NOR2x1_ASAP7_75t_SL g988 ( 
.A(n_939),
.B(n_910),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_936),
.B(n_908),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_939),
.A2(n_965),
.B(n_959),
.C(n_925),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_936),
.B(n_908),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_969),
.B(n_962),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_952),
.B(n_869),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_942),
.A2(n_889),
.B(n_925),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_939),
.A2(n_925),
.B(n_916),
.C(n_839),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_958),
.B(n_897),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_952),
.B(n_878),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_942),
.A2(n_925),
.B(n_907),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_953),
.B(n_878),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_953),
.B(n_888),
.Y(n_1000)
);

AO32x2_ASAP7_75t_L g1001 ( 
.A1(n_933),
.A2(n_893),
.A3(n_920),
.B1(n_758),
.B2(n_901),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_958),
.B(n_901),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_969),
.B(n_912),
.Y(n_1003)
);

AOI221xp5_ASAP7_75t_L g1004 ( 
.A1(n_960),
.A2(n_891),
.B1(n_888),
.B2(n_828),
.C(n_892),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_958),
.B(n_957),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_962),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_957),
.B(n_892),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_962),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_939),
.A2(n_884),
.B1(n_915),
.B2(n_879),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_967),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_967),
.B(n_920),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_950),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_934),
.B(n_920),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_992),
.B(n_934),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_1006),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_1003),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_992),
.B(n_968),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_987),
.B(n_968),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1008),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_1005),
.B(n_935),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_980),
.A2(n_960),
.B1(n_965),
.B2(n_959),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_1010),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_974),
.A2(n_960),
.B1(n_939),
.B2(n_959),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_985),
.B(n_935),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_997),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_993),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_999),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_987),
.B(n_968),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_1000),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_987),
.B(n_968),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_976),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_987),
.B(n_946),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_1001),
.B(n_946),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_980),
.A2(n_960),
.B1(n_959),
.B2(n_939),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_990),
.B(n_969),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1007),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1001),
.B(n_946),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_986),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1004),
.B(n_932),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1001),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1018),
.B(n_1013),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_1015),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1029),
.B(n_1004),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_1035),
.B(n_984),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_1032),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_1035),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1018),
.B(n_1002),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1032),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1032),
.Y(n_1049)
);

OAI33xp33_ASAP7_75t_L g1050 ( 
.A1(n_1039),
.A2(n_991),
.A3(n_989),
.B1(n_937),
.B2(n_940),
.B3(n_944),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1018),
.B(n_996),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_1014),
.B(n_969),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1033),
.Y(n_1053)
);

AOI33xp33_ASAP7_75t_L g1054 ( 
.A1(n_1021),
.A2(n_972),
.A3(n_977),
.B1(n_975),
.B2(n_1012),
.B3(n_1011),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_1040),
.B(n_932),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1028),
.B(n_1001),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_1014),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1015),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1022),
.Y(n_1059)
);

AOI221x1_ASAP7_75t_SL g1060 ( 
.A1(n_1040),
.A2(n_1009),
.B1(n_41),
.B2(n_42),
.C(n_43),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_1035),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1022),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1055),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1053),
.B(n_1028),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1046),
.B(n_1014),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1055),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_1054),
.B(n_1038),
.Y(n_1067)
);

INVxp67_ASAP7_75t_L g1068 ( 
.A(n_1042),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1055),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1046),
.B(n_1028),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1046),
.B(n_1030),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1046),
.B(n_1030),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1059),
.B(n_1031),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1042),
.Y(n_1074)
);

OAI22xp33_ASAP7_75t_SL g1075 ( 
.A1(n_1067),
.A2(n_1044),
.B1(n_1061),
.B2(n_1057),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_1068),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1065),
.B(n_1052),
.Y(n_1077)
);

AND2x4_ASAP7_75t_SL g1078 ( 
.A(n_1065),
.B(n_1044),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1068),
.B(n_1074),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1074),
.B(n_1056),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1070),
.B(n_1052),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_1070),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1078),
.B(n_1061),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1076),
.B(n_1073),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1082),
.Y(n_1085)
);

OAI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1080),
.A2(n_1023),
.B1(n_1044),
.B2(n_1061),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1077),
.B(n_1061),
.Y(n_1087)
);

OAI33xp33_ASAP7_75t_L g1088 ( 
.A1(n_1084),
.A2(n_1079),
.A3(n_1075),
.B1(n_1086),
.B2(n_1085),
.B3(n_1080),
.Y(n_1088)
);

OR2x2_ASAP7_75t_L g1089 ( 
.A(n_1084),
.B(n_1079),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_1083),
.A2(n_974),
.B(n_977),
.C(n_971),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_1087),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1085),
.B(n_1073),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_1086),
.B(n_1054),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1086),
.A2(n_1043),
.B(n_1044),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1085),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1085),
.B(n_1071),
.Y(n_1096)
);

XNOR2x1_ASAP7_75t_L g1097 ( 
.A(n_1086),
.B(n_904),
.Y(n_1097)
);

AOI322xp5_ASAP7_75t_L g1098 ( 
.A1(n_1086),
.A2(n_1056),
.A3(n_1072),
.B1(n_1071),
.B2(n_1064),
.C1(n_1040),
.C2(n_1048),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1084),
.B(n_1066),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1091),
.B(n_1081),
.Y(n_1100)
);

AOI221x1_ASAP7_75t_L g1101 ( 
.A1(n_1095),
.A2(n_1061),
.B1(n_1059),
.B2(n_1062),
.C(n_1058),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1093),
.A2(n_1044),
.B1(n_1061),
.B2(n_1023),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1089),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1092),
.Y(n_1104)
);

OAI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1088),
.A2(n_1044),
.B1(n_1060),
.B2(n_1043),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1097),
.A2(n_978),
.B(n_1021),
.Y(n_1106)
);

OAI32xp33_ASAP7_75t_L g1107 ( 
.A1(n_1096),
.A2(n_1040),
.A3(n_1060),
.B1(n_1056),
.B2(n_1045),
.Y(n_1107)
);

OAI221xp5_ASAP7_75t_L g1108 ( 
.A1(n_1094),
.A2(n_1098),
.B1(n_1099),
.B2(n_1090),
.C(n_1034),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1099),
.B(n_1072),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1092),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1095),
.Y(n_1111)
);

NAND2x1_ASAP7_75t_L g1112 ( 
.A(n_1095),
.B(n_1044),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1093),
.A2(n_978),
.B(n_1034),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1093),
.A2(n_972),
.B(n_995),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1092),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1103),
.B(n_1066),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_1103),
.Y(n_1117)
);

NAND2x1_ASAP7_75t_SL g1118 ( 
.A(n_1103),
.B(n_1064),
.Y(n_1118)
);

XOR2x2_ASAP7_75t_L g1119 ( 
.A(n_1114),
.B(n_950),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1111),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1111),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1100),
.Y(n_1122)
);

AOI222xp33_ASAP7_75t_L g1123 ( 
.A1(n_1105),
.A2(n_1050),
.B1(n_975),
.B2(n_994),
.C1(n_1039),
.C2(n_1064),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1105),
.B(n_877),
.Y(n_1124)
);

INVxp67_ASAP7_75t_SL g1125 ( 
.A(n_1113),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1100),
.Y(n_1126)
);

OAI222xp33_ASAP7_75t_L g1127 ( 
.A1(n_1108),
.A2(n_1057),
.B1(n_1069),
.B2(n_1063),
.C1(n_1035),
.C2(n_1062),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1104),
.B(n_1069),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_1106),
.B(n_877),
.Y(n_1129)
);

AOI222xp33_ASAP7_75t_L g1130 ( 
.A1(n_1107),
.A2(n_1050),
.B1(n_1030),
.B2(n_890),
.C1(n_1049),
.C2(n_1045),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1109),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1109),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1110),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1115),
.B(n_1041),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_1117),
.B(n_1102),
.Y(n_1135)
);

NOR3xp33_ASAP7_75t_L g1136 ( 
.A(n_1124),
.B(n_1112),
.C(n_881),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1122),
.B(n_904),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_1126),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1131),
.B(n_1101),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1133),
.B(n_903),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1124),
.A2(n_1038),
.B(n_1063),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1131),
.B(n_1063),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1132),
.B(n_1057),
.Y(n_1143)
);

AOI211xp5_ASAP7_75t_L g1144 ( 
.A1(n_1125),
.A2(n_1127),
.B(n_1129),
.C(n_1120),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1118),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1125),
.B(n_879),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1121),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1119),
.B(n_1057),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1123),
.B(n_1041),
.Y(n_1149)
);

NAND3xp33_ASAP7_75t_SL g1150 ( 
.A(n_1129),
.B(n_1130),
.C(n_1116),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1128),
.Y(n_1151)
);

AOI221xp5_ASAP7_75t_L g1152 ( 
.A1(n_1144),
.A2(n_1134),
.B1(n_1062),
.B2(n_1059),
.C(n_1058),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_SL g1153 ( 
.A1(n_1136),
.A2(n_1035),
.B(n_998),
.Y(n_1153)
);

OAI221xp5_ASAP7_75t_L g1154 ( 
.A1(n_1141),
.A2(n_884),
.B1(n_879),
.B2(n_1031),
.C(n_1058),
.Y(n_1154)
);

OAI221xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1145),
.A2(n_915),
.B1(n_1049),
.B2(n_1048),
.C(n_1045),
.Y(n_1155)
);

AOI32xp33_ASAP7_75t_L g1156 ( 
.A1(n_1148),
.A2(n_1035),
.A3(n_1041),
.B1(n_1048),
.B2(n_1049),
.Y(n_1156)
);

NAND4xp25_ASAP7_75t_L g1157 ( 
.A(n_1135),
.B(n_913),
.C(n_916),
.D(n_884),
.Y(n_1157)
);

NAND2xp33_ASAP7_75t_R g1158 ( 
.A(n_1146),
.B(n_1137),
.Y(n_1158)
);

AOI211xp5_ASAP7_75t_SL g1159 ( 
.A1(n_1138),
.A2(n_884),
.B(n_879),
.C(n_43),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1140),
.A2(n_1052),
.B1(n_1049),
.B2(n_1048),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1139),
.A2(n_1045),
.B(n_1053),
.C(n_1037),
.Y(n_1161)
);

OA211x2_ASAP7_75t_L g1162 ( 
.A1(n_1150),
.A2(n_39),
.B(n_41),
.C(n_44),
.Y(n_1162)
);

NAND4xp25_ASAP7_75t_L g1163 ( 
.A(n_1150),
.B(n_1016),
.C(n_922),
.D(n_1052),
.Y(n_1163)
);

OAI221xp5_ASAP7_75t_L g1164 ( 
.A1(n_1149),
.A2(n_1053),
.B1(n_912),
.B2(n_1036),
.C(n_1027),
.Y(n_1164)
);

AND4x1_ASAP7_75t_L g1165 ( 
.A(n_1147),
.B(n_44),
.C(n_45),
.D(n_47),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1151),
.B(n_1053),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_1142),
.Y(n_1167)
);

OAI211xp5_ASAP7_75t_L g1168 ( 
.A1(n_1143),
.A2(n_912),
.B(n_48),
.C(n_49),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1138),
.B(n_1047),
.Y(n_1169)
);

AOI221xp5_ASAP7_75t_L g1170 ( 
.A1(n_1144),
.A2(n_1033),
.B1(n_1037),
.B2(n_1036),
.C(n_1027),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1138),
.B(n_1047),
.Y(n_1171)
);

OAI21xp33_ASAP7_75t_L g1172 ( 
.A1(n_1149),
.A2(n_1052),
.B(n_1003),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1144),
.A2(n_1052),
.B1(n_1016),
.B2(n_1047),
.Y(n_1173)
);

AOI221xp5_ASAP7_75t_L g1174 ( 
.A1(n_1144),
.A2(n_1037),
.B1(n_1033),
.B2(n_983),
.C(n_960),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1138),
.B(n_1051),
.Y(n_1175)
);

NOR3xp33_ASAP7_75t_L g1176 ( 
.A(n_1157),
.B(n_1016),
.C(n_49),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1152),
.A2(n_1051),
.B(n_1029),
.C(n_51),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1173),
.A2(n_910),
.B1(n_912),
.B2(n_1016),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1162),
.A2(n_912),
.B1(n_1016),
.B2(n_1051),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1170),
.B(n_1029),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1165),
.Y(n_1181)
);

NAND4xp25_ASAP7_75t_L g1182 ( 
.A(n_1158),
.B(n_979),
.C(n_982),
.D(n_52),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1159),
.A2(n_894),
.B(n_1029),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1168),
.A2(n_988),
.B(n_942),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_1167),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1169),
.Y(n_1186)
);

NAND4xp25_ASAP7_75t_L g1187 ( 
.A(n_1163),
.B(n_47),
.C(n_50),
.D(n_53),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_SL g1188 ( 
.A1(n_1174),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.C(n_56),
.Y(n_1188)
);

NAND4xp25_ASAP7_75t_L g1189 ( 
.A(n_1171),
.B(n_55),
.C(n_57),
.D(n_981),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_SL g1190 ( 
.A(n_1155),
.B(n_917),
.Y(n_1190)
);

AOI221xp5_ASAP7_75t_SL g1191 ( 
.A1(n_1154),
.A2(n_1019),
.B1(n_970),
.B2(n_1025),
.C(n_939),
.Y(n_1191)
);

AOI211xp5_ASAP7_75t_L g1192 ( 
.A1(n_1153),
.A2(n_1164),
.B(n_1175),
.C(n_1166),
.Y(n_1192)
);

AOI21xp33_ASAP7_75t_SL g1193 ( 
.A1(n_1161),
.A2(n_68),
.B(n_69),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1172),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1156),
.A2(n_949),
.B(n_973),
.C(n_942),
.Y(n_1195)
);

OAI211xp5_ASAP7_75t_SL g1196 ( 
.A1(n_1160),
.A2(n_898),
.B(n_970),
.C(n_1024),
.Y(n_1196)
);

OAI211xp5_ASAP7_75t_SL g1197 ( 
.A1(n_1152),
.A2(n_898),
.B(n_970),
.C(n_1024),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1152),
.A2(n_1024),
.B(n_1025),
.Y(n_1198)
);

NAND4xp25_ASAP7_75t_SL g1199 ( 
.A(n_1152),
.B(n_1020),
.C(n_1017),
.D(n_1025),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1185),
.Y(n_1200)
);

XNOR2x1_ASAP7_75t_L g1201 ( 
.A(n_1181),
.B(n_71),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1194),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1186),
.Y(n_1203)
);

NOR2x1_ASAP7_75t_L g1204 ( 
.A(n_1189),
.B(n_1019),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1182),
.B(n_1187),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1192),
.Y(n_1206)
);

NAND2x1p5_ASAP7_75t_L g1207 ( 
.A(n_1179),
.B(n_959),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1176),
.Y(n_1208)
);

NOR2x1_ASAP7_75t_L g1209 ( 
.A(n_1177),
.B(n_898),
.Y(n_1209)
);

NAND3x1_ASAP7_75t_L g1210 ( 
.A(n_1178),
.B(n_1017),
.C(n_963),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1180),
.Y(n_1211)
);

INVxp33_ASAP7_75t_SL g1212 ( 
.A(n_1190),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1193),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1183),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1188),
.B(n_1025),
.Y(n_1215)
);

NAND4xp75_ASAP7_75t_L g1216 ( 
.A(n_1191),
.B(n_973),
.C(n_1017),
.D(n_836),
.Y(n_1216)
);

NAND2x1p5_ASAP7_75t_L g1217 ( 
.A(n_1184),
.B(n_959),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1199),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1198),
.B(n_1197),
.Y(n_1219)
);

NAND4xp75_ASAP7_75t_L g1220 ( 
.A(n_1195),
.B(n_944),
.C(n_940),
.D(n_937),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1196),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1212),
.A2(n_981),
.B1(n_917),
.B2(n_965),
.Y(n_1222)
);

NOR2x1p5_ASAP7_75t_L g1223 ( 
.A(n_1202),
.B(n_1208),
.Y(n_1223)
);

NOR2x1_ASAP7_75t_L g1224 ( 
.A(n_1200),
.B(n_84),
.Y(n_1224)
);

OAI221xp5_ASAP7_75t_L g1225 ( 
.A1(n_1218),
.A2(n_1206),
.B1(n_1213),
.B2(n_1217),
.C(n_1205),
.Y(n_1225)
);

NAND3xp33_ASAP7_75t_L g1226 ( 
.A(n_1203),
.B(n_1026),
.C(n_959),
.Y(n_1226)
);

AND4x1_ASAP7_75t_L g1227 ( 
.A(n_1214),
.B(n_93),
.C(n_95),
.D(n_104),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1218),
.B(n_1026),
.Y(n_1228)
);

NAND3xp33_ASAP7_75t_L g1229 ( 
.A(n_1214),
.B(n_1026),
.C(n_965),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1201),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_SL g1231 ( 
.A(n_1211),
.B(n_1026),
.C(n_1020),
.Y(n_1231)
);

OAI21xp33_ASAP7_75t_L g1232 ( 
.A1(n_1215),
.A2(n_1020),
.B(n_949),
.Y(n_1232)
);

NAND3x1_ASAP7_75t_L g1233 ( 
.A(n_1209),
.B(n_963),
.C(n_945),
.Y(n_1233)
);

AOI22x1_ASAP7_75t_L g1234 ( 
.A1(n_1207),
.A2(n_965),
.B1(n_118),
.B2(n_119),
.Y(n_1234)
);

AOI221xp5_ASAP7_75t_L g1235 ( 
.A1(n_1221),
.A2(n_965),
.B1(n_963),
.B2(n_945),
.C(n_947),
.Y(n_1235)
);

AOI221xp5_ASAP7_75t_L g1236 ( 
.A1(n_1219),
.A2(n_965),
.B1(n_963),
.B2(n_945),
.C(n_947),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1224),
.B(n_1204),
.Y(n_1237)
);

CKINVDCx14_ASAP7_75t_R g1238 ( 
.A(n_1230),
.Y(n_1238)
);

OAI21xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1223),
.A2(n_1220),
.B(n_1216),
.Y(n_1239)
);

AND3x1_ASAP7_75t_L g1240 ( 
.A(n_1228),
.B(n_1219),
.C(n_1210),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1227),
.B(n_963),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1225),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1232),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1231),
.A2(n_917),
.B1(n_945),
.B2(n_942),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_SL g1245 ( 
.A1(n_1222),
.A2(n_917),
.B1(n_942),
.B2(n_947),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_1234),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1229),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1226),
.A2(n_945),
.B1(n_942),
.B2(n_933),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1233),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1236),
.B(n_105),
.Y(n_1250)
);

AND3x1_ASAP7_75t_L g1251 ( 
.A(n_1235),
.B(n_124),
.C(n_125),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1238),
.A2(n_948),
.B1(n_938),
.B2(n_956),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1246),
.A2(n_948),
.B1(n_938),
.B2(n_956),
.Y(n_1253)
);

AO22x2_ASAP7_75t_L g1254 ( 
.A1(n_1242),
.A2(n_938),
.B1(n_964),
.B2(n_956),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1237),
.A2(n_938),
.B1(n_964),
.B2(n_956),
.Y(n_1255)
);

INVxp67_ASAP7_75t_SL g1256 ( 
.A(n_1247),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1240),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1243),
.A2(n_966),
.B1(n_964),
.B2(n_954),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_SL g1259 ( 
.A1(n_1251),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_1259)
);

AOI22xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1249),
.A2(n_131),
.B1(n_136),
.B2(n_137),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1239),
.A2(n_966),
.B1(n_964),
.B2(n_954),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1257),
.A2(n_1244),
.B1(n_1241),
.B2(n_1250),
.Y(n_1262)
);

XNOR2x1_ASAP7_75t_L g1263 ( 
.A(n_1256),
.B(n_1248),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1260),
.A2(n_1245),
.B(n_141),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1254),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1259),
.Y(n_1266)
);

NOR4xp75_ASAP7_75t_L g1267 ( 
.A(n_1258),
.B(n_139),
.C(n_142),
.D(n_145),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1266),
.A2(n_1261),
.B1(n_1252),
.B2(n_1253),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1263),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1264),
.A2(n_1255),
.B(n_147),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1267),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1270),
.A2(n_1262),
.B(n_1265),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1272),
.A2(n_1269),
.B(n_1271),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1273),
.A2(n_1268),
.B(n_149),
.Y(n_1274)
);

OAI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1274),
.A2(n_146),
.B1(n_150),
.B2(n_153),
.Y(n_1275)
);

AOI221xp5_ASAP7_75t_L g1276 ( 
.A1(n_1275),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.C(n_161),
.Y(n_1276)
);

AOI211xp5_ASAP7_75t_L g1277 ( 
.A1(n_1276),
.A2(n_163),
.B(n_165),
.C(n_167),
.Y(n_1277)
);


endmodule