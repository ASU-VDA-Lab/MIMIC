module fake_jpeg_29145_n_181 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_181);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_80),
.Y(n_94)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_85),
.Y(n_96)
);

INVx11_ASAP7_75t_SL g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_65),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_91),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_72),
.B1(n_68),
.B2(n_55),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_98),
.B1(n_99),
.B2(n_71),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_55),
.B1(n_60),
.B2(n_66),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_95),
.Y(n_103)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_76),
.C(n_75),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_68),
.B1(n_72),
.B2(n_61),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_72),
.B1(n_57),
.B2(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_63),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_108),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_73),
.B(n_51),
.C(n_70),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_103),
.C(n_116),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_52),
.B1(n_69),
.B2(n_62),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_120),
.B1(n_1),
.B2(n_2),
.Y(n_126)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_95),
.B(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_111),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_56),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_116),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_54),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_14),
.Y(n_123)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_53),
.B1(n_27),
.B2(n_28),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_0),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_49),
.B1(n_17),
.B2(n_30),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_128),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_114),
.A2(n_109),
.B1(n_115),
.B2(n_103),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_139),
.B1(n_121),
.B2(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_127),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_32),
.C(n_45),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_10),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_3),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_102),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_12),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_144)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_4),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_141),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_6),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_147),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_158),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_10),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_11),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_157),
.B(n_36),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_12),
.B1(n_13),
.B2(n_34),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_151),
.A2(n_38),
.B(n_39),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_134),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_130),
.B1(n_136),
.B2(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_156),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_13),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_35),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_42),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g168 ( 
.A(n_163),
.B(n_155),
.CI(n_158),
.CON(n_168),
.SN(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_145),
.B1(n_143),
.B2(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_162),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_142),
.B(n_161),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_172),
.B(n_171),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_171),
.C(n_168),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_167),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_165),
.B(n_170),
.Y(n_179)
);

OAI221xp5_ASAP7_75t_SL g180 ( 
.A1(n_179),
.A2(n_168),
.B1(n_166),
.B2(n_164),
.C(n_154),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_163),
.Y(n_181)
);


endmodule