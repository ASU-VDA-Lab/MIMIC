module fake_aes_2304_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
CKINVDCx5p33_ASAP7_75t_R g3 ( .A(n_1), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
INVx2_ASAP7_75t_SL g5 ( .A(n_2), .Y(n_5) );
BUFx6f_ASAP7_75t_L g6 ( .A(n_5), .Y(n_6) );
OAI22xp33_ASAP7_75t_L g7 ( .A1(n_3), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_8), .B(n_3), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
NAND2x1p5_ASAP7_75t_L g12 ( .A(n_10), .B(n_4), .Y(n_12) );
A2O1A1Ixp33_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_5), .B(n_4), .C(n_6), .Y(n_13) );
AOI22xp5_ASAP7_75t_L g14 ( .A1(n_12), .A2(n_7), .B1(n_4), .B2(n_6), .Y(n_14) );
AOI22xp5_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_12), .B1(n_6), .B2(n_10), .Y(n_15) );
NAND4xp75_ASAP7_75t_L g16 ( .A(n_13), .B(n_0), .C(n_1), .D(n_6), .Y(n_16) );
AOI22xp5_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_0), .B1(n_1), .B2(n_15), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_0), .Y(n_18) );
endmodule