module fake_jpeg_14973_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_65),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_69)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_61),
.B1(n_57),
.B2(n_3),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_0),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_48),
.B1(n_55),
.B2(n_49),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_80),
.Y(n_87)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_56),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_78),
.B(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_54),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_60),
.B1(n_51),
.B2(n_52),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_60),
.B1(n_52),
.B2(n_51),
.Y(n_92)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_90),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_102),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_57),
.B1(n_62),
.B2(n_50),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_99),
.B1(n_76),
.B2(n_25),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_62),
.B(n_2),
.C(n_4),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_30),
.C(n_11),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_100),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_9),
.B(n_13),
.C(n_14),
.Y(n_99)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_104),
.B(n_113),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_105),
.A2(n_111),
.B1(n_97),
.B2(n_112),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_95),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_94),
.B1(n_101),
.B2(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_118),
.B(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_115),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_107),
.C(n_111),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_110),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_119),
.C(n_110),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_126),
.A2(n_127),
.B(n_129),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_117),
.B1(n_110),
.B2(n_116),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_29),
.C(n_31),
.Y(n_132)
);

XNOR2x1_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_124),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_130),
.B1(n_34),
.B2(n_35),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_135),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_33),
.C(n_36),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_37),
.C(n_38),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_39),
.C(n_40),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_42),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_44),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_93),
.Y(n_144)
);

BUFx24_ASAP7_75t_SL g145 ( 
.A(n_144),
.Y(n_145)
);


endmodule