module fake_jpeg_31656_n_373 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_373);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_373;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_56),
.Y(n_93)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_15),
.B(n_14),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_15),
.B(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_62),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_70),
.Y(n_113)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_69),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_12),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_76),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_74),
.Y(n_126)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_73),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_40),
.CON(n_92),
.SN(n_92)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_31),
.B(n_23),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_77),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_22),
.B(n_12),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_35),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_113),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g157 ( 
.A1(n_92),
.A2(n_128),
.B1(n_109),
.B2(n_130),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_18),
.B1(n_16),
.B2(n_27),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_95),
.A2(n_108),
.B1(n_120),
.B2(n_123),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_49),
.A2(n_18),
.B1(n_27),
.B2(n_22),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_97),
.A2(n_110),
.B1(n_116),
.B2(n_121),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_41),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_101),
.B(n_107),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_41),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_18),
.B1(n_27),
.B2(n_37),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_18),
.B1(n_27),
.B2(n_35),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_73),
.A2(n_37),
.B1(n_39),
.B2(n_28),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_57),
.A2(n_30),
.B1(n_17),
.B2(n_34),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_114),
.B1(n_124),
.B2(n_50),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_45),
.A2(n_30),
.B1(n_17),
.B2(n_34),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_39),
.B1(n_28),
.B2(n_21),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_44),
.B(n_21),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_119),
.C(n_9),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_55),
.A2(n_36),
.B1(n_38),
.B2(n_65),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_38),
.B1(n_36),
.B2(n_3),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_59),
.A2(n_38),
.B1(n_36),
.B2(n_3),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_61),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_129),
.B1(n_77),
.B2(n_42),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_60),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_74),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_68),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_127),
.A2(n_98),
.B1(n_118),
.B2(n_87),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_80),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_133),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_134),
.B(n_135),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_88),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_137),
.A2(n_165),
.B1(n_143),
.B2(n_136),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_53),
.B1(n_52),
.B2(n_67),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_144),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_48),
.B1(n_43),
.B2(n_62),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_146),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_43),
.B1(n_62),
.B2(n_9),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_92),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_9),
.B1(n_102),
.B2(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_145),
.A2(n_151),
.B1(n_153),
.B2(n_155),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_102),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_147),
.A2(n_85),
.B(n_115),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_105),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_154),
.Y(n_180)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_97),
.A2(n_110),
.B1(n_122),
.B2(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_89),
.A2(n_98),
.B1(n_100),
.B2(n_83),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_116),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_94),
.B1(n_87),
.B2(n_111),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_160),
.Y(n_186)
);

AO22x1_ASAP7_75t_L g214 ( 
.A1(n_157),
.A2(n_169),
.B1(n_171),
.B2(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_93),
.B(n_126),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_90),
.B(n_103),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_162),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_99),
.B(n_83),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_91),
.B(n_89),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_168),
.Y(n_196)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_91),
.B(n_115),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_85),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_172),
.Y(n_208)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_128),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_174),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_177),
.B(n_192),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_147),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_181),
.B(n_184),
.C(n_190),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_134),
.B(n_158),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_183),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_175),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_139),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_175),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g231 ( 
.A(n_187),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_172),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_189),
.B(n_200),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_150),
.C(n_152),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_137),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_199),
.A2(n_173),
.B1(n_174),
.B2(n_133),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_135),
.B(n_163),
.C(n_159),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g203 ( 
.A(n_170),
.B(n_171),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_132),
.C(n_141),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_204),
.B(n_207),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_136),
.B(n_165),
.Y(n_207)
);

AO22x1_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_187),
.B1(n_208),
.B2(n_200),
.Y(n_238)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_215),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_228),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_217),
.A2(n_220),
.B1(n_233),
.B2(n_198),
.Y(n_261)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_138),
.B1(n_149),
.B2(n_189),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_138),
.B1(n_192),
.B2(n_184),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_221),
.A2(n_236),
.B1(n_234),
.B2(n_231),
.Y(n_268)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_183),
.A2(n_138),
.B(n_180),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_226),
.A2(n_234),
.B(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_203),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_229),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_191),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_232),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_188),
.B(n_186),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_193),
.A2(n_190),
.B1(n_214),
.B2(n_182),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_193),
.A2(n_177),
.B(n_214),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_201),
.A2(n_202),
.B1(n_196),
.B2(n_181),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_238),
.Y(n_260)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_243),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_212),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_241),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_204),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_212),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_245),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_185),
.A2(n_179),
.B(n_209),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_219),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_256),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_185),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_238),
.B(n_223),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_206),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_225),
.C(n_243),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_261),
.A2(n_263),
.B1(n_267),
.B2(n_240),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_220),
.A2(n_213),
.B1(n_205),
.B2(n_197),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_224),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_205),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_268),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_197),
.C(n_235),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_272),
.C(n_222),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_217),
.A2(n_233),
.B1(n_235),
.B2(n_238),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_222),
.A2(n_221),
.B(n_218),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_269),
.B(n_237),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_227),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_280),
.C(n_285),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_278),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_261),
.B1(n_260),
.B2(n_251),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_283),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_249),
.A2(n_245),
.B(n_241),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_282),
.A2(n_286),
.B(n_263),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_252),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_215),
.C(n_229),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_252),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_293),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_253),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_294),
.Y(n_307)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_253),
.Y(n_290)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_247),
.C(n_268),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_292),
.C(n_297),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_269),
.C(n_272),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_248),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_248),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_254),
.Y(n_295)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_259),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_296),
.B(n_250),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_255),
.C(n_260),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_298),
.A2(n_313),
.B1(n_278),
.B2(n_282),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_249),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_312),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_265),
.C(n_254),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_305),
.B(n_285),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_293),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_294),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_283),
.A2(n_273),
.B1(n_259),
.B2(n_262),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_310),
.A2(n_286),
.B1(n_295),
.B2(n_290),
.Y(n_320)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_311),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_262),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_279),
.A2(n_270),
.B1(n_250),
.B2(n_274),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_314),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_297),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_330),
.C(n_331),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_318),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_321),
.Y(n_337)
);

NAND3xp33_ASAP7_75t_SL g321 ( 
.A(n_300),
.B(n_307),
.C(n_316),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_316),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_324),
.Y(n_340)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_323),
.A2(n_315),
.B1(n_308),
.B2(n_304),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_277),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_329),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_303),
.B(n_280),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_299),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_310),
.A2(n_276),
.B(n_287),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_332),
.A2(n_302),
.B(n_308),
.Y(n_342)
);

FAx1_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_309),
.CI(n_305),
.CON(n_334),
.SN(n_334)
);

AO21x1_ASAP7_75t_L g352 ( 
.A1(n_334),
.A2(n_342),
.B(n_343),
.Y(n_352)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_335),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_326),
.B(n_277),
.Y(n_336)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_336),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_299),
.C(n_327),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_284),
.C(n_328),
.Y(n_353)
);

OAI21xp33_ASAP7_75t_L g341 ( 
.A1(n_325),
.A2(n_314),
.B(n_302),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_332),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_319),
.A2(n_313),
.B(n_304),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_323),
.Y(n_345)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_345),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_317),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_350),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_338),
.A2(n_301),
.B(n_291),
.Y(n_349)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_349),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_329),
.C(n_327),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_351),
.B(n_353),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_348),
.B(n_338),
.Y(n_355)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_355),
.Y(n_362)
);

AOI21xp33_ASAP7_75t_L g357 ( 
.A1(n_352),
.A2(n_337),
.B(n_334),
.Y(n_357)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_357),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_352),
.A2(n_343),
.B(n_342),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_358),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_360),
.B(n_353),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_365),
.C(n_359),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_351),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_364),
.A2(n_358),
.B1(n_346),
.B2(n_356),
.Y(n_366)
);

AOI322xp5_ASAP7_75t_L g369 ( 
.A1(n_366),
.A2(n_367),
.A3(n_363),
.B1(n_334),
.B2(n_289),
.C1(n_345),
.C2(n_344),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_339),
.C(n_344),
.Y(n_368)
);

OAI21xp33_ASAP7_75t_L g370 ( 
.A1(n_368),
.A2(n_284),
.B(n_363),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_370),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_270),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_320),
.C(n_274),
.Y(n_373)
);


endmodule