module fake_jpeg_20854_n_237 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_8),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_18),
.Y(n_70)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_24),
.B1(n_21),
.B2(n_26),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_68),
.B1(n_71),
.B2(n_73),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_34),
.B1(n_21),
.B2(n_20),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_57),
.B1(n_2),
.B2(n_3),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_34),
.B1(n_19),
.B2(n_31),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_39),
.B1(n_48),
.B2(n_36),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_59),
.B1(n_47),
.B2(n_49),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_33),
.B(n_25),
.C(n_18),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g103 ( 
.A(n_61),
.B(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_32),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_21),
.B1(n_26),
.B2(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_29),
.B1(n_33),
.B2(n_20),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_29),
.B1(n_20),
.B2(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_25),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_47),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_36),
.A2(n_30),
.B1(n_31),
.B2(n_19),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_77),
.B1(n_72),
.B2(n_60),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_30),
.B1(n_23),
.B2(n_32),
.Y(n_77)
);

OR2x2_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_22),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_79),
.B(n_87),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_80),
.B(n_93),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_44),
.B1(n_25),
.B2(n_47),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_83),
.A2(n_85),
.B1(n_86),
.B2(n_94),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_90),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_18),
.B1(n_35),
.B2(n_32),
.Y(n_86)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_42),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_18),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_18),
.B1(n_35),
.B2(n_38),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_14),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_102),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_104),
.B1(n_107),
.B2(n_65),
.Y(n_128)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_64),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_41),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_58),
.A2(n_35),
.B1(n_42),
.B2(n_38),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_109),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_61),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_114),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_41),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_118),
.C(n_122),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_64),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_63),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_80),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_63),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_134),
.Y(n_137)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_107),
.B(n_101),
.C(n_95),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_51),
.B1(n_66),
.B2(n_60),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_100),
.B1(n_89),
.B2(n_91),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_74),
.C(n_51),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_136),
.B(n_148),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_139),
.B(n_142),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_82),
.B1(n_99),
.B2(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_110),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_92),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_147),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_106),
.B1(n_88),
.B2(n_74),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_102),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_116),
.B(n_16),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_150),
.B(n_116),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_128),
.C(n_130),
.Y(n_162)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_55),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_155),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_126),
.B(n_120),
.C(n_113),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_100),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_89),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_157),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_91),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_161),
.B(n_176),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_166),
.A2(n_178),
.B(n_146),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_125),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_177),
.Y(n_181)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_112),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_138),
.B(n_114),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_158),
.A2(n_114),
.B1(n_133),
.B2(n_111),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_145),
.B(n_158),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_183),
.B(n_193),
.Y(n_205)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

AO21x1_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_157),
.B(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_173),
.B1(n_144),
.B2(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_140),
.B1(n_137),
.B2(n_147),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_190),
.Y(n_195)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_186),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_177),
.C(n_159),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_188),
.C(n_161),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_137),
.C(n_153),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_150),
.B1(n_154),
.B2(n_112),
.Y(n_190)
);

AO221x1_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_143),
.B1(n_115),
.B2(n_129),
.C(n_120),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_183),
.A2(n_167),
.B(n_174),
.C(n_170),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_197),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_194),
.B(n_172),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_200),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_170),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_178),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_187),
.C(n_188),
.Y(n_207)
);

AOI321xp33_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_164),
.A3(n_169),
.B1(n_175),
.B2(n_166),
.C(n_119),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_182),
.B(n_192),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_209),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_210),
.B1(n_204),
.B2(n_205),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_184),
.C(n_179),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_189),
.B1(n_191),
.B2(n_186),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_143),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_211),
.B(n_214),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_205),
.A2(n_191),
.B1(n_180),
.B2(n_193),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_216),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_115),
.C(n_16),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_198),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_203),
.Y(n_219)
);

AOI31xp33_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_196),
.A3(n_206),
.B(n_201),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_207),
.B(n_213),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_14),
.B1(n_4),
.B2(n_5),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_222),
.B(n_6),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_225),
.Y(n_231)
);

OAI221xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_213),
.B1(n_6),
.B2(n_7),
.C(n_10),
.Y(n_225)
);

AOI31xp33_ASAP7_75t_L g226 ( 
.A1(n_221),
.A2(n_2),
.A3(n_6),
.B(n_7),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_10),
.C(n_11),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_217),
.C(n_223),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_228),
.A2(n_217),
.B(n_10),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_230),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_231),
.C(n_232),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_236),
.Y(n_237)
);

AO21x1_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_11),
.B(n_230),
.Y(n_236)
);


endmodule