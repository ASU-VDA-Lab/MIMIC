module fake_aes_808_n_30 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_30);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_7;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g7 ( .A(n_6), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_4), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_5), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_1), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_4), .Y(n_11) );
O2A1O1Ixp33_ASAP7_75t_L g12 ( .A1(n_7), .A2(n_0), .B(n_1), .C(n_2), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_7), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
OAI22xp5_ASAP7_75t_L g15 ( .A1(n_11), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_16), .B(n_10), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_19), .B(n_16), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_17), .B(n_13), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
AOI221xp5_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_15), .B1(n_12), .B2(n_18), .C(n_9), .Y(n_24) );
NOR4xp75_ASAP7_75t_L g25 ( .A(n_23), .B(n_15), .C(n_12), .D(n_3), .Y(n_25) );
CKINVDCx20_ASAP7_75t_R g26 ( .A(n_25), .Y(n_26) );
AOI211xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_22), .B(n_2), .C(n_3), .Y(n_27) );
OAI22x1_ASAP7_75t_SL g28 ( .A1(n_26), .A2(n_0), .B1(n_3), .B2(n_4), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_5), .B1(n_6), .B2(n_0), .Y(n_29) );
AOI22xp33_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_5), .B1(n_6), .B2(n_28), .Y(n_30) );
endmodule