module fake_jpeg_3536_n_216 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_216);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_14),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_77),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_54),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx2_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

CKINVDCx12_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_66),
.B(n_63),
.C(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_69),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_60),
.B1(n_63),
.B2(n_75),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_95),
.B1(n_56),
.B2(n_68),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_72),
.Y(n_117)
);

CKINVDCx12_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_75),
.B1(n_56),
.B2(n_65),
.Y(n_95)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_64),
.Y(n_118)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_113),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_108),
.B1(n_112),
.B2(n_62),
.Y(n_125)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

OR2x2_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_109),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_68),
.B1(n_78),
.B2(n_64),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_98),
.A2(n_52),
.B1(n_73),
.B2(n_59),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_62),
.B1(n_71),
.B2(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_117),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_72),
.B1(n_52),
.B2(n_62),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_53),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_72),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_115),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_85),
.A2(n_67),
.B(n_74),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_97),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_51),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_0),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_24),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_114),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_150)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_71),
.B1(n_2),
.B2(n_3),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_135),
.B1(n_114),
.B2(n_5),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx6_ASAP7_75t_SL g145 ( 
.A(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_105),
.B1(n_107),
.B2(n_115),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_142),
.A2(n_161),
.B1(n_162),
.B2(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_148),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_150),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_4),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_149),
.B(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_6),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_152),
.Y(n_167)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_26),
.C(n_46),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_161),
.C(n_162),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_158),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_9),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_10),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_160),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_27),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_30),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_128),
.B(n_124),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_171),
.B(n_178),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_168),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_128),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_37),
.C(n_44),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_135),
.B(n_13),
.Y(n_171)
);

AO22x1_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_11),
.B1(n_15),
.B2(n_16),
.Y(n_173)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_16),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_21),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_150),
.B(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_140),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_181),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_191),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_19),
.B(n_20),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_189),
.C(n_177),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_40),
.C(n_45),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_164),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_196),
.C(n_165),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_181),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_174),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_198),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_182),
.B1(n_171),
.B2(n_175),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_188),
.A2(n_175),
.B(n_178),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_188),
.B(n_163),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_193),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_200),
.B(n_201),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_203),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_169),
.C(n_172),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_206),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_205),
.C(n_194),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_210),
.B(n_211),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_197),
.A3(n_190),
.B1(n_186),
.B2(n_184),
.C1(n_167),
.C2(n_173),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_212),
.B(n_208),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_208),
.A3(n_173),
.B1(n_35),
.B2(n_36),
.C1(n_42),
.C2(n_43),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_49),
.C(n_21),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_22),
.C(n_165),
.Y(n_216)
);


endmodule