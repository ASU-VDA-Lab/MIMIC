module fake_jpeg_15528_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_4),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_13),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_0),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_6),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_15),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_6),
.A2(n_1),
.B(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_19),
.C(n_21),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_7),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_24),
.B(n_10),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_14),
.B(n_8),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_9),
.B(n_12),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_9),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_23),
.C(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_5),
.B(n_11),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_30),
.B(n_34),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_30),
.Y(n_36)
);


endmodule