module fake_jpeg_18970_n_309 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_22),
.B(n_10),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_42),
.B(n_44),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_22),
.B(n_9),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_16),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_45),
.B(n_47),
.Y(n_113)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_64),
.Y(n_70)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g92 ( 
.A(n_60),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_62),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_29),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_29),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_69),
.B(n_74),
.Y(n_123)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_100),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_79),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_82),
.B(n_88),
.Y(n_125)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_84),
.B(n_106),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_23),
.Y(n_88)
);

CKINVDCx12_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_89),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_30),
.B1(n_35),
.B2(n_38),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_105),
.B1(n_109),
.B2(n_112),
.Y(n_117)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_35),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_97),
.B(n_111),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_98),
.Y(n_137)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_99),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_53),
.A2(n_28),
.B1(n_27),
.B2(n_29),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_58),
.C(n_63),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_28),
.C(n_25),
.Y(n_150)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_55),
.A2(n_26),
.B1(n_39),
.B2(n_38),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_59),
.A2(n_39),
.B1(n_37),
.B2(n_36),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_45),
.B(n_47),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_70),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_61),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_26),
.B(n_37),
.C(n_36),
.Y(n_127)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_67),
.A3(n_87),
.B1(n_105),
.B2(n_25),
.Y(n_166)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_40),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_98),
.B(n_61),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_138),
.A2(n_151),
.B(n_153),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_85),
.A2(n_57),
.B1(n_28),
.B2(n_27),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_100),
.B1(n_92),
.B2(n_115),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_62),
.A3(n_27),
.B1(n_17),
.B2(n_41),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_75),
.B(n_60),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_115),
.A2(n_27),
.B1(n_32),
.B2(n_41),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

OR2x2_ASAP7_75t_SL g146 ( 
.A(n_97),
.B(n_27),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_25),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_150),
.B(n_80),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_77),
.B(n_34),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_81),
.B(n_34),
.Y(n_153)
);

BUFx10_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_118),
.A2(n_117),
.B1(n_122),
.B2(n_150),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_177),
.B1(n_189),
.B2(n_186),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_112),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_160),
.B(n_167),
.Y(n_209)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_161),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_169),
.Y(n_194)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_103),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_103),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_190),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_172),
.A2(n_180),
.B1(n_187),
.B2(n_124),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_148),
.B(n_68),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_173),
.B(n_174),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_34),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_86),
.B1(n_91),
.B2(n_83),
.Y(n_177)
);

INVxp67_ASAP7_75t_SL g178 ( 
.A(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_130),
.A2(n_92),
.B1(n_86),
.B2(n_67),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_188),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_151),
.A2(n_87),
.B1(n_80),
.B2(n_104),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_182),
.A2(n_153),
.B(n_138),
.Y(n_198)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_192),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_125),
.B(n_33),
.Y(n_185)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_124),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_135),
.A2(n_99),
.B1(n_41),
.B2(n_32),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_119),
.A2(n_91),
.B1(n_68),
.B2(n_28),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_119),
.B(n_33),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_127),
.B(n_33),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_17),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_138),
.B(n_151),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_153),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_159),
.B(n_171),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_149),
.B1(n_141),
.B2(n_142),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_199),
.A2(n_212),
.B1(n_221),
.B2(n_170),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_162),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_201),
.B(n_222),
.Y(n_239)
);

AOI22x1_ASAP7_75t_SL g212 ( 
.A1(n_164),
.A2(n_17),
.B1(n_32),
.B2(n_99),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_141),
.B1(n_142),
.B2(n_126),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_179),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_157),
.B(n_134),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_217),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_135),
.Y(n_218)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_0),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_158),
.B(n_192),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_172),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_162),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_227),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_191),
.A2(n_137),
.B1(n_133),
.B2(n_2),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_225),
.Y(n_248)
);

AND2x6_ASAP7_75t_L g227 ( 
.A(n_163),
.B(n_158),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_235),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_230),
.B(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_234),
.A2(n_242),
.B1(n_226),
.B2(n_224),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_194),
.A2(n_168),
.B1(n_165),
.B2(n_181),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_155),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_240),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_155),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_250),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_139),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_195),
.Y(n_263)
);

NAND2x1_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_212),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_218),
.A2(n_194),
.B(n_198),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_193),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_196),
.B(n_0),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_203),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_251)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_247),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_268),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_218),
.B(n_197),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_265),
.B(n_229),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_227),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_269),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_263),
.B(n_244),
.Y(n_270)
);

AO21x1_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_245),
.B(n_248),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_222),
.B(n_210),
.Y(n_265)
);

OAI322xp33_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_228),
.A3(n_209),
.B1(n_200),
.B2(n_213),
.C1(n_226),
.C2(n_211),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_232),
.B(n_230),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_239),
.B(n_224),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_246),
.A2(n_207),
.B1(n_205),
.B2(n_211),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_272),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_236),
.B(n_237),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_271),
.A2(n_278),
.B(n_279),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_276),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_251),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_281),
.B(n_257),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_280),
.A2(n_262),
.B1(n_260),
.B2(n_256),
.Y(n_283)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_245),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_254),
.B(n_259),
.C(n_258),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_282),
.B(n_278),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_289),
.B(n_233),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_238),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_296),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_207),
.Y(n_296)
);

XOR2x2_ASAP7_75t_SL g298 ( 
.A(n_292),
.B(n_285),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_283),
.Y(n_299)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_299),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_290),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_8),
.B1(n_13),
.B2(n_14),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_298),
.B1(n_300),
.B2(n_287),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_304),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_302),
.B(n_14),
.Y(n_306)
);

AOI221xp5_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_1),
.B1(n_2),
.B2(n_274),
.C(n_227),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_307),
.Y(n_309)
);


endmodule