module real_jpeg_30689_n_19 (n_17, n_8, n_0, n_2, n_697, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_697;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_682;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_109;
wire n_686;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_667;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_602;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_694;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_690;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_659;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g289 ( 
.A(n_0),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_SL g348 ( 
.A(n_1),
.B(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_1),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_1),
.B(n_164),
.Y(n_411)
);

OAI32xp33_ASAP7_75t_L g438 ( 
.A1(n_1),
.A2(n_54),
.A3(n_439),
.B1(n_443),
.B2(n_450),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_1),
.A2(n_382),
.B1(n_483),
.B2(n_485),
.Y(n_482)
);

OAI32xp33_ASAP7_75t_L g490 ( 
.A1(n_1),
.A2(n_54),
.A3(n_439),
.B1(n_443),
.B2(n_450),
.Y(n_490)
);

OAI21xp33_ASAP7_75t_L g550 ( 
.A1(n_1),
.A2(n_95),
.B(n_551),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_2),
.A2(n_137),
.B1(n_141),
.B2(n_142),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_2),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_2),
.A2(n_141),
.B1(n_239),
.B2(n_242),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_2),
.A2(n_141),
.B1(n_292),
.B2(n_297),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_2),
.A2(n_141),
.B1(n_405),
.B2(n_409),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_3),
.Y(n_168)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_3),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_4),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_4),
.A2(n_64),
.B1(n_148),
.B2(n_153),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_4),
.A2(n_64),
.B1(n_329),
.B2(n_331),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_4),
.A2(n_64),
.B1(n_184),
.B2(n_602),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_5),
.Y(n_695)
);

AO22x1_ASAP7_75t_SL g86 ( 
.A1(n_6),
.A2(n_87),
.B1(n_92),
.B2(n_94),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_6),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_6),
.A2(n_94),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_6),
.A2(n_94),
.B1(n_614),
.B2(n_616),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_6),
.A2(n_94),
.B1(n_671),
.B2(n_673),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_7),
.A2(n_271),
.B1(n_272),
.B2(n_275),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_7),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_7),
.A2(n_271),
.B1(n_386),
.B2(n_390),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_7),
.A2(n_271),
.B1(n_474),
.B2(n_478),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_SL g497 ( 
.A1(n_7),
.A2(n_271),
.B1(n_498),
.B2(n_501),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_8),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_8),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_8),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_10),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_11),
.A2(n_179),
.B1(n_180),
.B2(n_184),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_11),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_11),
.A2(n_179),
.B1(n_317),
.B2(n_321),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g433 ( 
.A1(n_11),
.A2(n_179),
.B1(n_373),
.B2(n_434),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g507 ( 
.A1(n_11),
.A2(n_179),
.B1(n_508),
.B2(n_510),
.Y(n_507)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_13),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_13),
.A2(n_53),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_13),
.A2(n_53),
.B1(n_282),
.B2(n_285),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_13),
.A2(n_53),
.B1(n_379),
.B2(n_607),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_14),
.A2(n_103),
.B1(n_106),
.B2(n_109),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_14),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_14),
.A2(n_109),
.B1(n_205),
.B2(n_209),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_14),
.A2(n_109),
.B1(n_618),
.B2(n_622),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_14),
.A2(n_109),
.B1(n_656),
.B2(n_659),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_15),
.B(n_688),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_15),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_17),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_17),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_17),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_17),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_18),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_18),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_18),
.A2(n_160),
.B1(n_171),
.B2(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_18),
.A2(n_160),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_SL g460 ( 
.A1(n_18),
.A2(n_104),
.B1(n_160),
.B2(n_461),
.Y(n_460)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_682),
.B(n_686),
.C(n_690),
.Y(n_19)
);

INVxp67_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

AO21x2_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_593),
.B(n_676),
.Y(n_21)
);

NAND2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_419),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_359),
.B(n_415),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_25),
.B(n_590),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_246),
.B(n_300),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_26),
.B(n_246),
.Y(n_418)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_27),
.B(n_247),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_199),
.Y(n_27)
);

INVxp33_ASAP7_75t_SL g643 ( 
.A(n_28),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_110),
.C(n_154),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_30),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_80),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_31),
.B(n_80),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_48),
.B1(n_58),
.B2(n_69),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_32),
.A2(n_48),
.B1(n_69),
.B2(n_204),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_32),
.A2(n_58),
.B1(n_69),
.B2(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_32),
.A2(n_69),
.B1(n_433),
.B2(n_473),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_32),
.B(n_382),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_33),
.A2(n_203),
.B1(n_212),
.B2(n_213),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_33),
.A2(n_212),
.B1(n_371),
.B2(n_375),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_33),
.B(n_371),
.Y(n_436)
);

AO22x1_ASAP7_75t_L g576 ( 
.A1(n_33),
.A2(n_212),
.B1(n_371),
.B2(n_577),
.Y(n_576)
);

OA21x2_ASAP7_75t_L g625 ( 
.A1(n_33),
.A2(n_212),
.B(n_213),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_70),
.Y(n_69)
);

OAI22x1_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_42),
.B2(n_45),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_37),
.Y(n_522)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_44),
.Y(n_463)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_46),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_52),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_52),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_56),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_57),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_57),
.Y(n_544)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g296 ( 
.A(n_63),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_63),
.Y(n_455)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_69),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_SL g432 ( 
.A1(n_69),
.A2(n_433),
.B(n_436),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_74),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_78),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_79),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_85),
.B1(n_95),
.B2(n_102),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_84),
.Y(n_562)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_86),
.A2(n_96),
.B(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_91),
.Y(n_284)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_91),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_93),
.Y(n_332)
);

BUFx2_ASAP7_75t_SL g500 ( 
.A(n_93),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_95),
.A2(n_102),
.B1(n_280),
.B2(n_286),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_95),
.A2(n_286),
.B1(n_328),
.B2(n_404),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_95),
.A2(n_507),
.B(n_551),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_96),
.A2(n_281),
.B1(n_327),
.B2(n_333),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_96),
.B(n_460),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_96),
.A2(n_496),
.B1(n_504),
.B2(n_506),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_98),
.Y(n_330)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_98),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_98),
.Y(n_533)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_101),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_101),
.Y(n_335)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_101),
.Y(n_556)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_105),
.Y(n_285)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_108),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_110),
.A2(n_111),
.B1(n_154),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_136),
.B1(n_146),
.B2(n_147),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_112),
.A2(n_147),
.B1(n_219),
.B2(n_224),
.Y(n_218)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_112),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_112),
.A2(n_385),
.B1(n_392),
.B2(n_393),
.Y(n_384)
);

AO22x1_ASAP7_75t_SL g402 ( 
.A1(n_112),
.A2(n_146),
.B1(n_262),
.B2(n_385),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_112),
.A2(n_393),
.B1(n_613),
.B2(n_617),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_112),
.A2(n_219),
.B1(n_224),
.B2(n_617),
.Y(n_630)
);

OAI21xp33_ASAP7_75t_L g652 ( 
.A1(n_112),
.A2(n_146),
.B(n_613),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_122),
.Y(n_112)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_113),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_118),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_119),
.Y(n_214)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_127),
.B1(n_130),
.B2(n_133),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_125),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g621 ( 
.A(n_126),
.Y(n_621)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_136),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_140),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_140),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g320 ( 
.A(n_140),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_140),
.Y(n_355)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_145),
.Y(n_389)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_145),
.Y(n_445)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_145),
.Y(n_624)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_146),
.Y(n_225)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_152),
.Y(n_339)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_154),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_177),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_155),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_164),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_156),
.B(n_185),
.Y(n_236)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

BUFx4f_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g660 ( 
.A(n_158),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_159),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_159),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_159),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_159),
.Y(n_608)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_163),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_163),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_164),
.B(n_238),
.Y(n_237)
);

AO22x2_ASAP7_75t_SL g269 ( 
.A1(n_164),
.A2(n_178),
.B1(n_185),
.B2(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_164),
.B(n_270),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_164),
.Y(n_610)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_169),
.B1(n_171),
.B2(n_174),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_168),
.Y(n_342)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_170),
.Y(n_484)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_171),
.Y(n_616)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_172),
.Y(n_322)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_172),
.Y(n_615)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_185),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_183),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_185),
.B(n_378),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_185),
.Y(n_605)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_190),
.B1(n_192),
.B2(n_195),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_189),
.Y(n_274)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_198),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_227),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_200),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_226),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_218),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_218),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_208),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_212),
.B(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_217),
.Y(n_435)
);

BUFx4f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_223),
.Y(n_487)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22x1_ASAP7_75t_L g260 ( 
.A1(n_225),
.A2(n_261),
.B1(n_267),
.B2(n_268),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_225),
.B(n_382),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_226),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_227),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_SL g637 ( 
.A1(n_228),
.A2(n_256),
.B(n_638),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_229),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_231),
.Y(n_230)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_233),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_235),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_236),
.B(n_312),
.Y(n_311)
);

AOI22x1_ASAP7_75t_SL g627 ( 
.A1(n_238),
.A2(n_601),
.B1(n_605),
.B2(n_610),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.C(n_257),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_248),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_253),
.B(n_258),
.Y(n_302)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVxp33_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_269),
.C(n_278),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_260),
.B(n_269),
.Y(n_306)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_262),
.B(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_265),
.Y(n_442)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_267),
.A2(n_316),
.B(n_323),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_267),
.A2(n_323),
.B(n_482),
.Y(n_481)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_277),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_306),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_290),
.Y(n_278)
);

XNOR2x2_ASAP7_75t_L g368 ( 
.A(n_279),
.B(n_290),
.Y(n_368)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_285),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_286),
.A2(n_459),
.B(n_497),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_288),
.Y(n_505)
);

INVx8_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx8_ASAP7_75t_L g458 ( 
.A(n_289),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_291),
.Y(n_375)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_298),
.Y(n_372)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_299),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_301),
.B(n_303),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.C(n_309),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_305),
.B(n_308),
.Y(n_362)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_L g361 ( 
.A(n_309),
.B(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_313),
.C(n_325),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_310),
.A2(n_311),
.B1(n_314),
.B2(n_315),
.Y(n_366)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_324),
.Y(n_393)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_325),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_336),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_326),
.B(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

AOI32xp33_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_340),
.A3(n_343),
.B1(n_348),
.B2(n_351),
.Y(n_336)
);

AOI32xp33_ASAP7_75t_L g399 ( 
.A1(n_337),
.A2(n_340),
.A3(n_343),
.B1(n_348),
.B2(n_351),
.Y(n_399)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_348),
.Y(n_383)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_356),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.C(n_394),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

OAI21xp33_ASAP7_75t_L g590 ( 
.A1(n_361),
.A2(n_591),
.B(n_592),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_363),
.Y(n_591)
);

MAJx2_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_368),
.C(n_369),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_364),
.A2(n_365),
.B1(n_413),
.B2(n_414),
.Y(n_412)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

XNOR2x1_ASAP7_75t_L g413 ( 
.A(n_368),
.B(n_369),
.Y(n_413)
);

MAJx2_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_376),
.C(n_384),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_384),
.Y(n_397)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_397),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_379),
.A2(n_382),
.B(n_383),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx8_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_382),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_382),
.B(n_454),
.Y(n_537)
);

OAI21xp33_ASAP7_75t_SL g540 ( 
.A1(n_382),
.A2(n_537),
.B(n_541),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_382),
.B(n_559),
.Y(n_558)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_391),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_412),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_395),
.B(n_412),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_398),
.C(n_400),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_396),
.B(n_423),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_423),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_398),
.A2(n_400),
.B1(n_401),
.B2(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_398),
.Y(n_424)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.C(n_410),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_402),
.B(n_429),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_403),
.A2(n_410),
.B1(n_411),
.B2(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_403),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_404),
.A2(n_457),
.B(n_459),
.Y(n_456)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_413),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_417),
.B(n_418),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_589),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_464),
.B(n_588),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_425),
.B(n_426),
.Y(n_421)
);

NAND3xp33_ASAP7_75t_L g588 ( 
.A(n_422),
.B(n_425),
.C(n_426),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_431),
.C(n_437),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_428),
.B(n_467),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_431),
.A2(n_432),
.B1(n_437),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_436),
.B(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_437),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_456),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NAND2xp67_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_446),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx5_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_490),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_SL g551 ( 
.A(n_460),
.B(n_552),
.Y(n_551)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_461),
.Y(n_509)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

AOI21x1_ASAP7_75t_L g464 ( 
.A1(n_465),
.A2(n_492),
.B(n_587),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_SL g587 ( 
.A(n_466),
.B(n_469),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_488),
.B(n_491),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_480),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_471),
.B(n_480),
.Y(n_491)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_472),
.B(n_481),
.Y(n_571)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_473),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_477),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_489),
.B(n_571),
.Y(n_570)
);

OAI321xp33_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_569),
.A3(n_580),
.B1(n_585),
.B2(n_586),
.C(n_697),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_545),
.B(n_568),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_516),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_495),
.B(n_516),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_505),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_538),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_517),
.B(n_538),
.Y(n_581)
);

AOI21xp33_ASAP7_75t_L g517 ( 
.A1(n_518),
.A2(n_523),
.B(n_529),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_527),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_530),
.A2(n_534),
.B(n_537),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_535),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_542),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_546),
.A2(n_549),
.B(n_567),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_548),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_547),
.B(n_548),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_550),
.B(n_557),
.Y(n_549)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx3_ASAP7_75t_SL g553 ( 
.A(n_554),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g557 ( 
.A(n_558),
.B(n_563),
.Y(n_557)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_570),
.B(n_572),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_570),
.B(n_572),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_573),
.B(n_574),
.C(n_578),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_573),
.B(n_583),
.Y(n_582)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_575),
.A2(n_576),
.B1(n_579),
.B2(n_584),
.Y(n_583)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_579),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_581),
.B(n_582),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_581),
.B(n_582),
.Y(n_585)
);

NOR3xp33_ASAP7_75t_L g593 ( 
.A(n_594),
.B(n_647),
.C(n_668),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_595),
.B(n_639),
.Y(n_594)
);

A2O1A1Ixp33_ASAP7_75t_SL g678 ( 
.A1(n_595),
.A2(n_648),
.B(n_679),
.C(n_680),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_596),
.B(n_631),
.Y(n_595)
);

NOR2xp67_ASAP7_75t_SL g680 ( 
.A(n_596),
.B(n_631),
.Y(n_680)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_597),
.B(n_628),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_598),
.B(n_626),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_598),
.Y(n_667)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_599),
.B(n_611),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_599),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_600),
.A2(n_604),
.B1(n_606),
.B2(n_609),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_605),
.A2(n_610),
.B1(n_654),
.B2(n_655),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_605),
.A2(n_610),
.B1(n_655),
.B2(n_670),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_605),
.A2(n_610),
.B(n_670),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_606),
.Y(n_654)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_608),
.Y(n_672)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

XNOR2x1_ASAP7_75t_L g611 ( 
.A(n_612),
.B(n_625),
.Y(n_611)
);

INVxp33_ASAP7_75t_L g665 ( 
.A(n_612),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_623),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_624),
.Y(n_623)
);

MAJx2_ASAP7_75t_L g628 ( 
.A(n_625),
.B(n_627),
.C(n_629),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_625),
.A2(n_629),
.B1(n_630),
.B2(n_634),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_625),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_626),
.B(n_628),
.C(n_667),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_627),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_627),
.B(n_633),
.Y(n_632)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_632),
.B(n_635),
.C(n_636),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_632),
.B(n_645),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_SL g663 ( 
.A(n_634),
.B(n_664),
.C(n_665),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_635),
.A2(n_636),
.B1(n_637),
.B2(n_646),
.Y(n_645)
);

INVxp67_ASAP7_75t_SL g646 ( 
.A(n_635),
.Y(n_646)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_637),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_640),
.B(n_644),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_640),
.B(n_644),
.Y(n_679)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_641),
.B(n_642),
.C(n_643),
.Y(n_640)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_648),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_649),
.B(n_666),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_649),
.B(n_666),
.Y(n_677)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_650),
.B(n_663),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_SL g650 ( 
.A1(n_651),
.A2(n_653),
.B1(n_661),
.B2(n_662),
.Y(n_650)
);

CKINVDCx16_ASAP7_75t_R g661 ( 
.A(n_651),
.Y(n_661)
);

BUFx4_ASAP7_75t_R g651 ( 
.A(n_652),
.Y(n_651)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_653),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_653),
.B(n_661),
.C(n_663),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_657),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_658),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_658),
.Y(n_674)
);

INVx11_ASAP7_75t_L g659 ( 
.A(n_660),
.Y(n_659)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_668),
.A2(n_677),
.B(n_678),
.C(n_681),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_669),
.B(n_675),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_669),
.B(n_675),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_669),
.B(n_684),
.Y(n_683)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_669),
.Y(n_689)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_672),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_674),
.Y(n_673)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_683),
.Y(n_682)
);

CKINVDCx16_ASAP7_75t_R g684 ( 
.A(n_685),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_685),
.B(n_689),
.Y(n_688)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_687),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_691),
.B(n_695),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_692),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_693),
.Y(n_692)
);

BUFx12_ASAP7_75t_L g693 ( 
.A(n_694),
.Y(n_693)
);


endmodule