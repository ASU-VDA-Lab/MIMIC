module fake_jpeg_10882_n_557 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_557);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_557;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_11),
.B(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_60),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_61),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_62),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_63),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_64),
.B(n_66),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_15),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_65),
.B(n_93),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_25),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_68),
.Y(n_136)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx5_ASAP7_75t_SL g147 ( 
.A(n_73),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_74),
.A2(n_57),
.B1(n_54),
.B2(n_49),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_77),
.Y(n_176)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_83),
.B(n_88),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_84),
.Y(n_211)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_85),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_87),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_40),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_24),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_91),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_42),
.B(n_31),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_92),
.B(n_94),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_35),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_26),
.B(n_14),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g184 ( 
.A(n_95),
.Y(n_184)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_96),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_37),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_97),
.B(n_44),
.Y(n_153)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_35),
.B(n_1),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_33),
.Y(n_131)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_100),
.Y(n_172)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

BUFx10_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_104),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_52),
.B(n_1),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_107),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_29),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_29),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_114),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_37),
.Y(n_112)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_26),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_113),
.B(n_2),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_29),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_29),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_116),
.B(n_118),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_21),
.Y(n_118)
);

BUFx8_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_21),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_23),
.Y(n_175)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_32),
.Y(n_124)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_32),
.Y(n_125)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g236 ( 
.A(n_131),
.B(n_185),
.C(n_13),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_87),
.A2(n_23),
.B1(n_51),
.B2(n_45),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_134),
.A2(n_191),
.B1(n_197),
.B2(n_198),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_153),
.B(n_126),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_103),
.A2(n_44),
.B(n_34),
.Y(n_154)
);

OR2x2_ASAP7_75t_SL g221 ( 
.A(n_154),
.B(n_85),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_157),
.A2(n_173),
.B1(n_195),
.B2(n_203),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_91),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_167),
.B(n_170),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_89),
.B(n_44),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_74),
.A2(n_34),
.B1(n_54),
.B2(n_49),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_174),
.B(n_187),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_204),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_97),
.A2(n_19),
.B1(n_51),
.B2(n_30),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_177),
.A2(n_189),
.B(n_190),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_103),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_179),
.B(n_180),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_73),
.B(n_57),
.Y(n_180)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_68),
.A2(n_47),
.B(n_41),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_112),
.B(n_36),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_73),
.B(n_47),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_188),
.B(n_194),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_80),
.A2(n_19),
.B1(n_30),
.B2(n_45),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_61),
.A2(n_19),
.B1(n_39),
.B2(n_36),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_63),
.A2(n_41),
.B1(n_39),
.B2(n_33),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_82),
.B(n_4),
.C(n_5),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_193),
.B(n_206),
.C(n_177),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_89),
.B(n_4),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_58),
.A2(n_95),
.B1(n_75),
.B2(n_67),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_98),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_100),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_120),
.A2(n_121),
.B1(n_125),
.B2(n_117),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_200),
.A2(n_206),
.B1(n_84),
.B2(n_110),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_59),
.A2(n_14),
.B1(n_9),
.B2(n_10),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_96),
.B(n_8),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_104),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_81),
.B1(n_62),
.B2(n_60),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_120),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_206)
);

INVx6_ASAP7_75t_SL g212 ( 
.A(n_147),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_212),
.Y(n_332)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_213),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_147),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_214),
.B(n_220),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_146),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_215),
.B(n_233),
.Y(n_286)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_216),
.Y(n_321)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_171),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g294 ( 
.A1(n_221),
.A2(n_236),
.B(n_240),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_165),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_222),
.B(n_232),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_223),
.Y(n_318)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_224),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_225),
.A2(n_258),
.B1(n_260),
.B2(n_265),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_226),
.A2(n_231),
.B1(n_263),
.B2(n_276),
.Y(n_326)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_228),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_158),
.B(n_78),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_229),
.B(n_234),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_135),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_205),
.A2(n_102),
.B1(n_119),
.B2(n_86),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_135),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_137),
.B(n_105),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_176),
.B(n_12),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_153),
.A2(n_119),
.B(n_115),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_235),
.A2(n_276),
.B(n_244),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_148),
.B(n_14),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_237),
.B(n_242),
.Y(n_303)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_238),
.Y(n_327)
);

INVx2_ASAP7_75t_R g240 ( 
.A(n_136),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_168),
.B(n_199),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_127),
.B(n_149),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_243),
.B(n_247),
.Y(n_305)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_186),
.Y(n_244)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_245),
.Y(n_337)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_169),
.Y(n_246)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_246),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_128),
.B(n_183),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_181),
.B(n_196),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_248),
.B(n_264),
.Y(n_308)
);

BUFx8_ASAP7_75t_L g250 ( 
.A(n_135),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_250),
.Y(n_302)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_145),
.Y(n_251)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_252),
.Y(n_296)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_253),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_141),
.Y(n_254)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_186),
.A2(n_132),
.B1(n_184),
.B2(n_166),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_152),
.Y(n_256)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_256),
.Y(n_324)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_139),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_257),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_141),
.Y(n_258)
);

BUFx16f_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_259),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_132),
.A2(n_184),
.B1(n_144),
.B2(n_130),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_169),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_261),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_190),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_150),
.Y(n_264)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_126),
.Y(n_265)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_145),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_266),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_155),
.B(n_201),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_267),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_136),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_270),
.Y(n_310)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_207),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_144),
.A2(n_130),
.B1(n_159),
.B2(n_140),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_160),
.B(n_138),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_274),
.B(n_275),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_191),
.B(n_134),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_276),
.B(n_277),
.Y(n_320)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_211),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_278),
.A2(n_281),
.B1(n_254),
.B2(n_212),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_140),
.B(n_159),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_279),
.B(n_283),
.Y(n_322)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_211),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_189),
.B(n_208),
.C(n_161),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_282),
.B(n_235),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_208),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_262),
.A2(n_162),
.B1(n_164),
.B2(n_161),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_291),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_262),
.A2(n_162),
.B1(n_164),
.B2(n_143),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_275),
.A2(n_133),
.B1(n_178),
.B2(n_163),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_249),
.A2(n_163),
.B1(n_210),
.B2(n_277),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_234),
.A2(n_163),
.B1(n_210),
.B2(n_249),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_313),
.A2(n_315),
.B1(n_328),
.B2(n_330),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_221),
.A2(n_210),
.B1(n_282),
.B2(n_263),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_323),
.B(n_334),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_325),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_326),
.A2(n_329),
.B1(n_278),
.B2(n_281),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_280),
.A2(n_226),
.B1(n_242),
.B2(n_227),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_231),
.A2(n_248),
.B1(n_247),
.B2(n_243),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_229),
.A2(n_279),
.B1(n_239),
.B2(n_219),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_240),
.B(n_245),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_336),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_218),
.A2(n_228),
.B1(n_213),
.B2(n_238),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_333),
.A2(n_335),
.B1(n_257),
.B2(n_265),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_246),
.A2(n_261),
.B1(n_268),
.B2(n_251),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_264),
.B(n_270),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_336),
.Y(n_338)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_338),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_297),
.B(n_230),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_339),
.B(n_341),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_292),
.Y(n_340)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_300),
.B(n_241),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_322),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_343),
.Y(n_384)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_347),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_331),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_345),
.B(n_350),
.Y(n_381)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_285),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_292),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_348),
.B(n_349),
.Y(n_380)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_317),
.B(n_230),
.Y(n_350)
);

AND2x2_ASAP7_75t_SL g351 ( 
.A(n_320),
.B(n_250),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_324),
.Y(n_387)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_301),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_355),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_328),
.A2(n_266),
.B1(n_224),
.B2(n_272),
.Y(n_353)
);

OA22x2_ASAP7_75t_L g383 ( 
.A1(n_353),
.A2(n_359),
.B1(n_373),
.B2(n_377),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_319),
.B(n_334),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g392 ( 
.A1(n_354),
.A2(n_366),
.B(n_370),
.C(n_371),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_241),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_303),
.B(n_271),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_358),
.B(n_361),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_286),
.B(n_258),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_296),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_365),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_259),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_363),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_259),
.Y(n_364)
);

XNOR2x1_ASAP7_75t_L g409 ( 
.A(n_364),
.B(n_295),
.Y(n_409)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_367),
.A2(n_379),
.B1(n_312),
.B2(n_314),
.Y(n_393)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_309),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_370),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_291),
.A2(n_250),
.B1(n_315),
.B2(n_319),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_369),
.A2(n_372),
.B1(n_378),
.B2(n_327),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_305),
.B(n_289),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_305),
.B(n_289),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_371),
.B(n_375),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_307),
.A2(n_326),
.B1(n_329),
.B2(n_308),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_311),
.A2(n_333),
.B1(n_335),
.B2(n_321),
.Y(n_373)
);

OAI21xp33_ASAP7_75t_L g374 ( 
.A1(n_294),
.A2(n_308),
.B(n_310),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_374),
.A2(n_337),
.B(n_318),
.Y(n_397)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_309),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_310),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_376),
.Y(n_385)
);

AO21x2_ASAP7_75t_L g377 ( 
.A1(n_332),
.A2(n_298),
.B(n_316),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_311),
.A2(n_321),
.B1(n_284),
.B2(n_323),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_284),
.A2(n_314),
.B1(n_288),
.B2(n_324),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_354),
.A2(n_302),
.B(n_318),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_382),
.Y(n_418)
);

XNOR2x1_ASAP7_75t_L g432 ( 
.A(n_387),
.B(n_392),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_299),
.C(n_302),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_394),
.C(n_399),
.Y(n_417)
);

NAND2x1_ASAP7_75t_SL g391 ( 
.A(n_342),
.B(n_312),
.Y(n_391)
);

OAI21xp33_ASAP7_75t_L g442 ( 
.A1(n_391),
.A2(n_397),
.B(n_377),
.Y(n_442)
);

OAI22xp33_ASAP7_75t_L g420 ( 
.A1(n_393),
.A2(n_359),
.B1(n_346),
.B2(n_338),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_366),
.B(n_288),
.C(n_290),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_379),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_398),
.B(n_404),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_337),
.C(n_293),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_367),
.A2(n_301),
.B1(n_293),
.B2(n_327),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_401),
.A2(n_340),
.B1(n_360),
.B2(n_377),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_356),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_356),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_405),
.B(n_408),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_378),
.A2(n_295),
.B(n_287),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_407),
.B(n_360),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_377),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_410),
.A2(n_346),
.B1(n_347),
.B2(n_351),
.Y(n_426)
);

AO21x1_ASAP7_75t_L g412 ( 
.A1(n_357),
.A2(n_287),
.B(n_372),
.Y(n_412)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_412),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_364),
.B(n_351),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_362),
.C(n_375),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g465 ( 
.A(n_414),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_412),
.A2(n_357),
.B1(n_343),
.B2(n_369),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_415),
.A2(n_420),
.B1(n_428),
.B2(n_433),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_385),
.B(n_376),
.Y(n_419)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_419),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_385),
.B(n_345),
.Y(n_421)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_421),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_404),
.B(n_405),
.Y(n_422)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_422),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_381),
.B(n_344),
.Y(n_423)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_423),
.Y(n_456)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_390),
.Y(n_424)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_424),
.Y(n_463)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_390),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_425),
.B(n_429),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_426),
.A2(n_384),
.B1(n_389),
.B2(n_383),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_441),
.C(n_409),
.Y(n_453)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_390),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_386),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_435),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_412),
.A2(n_377),
.B1(n_365),
.B2(n_368),
.Y(n_433)
);

INVx13_ASAP7_75t_L g434 ( 
.A(n_402),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_434),
.Y(n_450)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_386),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g436 ( 
.A(n_406),
.Y(n_436)
);

NAND3xp33_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_406),
.C(n_411),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_396),
.B(n_340),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_437),
.B(n_438),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_380),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_396),
.B(n_348),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_439),
.B(n_443),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_440),
.B(n_387),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_352),
.C(n_349),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_442),
.A2(n_410),
.B1(n_382),
.B2(n_398),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_421),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_458),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_451),
.A2(n_418),
.B1(n_431),
.B2(n_430),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_426),
.A2(n_408),
.B1(n_400),
.B2(n_403),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_452),
.A2(n_460),
.B1(n_464),
.B2(n_467),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_455),
.C(n_441),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_399),
.C(n_394),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_457),
.B(n_434),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_388),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_462),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_416),
.A2(n_400),
.B1(n_403),
.B2(n_393),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_391),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_416),
.A2(n_384),
.B1(n_401),
.B2(n_389),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_432),
.B(n_391),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_468),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_427),
.B(n_392),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_433),
.A2(n_383),
.B1(n_411),
.B2(n_402),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_470),
.A2(n_431),
.B1(n_429),
.B2(n_425),
.Y(n_475)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_454),
.Y(n_472)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_472),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_473),
.A2(n_475),
.B1(n_476),
.B2(n_479),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_447),
.A2(n_470),
.B1(n_444),
.B2(n_451),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_444),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_477),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_478),
.B(n_480),
.C(n_481),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_447),
.A2(n_443),
.B1(n_422),
.B2(n_435),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_424),
.C(n_440),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_453),
.C(n_457),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_456),
.A2(n_419),
.B1(n_423),
.B2(n_437),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_483),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_465),
.B(n_395),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_484),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_446),
.A2(n_414),
.B(n_438),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_486),
.A2(n_446),
.B(n_462),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_449),
.A2(n_469),
.B1(n_445),
.B2(n_463),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_488),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_449),
.A2(n_415),
.B1(n_439),
.B2(n_428),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_461),
.B(n_380),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_489),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_468),
.B(n_397),
.C(n_407),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_460),
.C(n_383),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_469),
.Y(n_491)
);

INVx13_ASAP7_75t_L g497 ( 
.A(n_491),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_466),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_498),
.A2(n_477),
.B(n_482),
.Y(n_518)
);

BUFx24_ASAP7_75t_SL g499 ( 
.A(n_474),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_499),
.B(n_481),
.Y(n_515)
);

INVx13_ASAP7_75t_L g500 ( 
.A(n_491),
.Y(n_500)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_500),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_490),
.A2(n_450),
.B(n_464),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_501),
.A2(n_486),
.B(n_482),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_471),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_452),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_504),
.B(n_506),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_518),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_476),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_512),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_505),
.A2(n_479),
.B1(n_488),
.B2(n_473),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_511),
.A2(n_498),
.B1(n_472),
.B2(n_494),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_475),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_487),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_513),
.B(n_515),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_480),
.C(n_471),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_496),
.C(n_485),
.Y(n_523)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_493),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_519),
.A2(n_495),
.B1(n_489),
.B2(n_494),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_521),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_501),
.B(n_485),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_523),
.B(n_524),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_506),
.C(n_508),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_514),
.A2(n_503),
.B1(n_497),
.B2(n_500),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_525),
.B(n_528),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_527),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_514),
.A2(n_495),
.B1(n_507),
.B2(n_497),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_511),
.C(n_509),
.Y(n_533)
);

A2O1A1Ixp33_ASAP7_75t_L g532 ( 
.A1(n_518),
.A2(n_492),
.B(n_502),
.C(n_383),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_532),
.A2(n_521),
.B(n_519),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_533),
.B(n_534),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_530),
.A2(n_516),
.B(n_517),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_536),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_523),
.B(n_524),
.C(n_529),
.Y(n_536)
);

AOI21xp33_ASAP7_75t_L g539 ( 
.A1(n_526),
.A2(n_520),
.B(n_434),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_539),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_525),
.A2(n_529),
.B(n_522),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_540),
.B(n_537),
.Y(n_546)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_528),
.B(n_522),
.Y(n_542)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_542),
.Y(n_550)
);

NOR2x1_ASAP7_75t_L g544 ( 
.A(n_536),
.B(n_532),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_544),
.A2(n_546),
.B(n_534),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_548),
.B(n_549),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_547),
.A2(n_538),
.B(n_533),
.Y(n_549)
);

INVxp33_ASAP7_75t_SL g551 ( 
.A(n_545),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_551),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g554 ( 
.A(n_553),
.B(n_550),
.C(n_543),
.Y(n_554)
);

BUFx24_ASAP7_75t_SL g555 ( 
.A(n_554),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_552),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_537),
.Y(n_557)
);


endmodule