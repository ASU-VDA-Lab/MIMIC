module real_aes_17003_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1845;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_1383;
wire n_552;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_1787;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1760;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_1856;
wire n_676;
wire n_658;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1855;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_1838;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_1457;
wire n_1343;
wire n_719;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1176;
wire n_640;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_1777;
wire n_458;
wire n_444;
wire n_1200;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1868;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
XNOR2xp5_ASAP7_75t_L g893 ( .A(n_0), .B(n_894), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g1568 ( .A1(n_0), .A2(n_90), .B1(n_1525), .B2(n_1528), .Y(n_1568) );
OAI22xp33_ASAP7_75t_L g1051 ( .A1(n_1), .A2(n_334), .B1(n_462), .B2(n_842), .Y(n_1051) );
OAI22xp33_ASAP7_75t_SL g1064 ( .A1(n_1), .A2(n_334), .B1(n_505), .B2(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1323 ( .A(n_2), .Y(n_1323) );
INVx1_ASAP7_75t_L g389 ( .A(n_3), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_3), .B(n_399), .Y(n_547) );
AND2x2_ASAP7_75t_L g1732 ( .A(n_3), .B(n_465), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1735 ( .A(n_3), .B(n_268), .Y(n_1735) );
CKINVDCx5p33_ASAP7_75t_R g1180 ( .A(n_4), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_5), .A2(n_273), .B1(n_991), .B2(n_1287), .Y(n_1286) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_5), .A2(n_210), .B1(n_967), .B2(n_978), .Y(n_1303) );
INVx1_ASAP7_75t_L g745 ( .A(n_6), .Y(n_745) );
INVx1_ASAP7_75t_L g1092 ( .A(n_7), .Y(n_1092) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_8), .A2(n_56), .B1(n_391), .B2(n_462), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g646 ( .A1(n_8), .A2(n_56), .B1(n_507), .B2(n_647), .Y(n_646) );
OAI22xp5_ASAP7_75t_SL g1107 ( .A1(n_9), .A2(n_237), .B1(n_489), .B2(n_834), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_9), .A2(n_237), .B1(n_940), .B2(n_1111), .Y(n_1110) );
INVx1_ASAP7_75t_L g1861 ( .A(n_10), .Y(n_1861) );
OAI22xp33_ASAP7_75t_SL g1202 ( .A1(n_11), .A2(n_358), .B1(n_842), .B2(n_1010), .Y(n_1202) );
OAI22xp33_ASAP7_75t_L g1214 ( .A1(n_11), .A2(n_195), .B1(n_505), .B2(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_L g1083 ( .A(n_12), .Y(n_1083) );
INVx1_ASAP7_75t_L g1277 ( .A(n_13), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g1308 ( .A1(n_13), .A2(n_273), .B1(n_978), .B2(n_1309), .Y(n_1308) );
INVx1_ASAP7_75t_L g1740 ( .A(n_14), .Y(n_1740) );
OAI22xp5_ASAP7_75t_L g1782 ( .A1(n_14), .A2(n_362), .B1(n_1783), .B2(n_1787), .Y(n_1782) );
OAI22xp5_ASAP7_75t_L g1862 ( .A1(n_15), .A2(n_159), .B1(n_391), .B2(n_462), .Y(n_1862) );
OAI22xp5_ASAP7_75t_L g1864 ( .A1(n_15), .A2(n_159), .B1(n_503), .B2(n_1215), .Y(n_1864) );
OAI22xp33_ASAP7_75t_L g1108 ( .A1(n_16), .A2(n_158), .B1(n_391), .B2(n_462), .Y(n_1108) );
OAI22xp33_ASAP7_75t_L g1117 ( .A1(n_16), .A2(n_158), .B1(n_507), .B2(n_739), .Y(n_1117) );
INVx1_ASAP7_75t_L g1364 ( .A(n_17), .Y(n_1364) );
OAI221xp5_ASAP7_75t_L g1373 ( .A1(n_17), .A2(n_315), .B1(n_623), .B2(n_1374), .C(n_1375), .Y(n_1373) );
CKINVDCx5p33_ASAP7_75t_R g1223 ( .A(n_18), .Y(n_1223) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_19), .A2(n_317), .B1(n_1061), .B2(n_1062), .Y(n_1060) );
OAI22xp33_ASAP7_75t_L g1069 ( .A1(n_19), .A2(n_317), .B1(n_532), .B2(n_535), .Y(n_1069) );
INVx2_ASAP7_75t_L g441 ( .A(n_20), .Y(n_441) );
OAI22xp33_ASAP7_75t_SL g1421 ( .A1(n_21), .A2(n_285), .B1(n_505), .B2(n_1215), .Y(n_1421) );
OAI22xp33_ASAP7_75t_L g1428 ( .A1(n_21), .A2(n_285), .B1(n_842), .B2(n_873), .Y(n_1428) );
INVx1_ASAP7_75t_L g857 ( .A(n_22), .Y(n_857) );
INVx1_ASAP7_75t_L g1152 ( .A(n_23), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_24), .A2(n_192), .B1(n_971), .B2(n_972), .Y(n_970) );
AOI22xp33_ASAP7_75t_SL g1002 ( .A1(n_24), .A2(n_142), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1380 ( .A1(n_25), .A2(n_300), .B1(n_1381), .B2(n_1383), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_25), .A2(n_165), .B1(n_1390), .B2(n_1392), .Y(n_1389) );
AOI22xp33_ASAP7_75t_SL g1840 ( .A1(n_26), .A2(n_177), .B1(n_991), .B2(n_1841), .Y(n_1840) );
AOI22xp33_ASAP7_75t_L g1850 ( .A1(n_26), .A2(n_221), .B1(n_616), .B2(n_1392), .Y(n_1850) );
INVx1_ASAP7_75t_L g790 ( .A(n_27), .Y(n_790) );
XOR2xp5_ASAP7_75t_L g1828 ( .A(n_28), .B(n_1829), .Y(n_1828) );
INVx1_ASAP7_75t_L g853 ( .A(n_29), .Y(n_853) );
OAI211xp5_ASAP7_75t_L g874 ( .A1(n_30), .A2(n_585), .B(n_875), .C(n_878), .Y(n_874) );
INVx1_ASAP7_75t_L g888 ( .A(n_30), .Y(n_888) );
INVx1_ASAP7_75t_L g1436 ( .A(n_31), .Y(n_1436) );
OAI221xp5_ASAP7_75t_L g1334 ( .A1(n_32), .A2(n_87), .B1(n_535), .B2(n_1215), .C(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1348 ( .A(n_32), .Y(n_1348) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_33), .Y(n_384) );
AND2x2_ASAP7_75t_L g1519 ( .A(n_33), .B(n_382), .Y(n_1519) );
INVx1_ASAP7_75t_L g908 ( .A(n_34), .Y(n_908) );
OAI22xp33_ASAP7_75t_SL g730 ( .A1(n_35), .A2(n_184), .B1(n_489), .B2(n_491), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_35), .A2(n_184), .B1(n_530), .B2(n_720), .Y(n_733) );
OAI222xp33_ASAP7_75t_L g956 ( .A1(n_36), .A2(n_218), .B1(n_356), .B2(n_606), .C1(n_957), .C2(n_958), .Y(n_956) );
OAI222xp33_ASAP7_75t_L g1012 ( .A1(n_36), .A2(n_218), .B1(n_356), .B2(n_633), .C1(n_839), .C2(n_1013), .Y(n_1012) );
CKINVDCx5p33_ASAP7_75t_R g1484 ( .A(n_37), .Y(n_1484) );
AOI22xp33_ASAP7_75t_L g1567 ( .A1(n_38), .A2(n_66), .B1(n_1518), .B2(n_1522), .Y(n_1567) );
INVx1_ASAP7_75t_L g1105 ( .A(n_39), .Y(n_1105) );
INVx1_ASAP7_75t_L g686 ( .A(n_40), .Y(n_686) );
INVx1_ASAP7_75t_L g1141 ( .A(n_41), .Y(n_1141) );
INVx1_ASAP7_75t_L g418 ( .A(n_42), .Y(n_418) );
INVx1_ASAP7_75t_L g612 ( .A(n_43), .Y(n_612) );
INVx1_ASAP7_75t_L g825 ( .A(n_44), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_44), .A2(n_366), .B1(n_594), .B2(n_834), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g1749 ( .A1(n_45), .A2(n_200), .B1(n_1750), .B2(n_1752), .Y(n_1749) );
AOI22xp33_ASAP7_75t_SL g1803 ( .A1(n_45), .A2(n_335), .B1(n_450), .B2(n_821), .Y(n_1803) );
XNOR2x1_ASAP7_75t_L g1399 ( .A(n_46), .B(n_1400), .Y(n_1399) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_47), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g1275 ( .A(n_48), .Y(n_1275) );
INVx1_ASAP7_75t_L g911 ( .A(n_49), .Y(n_911) );
INVx1_ASAP7_75t_L g1035 ( .A(n_50), .Y(n_1035) );
AOI22xp33_ASAP7_75t_SL g1833 ( .A1(n_51), .A2(n_221), .B1(n_1058), .B2(n_1834), .Y(n_1833) );
AOI22xp33_ASAP7_75t_L g1844 ( .A1(n_51), .A2(n_177), .B1(n_1805), .B2(n_1845), .Y(n_1844) );
INVx1_ASAP7_75t_L g1326 ( .A(n_52), .Y(n_1326) );
AOI22xp5_ASAP7_75t_L g1543 ( .A1(n_53), .A2(n_118), .B1(n_1518), .B2(n_1522), .Y(n_1543) );
XOR2x2_ASAP7_75t_L g1725 ( .A(n_53), .B(n_1726), .Y(n_1725) );
AOI22xp33_ASAP7_75t_L g1826 ( .A1(n_53), .A2(n_1827), .B1(n_1868), .B2(n_1870), .Y(n_1826) );
AOI22xp5_ASAP7_75t_L g1533 ( .A1(n_54), .A2(n_277), .B1(n_1518), .B2(n_1522), .Y(n_1533) );
INVx1_ASAP7_75t_L g779 ( .A(n_55), .Y(n_779) );
INVx1_ASAP7_75t_L g1091 ( .A(n_57), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_58), .B(n_523), .Y(n_1336) );
INVxp67_ASAP7_75t_SL g1343 ( .A(n_58), .Y(n_1343) );
OAI211xp5_ASAP7_75t_L g1123 ( .A1(n_59), .A2(n_715), .B(n_1124), .C(n_1126), .Y(n_1123) );
INVx1_ASAP7_75t_L g1133 ( .A(n_59), .Y(n_1133) );
OAI211xp5_ASAP7_75t_L g1195 ( .A1(n_60), .A2(n_567), .B(n_1196), .C(n_1199), .Y(n_1195) );
INVx1_ASAP7_75t_L g1213 ( .A(n_60), .Y(n_1213) );
INVx1_ASAP7_75t_L g1089 ( .A(n_61), .Y(n_1089) );
CKINVDCx5p33_ASAP7_75t_R g1171 ( .A(n_62), .Y(n_1171) );
OAI222xp33_ASAP7_75t_L g1263 ( .A1(n_63), .A2(n_198), .B1(n_572), .B2(n_591), .C1(n_1264), .C2(n_1266), .Y(n_1263) );
OAI222xp33_ASAP7_75t_L g1293 ( .A1(n_63), .A2(n_198), .B1(n_238), .B2(n_1294), .C1(n_1295), .C2(n_1296), .Y(n_1293) );
OAI22xp5_ASAP7_75t_L g1369 ( .A1(n_64), .A2(n_126), .B1(n_1061), .B2(n_1242), .Y(n_1369) );
OAI22xp5_ASAP7_75t_L g1376 ( .A1(n_64), .A2(n_126), .B1(n_532), .B2(n_535), .Y(n_1376) );
OAI211xp5_ASAP7_75t_L g468 ( .A1(n_65), .A2(n_469), .B(n_474), .C(n_479), .Y(n_468) );
INVx1_ASAP7_75t_L g528 ( .A(n_65), .Y(n_528) );
OAI22xp33_ASAP7_75t_L g709 ( .A1(n_67), .A2(n_319), .B1(n_391), .B2(n_462), .Y(n_709) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_67), .A2(n_319), .B1(n_507), .B2(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g880 ( .A(n_68), .Y(n_880) );
OAI211xp5_ASAP7_75t_L g885 ( .A1(n_68), .A2(n_517), .B(n_650), .C(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g1031 ( .A(n_69), .Y(n_1031) );
OAI22xp33_ASAP7_75t_L g1339 ( .A1(n_70), .A2(n_202), .B1(n_505), .B2(n_954), .Y(n_1339) );
INVxp67_ASAP7_75t_SL g1345 ( .A(n_70), .Y(n_1345) );
INVx1_ASAP7_75t_L g1856 ( .A(n_71), .Y(n_1856) );
INVx1_ASAP7_75t_L g1151 ( .A(n_72), .Y(n_1151) );
CKINVDCx5p33_ASAP7_75t_R g1234 ( .A(n_73), .Y(n_1234) );
INVx1_ASAP7_75t_L g1147 ( .A(n_74), .Y(n_1147) );
CKINVDCx5p33_ASAP7_75t_R g1449 ( .A(n_75), .Y(n_1449) );
AOI22xp33_ASAP7_75t_L g1555 ( .A1(n_76), .A2(n_260), .B1(n_1518), .B2(n_1522), .Y(n_1555) );
INVx1_ASAP7_75t_L g1414 ( .A(n_77), .Y(n_1414) );
AOI22xp5_ASAP7_75t_L g1537 ( .A1(n_78), .A2(n_266), .B1(n_1525), .B2(n_1528), .Y(n_1537) );
XNOR2xp5_ASAP7_75t_L g1353 ( .A(n_79), .B(n_1354), .Y(n_1353) );
INVx1_ASAP7_75t_L g1325 ( .A(n_80), .Y(n_1325) );
INVx1_ASAP7_75t_L g757 ( .A(n_81), .Y(n_757) );
INVx1_ASAP7_75t_L g904 ( .A(n_82), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g1538 ( .A1(n_83), .A2(n_104), .B1(n_1518), .B2(n_1539), .Y(n_1538) );
OAI22xp33_ASAP7_75t_L g1426 ( .A1(n_84), .A2(n_117), .B1(n_532), .B2(n_535), .Y(n_1426) );
OAI22xp5_ASAP7_75t_L g1432 ( .A1(n_84), .A2(n_117), .B1(n_1061), .B2(n_1242), .Y(n_1432) );
AO22x1_ASAP7_75t_L g1561 ( .A1(n_85), .A2(n_278), .B1(n_1525), .B2(n_1528), .Y(n_1561) );
XNOR2xp5_ASAP7_75t_L g1473 ( .A(n_86), .B(n_1474), .Y(n_1473) );
OAI22xp33_ASAP7_75t_L g1350 ( .A1(n_87), .A2(n_202), .B1(n_842), .B2(n_873), .Y(n_1350) );
INVx1_ASAP7_75t_L g859 ( .A(n_88), .Y(n_859) );
INVx1_ASAP7_75t_L g1464 ( .A(n_89), .Y(n_1464) );
OAI211xp5_ASAP7_75t_L g1469 ( .A1(n_89), .A2(n_715), .B(n_760), .C(n_1470), .Y(n_1469) );
OAI22xp5_ASAP7_75t_L g1241 ( .A1(n_91), .A2(n_289), .B1(n_842), .B2(n_1242), .Y(n_1241) );
OAI22xp5_ASAP7_75t_SL g1250 ( .A1(n_91), .A2(n_138), .B1(n_505), .B2(n_532), .Y(n_1250) );
INVx1_ASAP7_75t_L g1338 ( .A(n_92), .Y(n_1338) );
INVx1_ASAP7_75t_L g1128 ( .A(n_93), .Y(n_1128) );
OAI211xp5_ASAP7_75t_L g1131 ( .A1(n_93), .A2(n_806), .B(n_836), .C(n_1132), .Y(n_1131) );
CKINVDCx5p33_ASAP7_75t_R g1245 ( .A(n_94), .Y(n_1245) );
CKINVDCx5p33_ASAP7_75t_R g1222 ( .A(n_95), .Y(n_1222) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_96), .A2(n_173), .B1(n_391), .B2(n_873), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_96), .A2(n_173), .B1(n_647), .B2(n_884), .Y(n_883) );
CKINVDCx5p33_ASAP7_75t_R g1170 ( .A(n_97), .Y(n_1170) );
AOI22xp33_ASAP7_75t_SL g1842 ( .A1(n_98), .A2(n_373), .B1(n_1058), .B2(n_1834), .Y(n_1842) );
AOI22xp33_ASAP7_75t_L g1852 ( .A1(n_98), .A2(n_100), .B1(n_1811), .B2(n_1847), .Y(n_1852) );
OAI22xp33_ASAP7_75t_SL g593 ( .A1(n_99), .A2(n_288), .B1(n_594), .B2(n_595), .Y(n_593) );
OAI22xp33_ASAP7_75t_L g653 ( .A1(n_99), .A2(n_288), .B1(n_533), .B2(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g1837 ( .A1(n_100), .A2(n_336), .B1(n_991), .B2(n_1838), .Y(n_1837) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_101), .A2(n_263), .B1(n_998), .B2(n_1381), .Y(n_1384) );
AOI22xp33_ASAP7_75t_L g1393 ( .A1(n_101), .A2(n_181), .B1(n_450), .B2(n_968), .Y(n_1393) );
XOR2xp5_ASAP7_75t_L g1165 ( .A(n_102), .B(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1022 ( .A(n_103), .Y(n_1022) );
INVx1_ASAP7_75t_L g909 ( .A(n_105), .Y(n_909) );
CKINVDCx5p33_ASAP7_75t_R g1487 ( .A(n_106), .Y(n_1487) );
INVx1_ASAP7_75t_L g1146 ( .A(n_107), .Y(n_1146) );
CKINVDCx5p33_ASAP7_75t_R g1230 ( .A(n_108), .Y(n_1230) );
OAI22xp33_ASAP7_75t_L g932 ( .A1(n_109), .A2(n_149), .B1(n_462), .B2(n_842), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_109), .A2(n_135), .B1(n_505), .B2(n_720), .Y(n_934) );
INVx1_ASAP7_75t_L g900 ( .A(n_110), .Y(n_900) );
INVx1_ASAP7_75t_L g913 ( .A(n_111), .Y(n_913) );
INVx1_ASAP7_75t_L g692 ( .A(n_112), .Y(n_692) );
OAI211xp5_ASAP7_75t_L g1461 ( .A1(n_113), .A2(n_697), .B(n_1196), .C(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1471 ( .A(n_113), .Y(n_1471) );
INVx1_ASAP7_75t_L g382 ( .A(n_114), .Y(n_382) );
INVx1_ASAP7_75t_L g624 ( .A(n_115), .Y(n_624) );
INVx1_ASAP7_75t_L g1086 ( .A(n_116), .Y(n_1086) );
AO221x2_ASAP7_75t_L g1628 ( .A1(n_119), .A2(n_348), .B1(n_1525), .B2(n_1528), .C(n_1629), .Y(n_1628) );
OAI22xp33_ASAP7_75t_L g1466 ( .A1(n_120), .A2(n_313), .B1(n_462), .B2(n_490), .Y(n_1466) );
OAI22xp33_ASAP7_75t_L g1472 ( .A1(n_120), .A2(n_168), .B1(n_532), .B2(n_535), .Y(n_1472) );
XOR2xp5_ASAP7_75t_L g1256 ( .A(n_121), .B(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1407 ( .A(n_122), .Y(n_1407) );
INVx1_ASAP7_75t_L g1404 ( .A(n_123), .Y(n_1404) );
INVx1_ASAP7_75t_L g728 ( .A(n_124), .Y(n_728) );
CKINVDCx5p33_ASAP7_75t_R g928 ( .A(n_125), .Y(n_928) );
INVx1_ASAP7_75t_L g674 ( .A(n_127), .Y(n_674) );
INVx1_ASAP7_75t_L g589 ( .A(n_128), .Y(n_589) );
INVxp67_ASAP7_75t_SL g1756 ( .A(n_129), .Y(n_1756) );
AOI22xp33_ASAP7_75t_L g1804 ( .A1(n_129), .A2(n_280), .B1(n_1805), .B2(n_1806), .Y(n_1804) );
INVx1_ASAP7_75t_L g748 ( .A(n_130), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_131), .A2(n_207), .B1(n_449), .B2(n_452), .Y(n_448) );
INVx1_ASAP7_75t_L g551 ( .A(n_131), .Y(n_551) );
INVx1_ASAP7_75t_L g1039 ( .A(n_132), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_133), .A2(n_271), .B1(n_953), .B2(n_954), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_133), .A2(n_271), .B1(n_594), .B2(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1127 ( .A(n_134), .Y(n_1127) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_135), .A2(n_232), .B1(n_594), .B2(n_931), .Y(n_930) );
OAI22xp33_ASAP7_75t_SL g1247 ( .A1(n_136), .A2(n_138), .B1(n_873), .B2(n_1061), .Y(n_1247) );
OAI22xp5_ASAP7_75t_L g1254 ( .A1(n_136), .A2(n_141), .B1(n_1210), .B2(n_1211), .Y(n_1254) );
INVx1_ASAP7_75t_L g1737 ( .A(n_137), .Y(n_1737) );
OAI22xp33_ASAP7_75t_L g1812 ( .A1(n_137), .A2(n_190), .B1(n_1813), .B2(n_1816), .Y(n_1812) );
INVx1_ASAP7_75t_L g1054 ( .A(n_139), .Y(n_1054) );
INVxp67_ASAP7_75t_SL g1748 ( .A(n_140), .Y(n_1748) );
AOI22xp33_ASAP7_75t_SL g1807 ( .A1(n_140), .A2(n_212), .B1(n_1390), .B2(n_1808), .Y(n_1807) );
INVx1_ASAP7_75t_L g1246 ( .A(n_141), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_142), .A2(n_310), .B1(n_980), .B2(n_981), .Y(n_979) );
INVx1_ASAP7_75t_L g1144 ( .A(n_143), .Y(n_1144) );
INVx1_ASAP7_75t_L g1357 ( .A(n_144), .Y(n_1357) );
AO22x1_ASAP7_75t_L g1524 ( .A1(n_145), .A2(n_352), .B1(n_1525), .B2(n_1528), .Y(n_1524) );
INVx1_ASAP7_75t_L g1425 ( .A(n_146), .Y(n_1425) );
OAI211xp5_ASAP7_75t_L g1429 ( .A1(n_146), .A2(n_1023), .B(n_1196), .C(n_1430), .Y(n_1429) );
CKINVDCx5p33_ASAP7_75t_R g1424 ( .A(n_147), .Y(n_1424) );
INVx1_ASAP7_75t_L g854 ( .A(n_148), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_149), .A2(n_232), .B1(n_507), .B2(n_940), .Y(n_939) );
CKINVDCx5p33_ASAP7_75t_R g1485 ( .A(n_150), .Y(n_1485) );
OAI22xp33_ASAP7_75t_L g1500 ( .A1(n_151), .A2(n_204), .B1(n_462), .B2(n_1061), .Y(n_1500) );
OAI22xp33_ASAP7_75t_L g1506 ( .A1(n_151), .A2(n_191), .B1(n_532), .B2(n_535), .Y(n_1506) );
CKINVDCx5p33_ASAP7_75t_R g1478 ( .A(n_152), .Y(n_1478) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_153), .A2(n_171), .B1(n_739), .B2(n_741), .Y(n_1129) );
OAI22xp33_ASAP7_75t_L g1136 ( .A1(n_153), .A2(n_171), .B1(n_462), .B2(n_842), .Y(n_1136) );
OAI211xp5_ASAP7_75t_L g726 ( .A1(n_154), .A2(n_469), .B(n_474), .C(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g737 ( .A(n_154), .Y(n_737) );
CKINVDCx5p33_ASAP7_75t_R g1226 ( .A(n_155), .Y(n_1226) );
INVx1_ASAP7_75t_L g729 ( .A(n_156), .Y(n_729) );
OAI211xp5_ASAP7_75t_L g734 ( .A1(n_156), .A2(n_715), .B(n_735), .C(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g1025 ( .A(n_157), .Y(n_1025) );
INVx1_ASAP7_75t_L g860 ( .A(n_160), .Y(n_860) );
INVx1_ASAP7_75t_L g746 ( .A(n_161), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g1173 ( .A(n_162), .Y(n_1173) );
OAI211xp5_ASAP7_75t_L g704 ( .A1(n_163), .A2(n_471), .B(n_474), .C(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g718 ( .A(n_163), .Y(n_718) );
INVx1_ASAP7_75t_L g902 ( .A(n_164), .Y(n_902) );
AOI22xp33_ASAP7_75t_SL g1385 ( .A1(n_165), .A2(n_222), .B1(n_1386), .B2(n_1387), .Y(n_1385) );
INVx1_ASAP7_75t_L g706 ( .A(n_166), .Y(n_706) );
INVx1_ASAP7_75t_L g1860 ( .A(n_167), .Y(n_1860) );
OAI22xp33_ASAP7_75t_L g1465 ( .A1(n_168), .A2(n_292), .B1(n_596), .B2(n_842), .Y(n_1465) );
INVx1_ASAP7_75t_L g1498 ( .A(n_169), .Y(n_1498) );
OAI211xp5_ASAP7_75t_L g1503 ( .A1(n_169), .A2(n_715), .B(n_760), .C(n_1504), .Y(n_1503) );
CKINVDCx5p33_ASAP7_75t_R g1441 ( .A(n_170), .Y(n_1441) );
AO22x1_ASAP7_75t_L g1559 ( .A1(n_172), .A2(n_353), .B1(n_1518), .B2(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1321 ( .A(n_174), .Y(n_1321) );
CKINVDCx16_ASAP7_75t_R g1630 ( .A(n_175), .Y(n_1630) );
OAI211xp5_ASAP7_75t_SL g1103 ( .A1(n_176), .A2(n_474), .B(n_875), .C(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1116 ( .A(n_176), .Y(n_1116) );
INVx1_ASAP7_75t_L g592 ( .A(n_178), .Y(n_592) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_178), .A2(n_517), .B(n_650), .C(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g1359 ( .A(n_179), .Y(n_1359) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_180), .A2(n_309), .B1(n_489), .B2(n_491), .Y(n_708) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_180), .A2(n_309), .B1(n_530), .B2(n_720), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_181), .A2(n_281), .B1(n_1003), .B2(n_1004), .Y(n_1379) );
INVx1_ASAP7_75t_L g1143 ( .A(n_182), .Y(n_1143) );
OAI211xp5_ASAP7_75t_L g1495 ( .A1(n_183), .A2(n_697), .B(n_1196), .C(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1505 ( .A(n_183), .Y(n_1505) );
CKINVDCx5p33_ASAP7_75t_R g1177 ( .A(n_185), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g1363 ( .A(n_186), .Y(n_1363) );
INVx1_ASAP7_75t_L g756 ( .A(n_187), .Y(n_756) );
INVx1_ASAP7_75t_L g691 ( .A(n_188), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g1499 ( .A1(n_189), .A2(n_191), .B1(n_596), .B2(n_842), .Y(n_1499) );
OAI22xp33_ASAP7_75t_L g1502 ( .A1(n_189), .A2(n_204), .B1(n_505), .B2(n_1215), .Y(n_1502) );
INVx1_ASAP7_75t_L g1733 ( .A(n_190), .Y(n_1733) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_192), .A2(n_310), .B1(n_994), .B2(n_998), .Y(n_993) );
OAI211xp5_ASAP7_75t_L g1422 ( .A1(n_193), .A2(n_622), .B(n_715), .C(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g1431 ( .A(n_193), .Y(n_1431) );
INVx1_ASAP7_75t_L g610 ( .A(n_194), .Y(n_610) );
OAI22xp33_ASAP7_75t_SL g1203 ( .A1(n_195), .A2(n_322), .B1(n_462), .B2(n_490), .Y(n_1203) );
INVx1_ASAP7_75t_L g605 ( .A(n_196), .Y(n_605) );
INVx1_ASAP7_75t_L g665 ( .A(n_197), .Y(n_665) );
INVx2_ASAP7_75t_L g1521 ( .A(n_199), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_199), .B(n_316), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1529 ( .A(n_199), .B(n_1527), .Y(n_1529) );
AOI22xp33_ASAP7_75t_SL g1810 ( .A1(n_200), .A2(n_368), .B1(n_450), .B2(n_1811), .Y(n_1810) );
AO22x2_ASAP7_75t_L g1015 ( .A1(n_201), .A2(n_1016), .B1(n_1071), .B2(n_1072), .Y(n_1015) );
INVx1_ASAP7_75t_L g1071 ( .A(n_201), .Y(n_1071) );
INVx1_ASAP7_75t_L g621 ( .A(n_203), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g1482 ( .A(n_205), .Y(n_1482) );
CKINVDCx5p33_ASAP7_75t_R g1229 ( .A(n_206), .Y(n_1229) );
INVx1_ASAP7_75t_L g569 ( .A(n_207), .Y(n_569) );
XNOR2xp5_ASAP7_75t_L g1077 ( .A(n_208), .B(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g929 ( .A(n_209), .Y(n_929) );
OAI211xp5_ASAP7_75t_L g935 ( .A1(n_209), .A2(n_715), .B(n_936), .C(n_937), .Y(n_935) );
INVx1_ASAP7_75t_L g1278 ( .A(n_210), .Y(n_1278) );
XOR2xp5_ASAP7_75t_L g1310 ( .A(n_211), .B(n_1311), .Y(n_1310) );
INVxp67_ASAP7_75t_SL g1758 ( .A(n_212), .Y(n_1758) );
INVx1_ASAP7_75t_L g827 ( .A(n_213), .Y(n_827) );
OAI22xp33_ASAP7_75t_L g841 ( .A1(n_213), .A2(n_247), .B1(n_462), .B2(n_842), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_214), .A2(n_343), .B1(n_964), .B2(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_214), .A2(n_262), .B1(n_994), .B2(n_998), .Y(n_1001) );
XNOR2x2_ASAP7_75t_L g847 ( .A(n_215), .B(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g1316 ( .A(n_216), .Y(n_1316) );
NOR2xp33_ASAP7_75t_L g1763 ( .A(n_217), .B(n_1764), .Y(n_1763) );
INVx1_ASAP7_75t_L g1798 ( .A(n_217), .Y(n_1798) );
CKINVDCx5p33_ASAP7_75t_R g1447 ( .A(n_219), .Y(n_1447) );
INVx1_ASAP7_75t_L g480 ( .A(n_220), .Y(n_480) );
AOI22xp33_ASAP7_75t_SL g1395 ( .A1(n_222), .A2(n_300), .B1(n_411), .B2(n_1392), .Y(n_1395) );
INVx1_ASAP7_75t_L g1088 ( .A(n_223), .Y(n_1088) );
OAI211xp5_ASAP7_75t_L g1259 ( .A1(n_224), .A2(n_1260), .B(n_1261), .C(n_1270), .Y(n_1259) );
INVx1_ASAP7_75t_L g1299 ( .A(n_224), .Y(n_1299) );
INVx1_ASAP7_75t_L g676 ( .A(n_225), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_226), .A2(n_250), .B1(n_720), .B2(n_940), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_226), .A2(n_250), .B1(n_594), .B2(n_834), .Y(n_1135) );
INVx1_ASAP7_75t_L g1319 ( .A(n_227), .Y(n_1319) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_228), .A2(n_311), .B1(n_391), .B2(n_462), .Y(n_725) );
OAI22xp33_ASAP7_75t_L g738 ( .A1(n_228), .A2(n_311), .B1(n_739), .B2(n_741), .Y(n_738) );
INVx2_ASAP7_75t_L g440 ( .A(n_229), .Y(n_440) );
INVx1_ASAP7_75t_L g459 ( .A(n_229), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g1777 ( .A(n_229), .B(n_441), .Y(n_1777) );
CKINVDCx5p33_ASAP7_75t_R g1442 ( .A(n_230), .Y(n_1442) );
XNOR2xp5_ASAP7_75t_L g579 ( .A(n_231), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g794 ( .A(n_233), .Y(n_794) );
INVx1_ASAP7_75t_L g1411 ( .A(n_234), .Y(n_1411) );
XOR2xp5_ASAP7_75t_L g945 ( .A(n_235), .B(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g1269 ( .A(n_236), .Y(n_1269) );
OAI22xp5_ASAP7_75t_L g1297 ( .A1(n_236), .A2(n_267), .B1(n_532), .B2(n_535), .Y(n_1297) );
INVx1_ASAP7_75t_L g1262 ( .A(n_238), .Y(n_1262) );
INVx1_ASAP7_75t_L g819 ( .A(n_239), .Y(n_819) );
OA211x2_ASAP7_75t_L g835 ( .A1(n_239), .A2(n_633), .B(n_836), .C(n_837), .Y(n_835) );
BUFx3_ASAP7_75t_L g417 ( .A(n_240), .Y(n_417) );
INVx1_ASAP7_75t_L g1405 ( .A(n_241), .Y(n_1405) );
CKINVDCx5p33_ASAP7_75t_R g1452 ( .A(n_242), .Y(n_1452) );
OAI22xp33_ASAP7_75t_L g461 ( .A1(n_243), .A2(n_363), .B1(n_391), .B2(n_462), .Y(n_461) );
OAI22xp33_ASAP7_75t_L g502 ( .A1(n_243), .A2(n_363), .B1(n_503), .B2(n_507), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g1488 ( .A(n_244), .Y(n_1488) );
OAI22xp5_ASAP7_75t_SL g770 ( .A1(n_245), .A2(n_771), .B1(n_831), .B2(n_844), .Y(n_770) );
NAND4xp25_ASAP7_75t_L g771 ( .A(n_245), .B(n_772), .C(n_797), .D(n_812), .Y(n_771) );
XOR2xp5_ASAP7_75t_L g659 ( .A(n_246), .B(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g1556 ( .A1(n_246), .A2(n_252), .B1(n_1525), .B2(n_1528), .Y(n_1556) );
INVx1_ASAP7_75t_L g823 ( .A(n_247), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_248), .A2(n_262), .B1(n_964), .B2(n_968), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_248), .A2(n_343), .B1(n_986), .B2(n_990), .Y(n_985) );
INVx1_ASAP7_75t_L g484 ( .A(n_249), .Y(n_484) );
OAI211xp5_ASAP7_75t_L g510 ( .A1(n_249), .A2(n_511), .B(n_517), .C(n_519), .Y(n_510) );
OA22x2_ASAP7_75t_L g1119 ( .A1(n_251), .A2(n_1120), .B1(n_1159), .B2(n_1160), .Y(n_1119) );
INVxp67_ASAP7_75t_L g1160 ( .A(n_251), .Y(n_1160) );
INVx1_ASAP7_75t_L g1859 ( .A(n_253), .Y(n_1859) );
INVx1_ASAP7_75t_L g1274 ( .A(n_254), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_254), .B(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1056 ( .A(n_255), .Y(n_1056) );
INVx1_ASAP7_75t_L g669 ( .A(n_256), .Y(n_669) );
INVx1_ASAP7_75t_L g782 ( .A(n_257), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g1481 ( .A(n_258), .Y(n_1481) );
CKINVDCx5p33_ASAP7_75t_R g1444 ( .A(n_259), .Y(n_1444) );
INVx1_ASAP7_75t_L g749 ( .A(n_261), .Y(n_749) );
AOI221xp5_ASAP7_75t_L g1396 ( .A1(n_263), .A2(n_281), .B1(n_450), .B2(n_1397), .C(n_1398), .Y(n_1396) );
INVx1_ASAP7_75t_L g1020 ( .A(n_264), .Y(n_1020) );
INVx1_ASAP7_75t_L g1410 ( .A(n_265), .Y(n_1410) );
XOR2xp5_ASAP7_75t_L g1217 ( .A(n_266), .B(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1271 ( .A(n_267), .Y(n_1271) );
BUFx3_ASAP7_75t_L g399 ( .A(n_268), .Y(n_399) );
INVx1_ASAP7_75t_L g465 ( .A(n_268), .Y(n_465) );
INVx1_ASAP7_75t_L g879 ( .A(n_269), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g1632 ( .A(n_270), .Y(n_1632) );
AOI22xp5_ASAP7_75t_L g1532 ( .A1(n_272), .A2(n_290), .B1(n_1525), .B2(n_1528), .Y(n_1532) );
INVx1_ASAP7_75t_L g817 ( .A(n_274), .Y(n_817) );
INVx1_ASAP7_75t_L g1315 ( .A(n_275), .Y(n_1315) );
INVx1_ASAP7_75t_L g796 ( .A(n_276), .Y(n_796) );
XNOR2x1_ASAP7_75t_L g405 ( .A(n_278), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g863 ( .A(n_279), .Y(n_863) );
AOI21xp5_ASAP7_75t_L g1753 ( .A1(n_280), .A2(n_994), .B(n_1754), .Y(n_1753) );
INVx1_ASAP7_75t_L g423 ( .A(n_282), .Y(n_423) );
INVx1_ASAP7_75t_L g950 ( .A(n_283), .Y(n_950) );
OAI211xp5_ASAP7_75t_L g583 ( .A1(n_284), .A2(n_584), .B(n_585), .C(n_586), .Y(n_583) );
INVx1_ASAP7_75t_L g652 ( .A(n_284), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_286), .A2(n_367), .B1(n_425), .B2(n_430), .Y(n_424) );
INVxp33_ASAP7_75t_SL g549 ( .A(n_286), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g1175 ( .A(n_287), .Y(n_1175) );
NOR2xp33_ASAP7_75t_L g1249 ( .A(n_289), .B(n_535), .Y(n_1249) );
CKINVDCx5p33_ASAP7_75t_R g1233 ( .A(n_291), .Y(n_1233) );
OAI22xp33_ASAP7_75t_L g1468 ( .A1(n_292), .A2(n_313), .B1(n_505), .B2(n_1215), .Y(n_1468) );
CKINVDCx5p33_ASAP7_75t_R g1178 ( .A(n_293), .Y(n_1178) );
INVx1_ASAP7_75t_L g789 ( .A(n_294), .Y(n_789) );
XOR2x2_ASAP7_75t_L g722 ( .A(n_295), .B(n_723), .Y(n_722) );
CKINVDCx5p33_ASAP7_75t_R g1479 ( .A(n_296), .Y(n_1479) );
AOI22xp5_ASAP7_75t_L g1542 ( .A1(n_297), .A2(n_361), .B1(n_1525), .B2(n_1528), .Y(n_1542) );
AO22x1_ASAP7_75t_L g1517 ( .A1(n_298), .A2(n_304), .B1(n_1518), .B2(n_1522), .Y(n_1517) );
INVx1_ASAP7_75t_L g1857 ( .A(n_299), .Y(n_1857) );
INVx1_ASAP7_75t_L g415 ( .A(n_301), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_301), .Y(n_422) );
INVx1_ASAP7_75t_L g862 ( .A(n_302), .Y(n_862) );
INVx1_ASAP7_75t_L g856 ( .A(n_303), .Y(n_856) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_305), .A2(n_350), .B1(n_489), .B2(n_491), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_305), .A2(n_350), .B1(n_530), .B2(n_533), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_306), .A2(n_351), .B1(n_594), .B2(n_834), .Y(n_881) );
OAI22xp33_ASAP7_75t_L g889 ( .A1(n_306), .A2(n_351), .B1(n_654), .B2(n_720), .Y(n_889) );
INVx1_ASAP7_75t_L g785 ( .A(n_307), .Y(n_785) );
INVx1_ASAP7_75t_L g446 ( .A(n_308), .Y(n_446) );
INVx1_ASAP7_75t_L g1200 ( .A(n_312), .Y(n_1200) );
OAI211xp5_ASAP7_75t_SL g1206 ( .A1(n_312), .A2(n_517), .B(n_957), .C(n_1207), .Y(n_1206) );
INVx1_ASAP7_75t_L g1318 ( .A(n_314), .Y(n_1318) );
INVx1_ASAP7_75t_L g1368 ( .A(n_315), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_316), .B(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1527 ( .A(n_316), .Y(n_1527) );
OAI211xp5_ASAP7_75t_SL g1742 ( .A1(n_318), .A2(n_1743), .B(n_1747), .C(n_1755), .Y(n_1742) );
INVx1_ASAP7_75t_L g1795 ( .A(n_318), .Y(n_1795) );
INVx1_ASAP7_75t_L g1413 ( .A(n_320), .Y(n_1413) );
CKINVDCx5p33_ASAP7_75t_R g1445 ( .A(n_321), .Y(n_1445) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_322), .A2(n_358), .B1(n_532), .B2(n_535), .Y(n_1205) );
INVx1_ASAP7_75t_L g949 ( .A(n_323), .Y(n_949) );
CKINVDCx5p33_ASAP7_75t_R g1497 ( .A(n_324), .Y(n_1497) );
INVx1_ASAP7_75t_L g1037 ( .A(n_325), .Y(n_1037) );
CKINVDCx5p33_ASAP7_75t_R g1280 ( .A(n_326), .Y(n_1280) );
OAI211xp5_ASAP7_75t_SL g1243 ( .A1(n_327), .A2(n_567), .B(n_1196), .C(n_1244), .Y(n_1243) );
OAI211xp5_ASAP7_75t_SL g1251 ( .A1(n_327), .A2(n_517), .B(n_1252), .C(n_1253), .Y(n_1251) );
INVx1_ASAP7_75t_L g1408 ( .A(n_328), .Y(n_1408) );
INVx1_ASAP7_75t_L g1106 ( .A(n_329), .Y(n_1106) );
OAI211xp5_ASAP7_75t_SL g1112 ( .A1(n_329), .A2(n_517), .B(n_1113), .C(n_1115), .Y(n_1112) );
INVx1_ASAP7_75t_L g1337 ( .A(n_330), .Y(n_1337) );
INVx1_ASAP7_75t_L g447 ( .A(n_331), .Y(n_447) );
INVx1_ASAP7_75t_L g617 ( .A(n_332), .Y(n_617) );
OAI211xp5_ASAP7_75t_L g925 ( .A1(n_333), .A2(n_836), .B(n_926), .C(n_927), .Y(n_925) );
INVx1_ASAP7_75t_L g938 ( .A(n_333), .Y(n_938) );
AOI221xp5_ASAP7_75t_L g1759 ( .A1(n_335), .A2(n_368), .B1(n_1058), .B2(n_1760), .C(n_1762), .Y(n_1759) );
AOI22xp33_ASAP7_75t_SL g1846 ( .A1(n_336), .A2(n_373), .B1(n_1811), .B2(n_1847), .Y(n_1846) );
INVx1_ASAP7_75t_L g707 ( .A(n_337), .Y(n_707) );
OAI211xp5_ASAP7_75t_L g714 ( .A1(n_337), .A2(n_511), .B(n_715), .C(n_716), .Y(n_714) );
INVx1_ASAP7_75t_L g601 ( .A(n_338), .Y(n_601) );
INVx1_ASAP7_75t_L g1140 ( .A(n_339), .Y(n_1140) );
CKINVDCx5p33_ASAP7_75t_R g1181 ( .A(n_340), .Y(n_1181) );
INVx1_ASAP7_75t_L g776 ( .A(n_341), .Y(n_776) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_342), .Y(n_395) );
INVx1_ASAP7_75t_L g753 ( .A(n_344), .Y(n_753) );
INVx1_ASAP7_75t_L g1027 ( .A(n_345), .Y(n_1027) );
INVx1_ASAP7_75t_L g1781 ( .A(n_346), .Y(n_1781) );
INVx1_ASAP7_75t_L g682 ( .A(n_347), .Y(n_682) );
CKINVDCx5p33_ASAP7_75t_R g1463 ( .A(n_349), .Y(n_1463) );
CKINVDCx5p33_ASAP7_75t_R g1201 ( .A(n_354), .Y(n_1201) );
CKINVDCx5p33_ASAP7_75t_R g1225 ( .A(n_355), .Y(n_1225) );
INVx1_ASAP7_75t_L g1059 ( .A(n_357), .Y(n_1059) );
INVx1_ASAP7_75t_L g438 ( .A(n_359), .Y(n_438) );
INVx1_ASAP7_75t_L g458 ( .A(n_359), .Y(n_458) );
INVx2_ASAP7_75t_L g546 ( .A(n_359), .Y(n_546) );
INVx1_ASAP7_75t_L g898 ( .A(n_360), .Y(n_898) );
INVx1_ASAP7_75t_L g608 ( .A(n_364), .Y(n_608) );
INVx1_ASAP7_75t_L g1082 ( .A(n_365), .Y(n_1082) );
INVx1_ASAP7_75t_L g828 ( .A(n_366), .Y(n_828) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_367), .Y(n_566) );
INVx1_ASAP7_75t_L g1085 ( .A(n_369), .Y(n_1085) );
INVx1_ASAP7_75t_L g754 ( .A(n_370), .Y(n_754) );
AOI21xp33_ASAP7_75t_L g1281 ( .A1(n_371), .A2(n_1282), .B(n_1284), .Y(n_1281) );
INVx1_ASAP7_75t_L g1302 ( .A(n_371), .Y(n_1302) );
INVx1_ASAP7_75t_L g820 ( .A(n_372), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g1453 ( .A(n_374), .Y(n_1453) );
CKINVDCx5p33_ASAP7_75t_R g1267 ( .A(n_375), .Y(n_1267) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_400), .B(n_1509), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_385), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g1825 ( .A(n_379), .B(n_388), .Y(n_1825) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g1869 ( .A(n_381), .B(n_384), .Y(n_1869) );
INVx1_ASAP7_75t_L g1871 ( .A(n_381), .Y(n_1871) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g1873 ( .A(n_384), .B(n_1871), .Y(n_1873) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g498 ( .A(n_388), .B(n_499), .Y(n_498) );
AOI21xp5_ASAP7_75t_SL g1258 ( .A1(n_388), .A2(n_1259), .B(n_1272), .Y(n_1258) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g576 ( .A(n_389), .B(n_399), .Y(n_576) );
AND2x4_ASAP7_75t_L g1285 ( .A(n_389), .B(n_398), .Y(n_1285) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_390), .A2(n_463), .B1(n_949), .B2(n_950), .Y(n_1007) );
AND2x4_ASAP7_75t_SL g1824 ( .A(n_390), .B(n_1825), .Y(n_1824) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_397), .Y(n_391) );
OR2x6_ASAP7_75t_L g490 ( .A(n_392), .B(n_464), .Y(n_490) );
BUFx4f_ASAP7_75t_L g550 ( .A(n_392), .Y(n_550) );
OR2x2_ASAP7_75t_L g1061 ( .A(n_392), .B(n_464), .Y(n_1061) );
INVx1_ASAP7_75t_L g1192 ( .A(n_392), .Y(n_1192) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g572 ( .A(n_393), .Y(n_572) );
BUFx4f_ASAP7_75t_L g630 ( .A(n_393), .Y(n_630) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
AND2x2_ASAP7_75t_L g466 ( .A(n_395), .B(n_467), .Y(n_466) );
NAND2x1_ASAP7_75t_L g473 ( .A(n_395), .B(n_396), .Y(n_473) );
AND2x2_ASAP7_75t_L g478 ( .A(n_395), .B(n_396), .Y(n_478) );
INVx1_ASAP7_75t_L g487 ( .A(n_395), .Y(n_487) );
INVx2_ASAP7_75t_L g496 ( .A(n_395), .Y(n_496) );
INVx2_ASAP7_75t_L g560 ( .A(n_395), .Y(n_560) );
INVx2_ASAP7_75t_L g467 ( .A(n_396), .Y(n_467) );
BUFx2_ASAP7_75t_L g483 ( .A(n_396), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_396), .B(n_496), .Y(n_495) );
OR2x2_ASAP7_75t_L g559 ( .A(n_396), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g989 ( .A(n_396), .Y(n_989) );
AND2x2_ASAP7_75t_L g992 ( .A(n_396), .B(n_496), .Y(n_992) );
OR2x6_ASAP7_75t_L g842 ( .A(n_397), .B(n_572), .Y(n_842) );
AOI22xp5_ASAP7_75t_L g1266 ( .A1(n_397), .A2(n_1267), .B1(n_1268), .B2(n_1269), .Y(n_1266) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g476 ( .A(n_398), .Y(n_476) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g482 ( .A(n_399), .Y(n_482) );
AND2x4_ASAP7_75t_L g485 ( .A(n_399), .B(n_486), .Y(n_485) );
XNOR2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_942), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_845), .B2(n_941), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
XOR2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_656), .Y(n_403) );
XNOR2x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_579), .Y(n_404) );
NAND4xp75_ASAP7_75t_L g406 ( .A(n_407), .B(n_460), .C(n_501), .D(n_541), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_433), .B1(n_442), .B2(n_453), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_418), .B1(n_419), .B2(n_423), .C(n_424), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_410), .A2(n_419), .B1(n_902), .B2(n_911), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g1157 ( .A1(n_410), .A2(n_419), .B1(n_1144), .B2(n_1152), .Y(n_1157) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g1448 ( .A(n_411), .Y(n_1448) );
INVx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g781 ( .A(n_412), .Y(n_781) );
INVx1_ASAP7_75t_L g980 ( .A(n_412), .Y(n_980) );
BUFx2_ASAP7_75t_L g1307 ( .A(n_412), .Y(n_1307) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_413), .Y(n_445) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_413), .Y(n_616) );
BUFx8_ASAP7_75t_L g788 ( .A(n_413), .Y(n_788) );
AND2x4_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g429 ( .A(n_415), .Y(n_429) );
AND2x4_ASAP7_75t_L g427 ( .A(n_416), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_417), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g431 ( .A(n_417), .B(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g506 ( .A(n_417), .B(n_429), .Y(n_506) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_417), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_418), .A2(n_446), .B1(n_556), .B2(n_561), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g442 ( .A1(n_419), .A2(n_443), .B1(n_446), .B2(n_447), .C(n_448), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_419), .A2(n_608), .B1(n_609), .B2(n_610), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_419), .A2(n_612), .B1(n_613), .B2(n_617), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_419), .A2(n_763), .B1(n_857), .B2(n_863), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_419), .A2(n_1085), .B1(n_1091), .B2(n_1097), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1099 ( .A1(n_419), .A2(n_1086), .B1(n_1092), .B2(n_1100), .Y(n_1099) );
BUFx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OR2x6_ASAP7_75t_L g532 ( .A(n_420), .B(n_456), .Y(n_532) );
INVx1_ASAP7_75t_L g679 ( .A(n_420), .Y(n_679) );
BUFx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g685 ( .A(n_421), .Y(n_685) );
INVx2_ASAP7_75t_L g432 ( .A(n_422), .Y(n_432) );
INVx1_ASAP7_75t_L g515 ( .A(n_422), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_423), .A2(n_447), .B1(n_571), .B2(n_573), .Y(n_570) );
BUFx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g1848 ( .A(n_426), .Y(n_1848) );
BUFx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx8_ASAP7_75t_L g451 ( .A(n_427), .Y(n_451) );
BUFx3_ASAP7_75t_L g967 ( .A(n_427), .Y(n_967) );
NAND2x1p5_ASAP7_75t_L g1788 ( .A(n_427), .B(n_1789), .Y(n_1788) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI222xp33_ASAP7_75t_L g1335 ( .A1(n_430), .A2(n_818), .B1(n_1212), .B2(n_1336), .C1(n_1337), .C2(n_1338), .Y(n_1335) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g452 ( .A(n_431), .Y(n_452) );
AND2x4_ASAP7_75t_L g518 ( .A(n_431), .B(n_456), .Y(n_518) );
BUFx2_ASAP7_75t_L g821 ( .A(n_431), .Y(n_821) );
INVx2_ASAP7_75t_L g969 ( .A(n_431), .Y(n_969) );
BUFx2_ASAP7_75t_L g978 ( .A(n_431), .Y(n_978) );
BUFx3_ASAP7_75t_L g1397 ( .A(n_431), .Y(n_1397) );
INVx1_ASAP7_75t_L g975 ( .A(n_432), .Y(n_975) );
BUFx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI33xp33_ASAP7_75t_L g599 ( .A1(n_434), .A2(n_600), .A3(n_607), .B1(n_611), .B2(n_618), .B3(n_619), .Y(n_599) );
OAI33xp33_ASAP7_75t_L g1168 ( .A1(n_434), .A2(n_1169), .A3(n_1172), .B1(n_1176), .B2(n_1179), .B3(n_1182), .Y(n_1168) );
OAI33xp33_ASAP7_75t_L g1220 ( .A1(n_434), .A2(n_1182), .A3(n_1221), .B1(n_1224), .B2(n_1228), .B3(n_1232), .Y(n_1220) );
OAI33xp33_ASAP7_75t_L g1402 ( .A1(n_434), .A2(n_1182), .A3(n_1403), .B1(n_1406), .B2(n_1409), .B3(n_1412), .Y(n_1402) );
OAI33xp33_ASAP7_75t_L g1439 ( .A1(n_434), .A2(n_1182), .A3(n_1440), .B1(n_1443), .B2(n_1446), .B3(n_1450), .Y(n_1439) );
OAI33xp33_ASAP7_75t_L g1489 ( .A1(n_434), .A2(n_1182), .A3(n_1490), .B1(n_1491), .B2(n_1492), .B3(n_1493), .Y(n_1489) );
BUFx4f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx4f_ASAP7_75t_L g663 ( .A(n_435), .Y(n_663) );
BUFx2_ASAP7_75t_L g774 ( .A(n_435), .Y(n_774) );
BUFx8_ASAP7_75t_L g915 ( .A(n_435), .Y(n_915) );
OR2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_439), .Y(n_435) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_436), .Y(n_540) );
INVx1_ASAP7_75t_L g578 ( .A(n_436), .Y(n_578) );
AND2x2_ASAP7_75t_SL g809 ( .A(n_436), .B(n_576), .Y(n_809) );
OR2x2_ASAP7_75t_L g1776 ( .A(n_436), .B(n_1777), .Y(n_1776) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g500 ( .A(n_437), .Y(n_500) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND2xp33_ASAP7_75t_SL g439 ( .A(n_440), .B(n_441), .Y(n_439) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_440), .Y(n_538) );
AND3x4_ASAP7_75t_L g961 ( .A(n_440), .B(n_523), .C(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g1790 ( .A(n_440), .Y(n_1790) );
INVx3_ASAP7_75t_L g456 ( .A(n_441), .Y(n_456) );
BUFx3_ASAP7_75t_L g523 ( .A(n_441), .Y(n_523) );
OAI22xp33_ASAP7_75t_L g1156 ( .A1(n_443), .A2(n_683), .B1(n_1143), .B2(n_1151), .Y(n_1156) );
OAI211xp5_ASAP7_75t_L g1301 ( .A1(n_443), .A2(n_1302), .B(n_1303), .C(n_1304), .Y(n_1301) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g508 ( .A(n_445), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g609 ( .A(n_445), .Y(n_609) );
AND2x2_ASAP7_75t_L g824 ( .A(n_445), .B(n_509), .Y(n_824) );
INVx2_ASAP7_75t_L g921 ( .A(n_445), .Y(n_921) );
BUFx6f_ASAP7_75t_L g1098 ( .A(n_445), .Y(n_1098) );
INVx2_ASAP7_75t_L g1100 ( .A(n_445), .Y(n_1100) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx8_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g1309 ( .A(n_451), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_452), .B(n_1056), .Y(n_1068) );
OAI33xp33_ASAP7_75t_L g914 ( .A1(n_453), .A2(n_915), .A3(n_916), .B1(n_919), .B2(n_920), .B3(n_922), .Y(n_914) );
OAI33xp33_ASAP7_75t_L g1153 ( .A1(n_453), .A2(n_774), .A3(n_1154), .B1(n_1156), .B2(n_1157), .B3(n_1158), .Y(n_1153) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g618 ( .A(n_454), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_454), .Y(n_765) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx3_ASAP7_75t_L g689 ( .A(n_455), .Y(n_689) );
NAND3x1_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .C(n_459), .Y(n_455) );
OR2x4_ASAP7_75t_L g505 ( .A(n_456), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g509 ( .A(n_456), .Y(n_509) );
NAND2x1p5_ASAP7_75t_L g792 ( .A(n_456), .B(n_459), .Y(n_792) );
AND2x4_ASAP7_75t_L g1789 ( .A(n_456), .B(n_1790), .Y(n_1789) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g1779 ( .A(n_458), .Y(n_1779) );
OAI31xp33_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_468), .A3(n_488), .B(n_497), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_463), .Y(n_462) );
INVx4_ASAP7_75t_L g873 ( .A(n_463), .Y(n_873) );
INVx3_ASAP7_75t_SL g1260 ( .A(n_463), .Y(n_1260) );
AOI22xp5_ASAP7_75t_L g1356 ( .A1(n_463), .A2(n_1357), .B1(n_1358), .B2(n_1359), .Y(n_1356) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g997 ( .A(n_466), .Y(n_997) );
BUFx6f_ASAP7_75t_L g1283 ( .A(n_466), .Y(n_1283) );
BUFx3_ASAP7_75t_L g1836 ( .A(n_466), .Y(n_1836) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g584 ( .A(n_471), .Y(n_584) );
BUFx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_SL g561 ( .A(n_472), .Y(n_561) );
INVx2_ASAP7_75t_SL g634 ( .A(n_472), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_472), .A2(n_638), .B1(n_856), .B2(n_857), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g1458 ( .A1(n_472), .A2(n_805), .B1(n_1442), .B2(n_1453), .Y(n_1458) );
OAI22xp5_ASAP7_75t_L g1480 ( .A1(n_472), .A2(n_1457), .B1(n_1481), .B2(n_1482), .Y(n_1480) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_473), .Y(n_568) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g585 ( .A(n_475), .Y(n_585) );
INVx3_ASAP7_75t_L g836 ( .A(n_475), .Y(n_836) );
NOR3xp33_ASAP7_75t_L g1008 ( .A(n_475), .B(n_1009), .C(n_1012), .Y(n_1008) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_476), .B(n_1198), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_476), .B(n_494), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_476), .B(n_483), .Y(n_1265) );
BUFx3_ASAP7_75t_L g1058 ( .A(n_477), .Y(n_1058) );
AND2x6_ASAP7_75t_L g1734 ( .A(n_477), .B(n_1735), .Y(n_1734) );
AND2x4_ASAP7_75t_SL g1767 ( .A(n_477), .B(n_1732), .Y(n_1767) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g1000 ( .A(n_478), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_484), .B2(n_485), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_480), .A2(n_520), .B1(n_525), .B2(n_528), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_481), .A2(n_1054), .B1(n_1055), .B2(n_1056), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_481), .A2(n_1127), .B1(n_1133), .B2(n_1134), .Y(n_1132) );
AOI22xp5_ASAP7_75t_L g1199 ( .A1(n_481), .A2(n_590), .B1(n_1200), .B2(n_1201), .Y(n_1199) );
AOI222xp33_ASAP7_75t_L g1342 ( .A1(n_481), .A2(n_1055), .B1(n_1058), .B2(n_1337), .C1(n_1338), .C2(n_1343), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_481), .A2(n_590), .B1(n_1424), .B2(n_1431), .Y(n_1430) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
OR2x2_ASAP7_75t_L g493 ( .A(n_482), .B(n_494), .Y(n_493) );
AND2x4_ASAP7_75t_L g588 ( .A(n_482), .B(n_483), .Y(n_588) );
O2A1O1Ixp33_ASAP7_75t_L g1261 ( .A1(n_482), .A2(n_1058), .B(n_1262), .C(n_1263), .Y(n_1261) );
INVx1_ASAP7_75t_L g1268 ( .A(n_482), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_482), .B(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g1745 ( .A(n_483), .Y(n_1745) );
INVx2_ASAP7_75t_L g591 ( .A(n_485), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_485), .A2(n_588), .B1(n_728), .B2(n_729), .Y(n_727) );
INVx2_ASAP7_75t_L g839 ( .A(n_485), .Y(n_839) );
BUFx3_ASAP7_75t_L g1055 ( .A(n_485), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_485), .A2(n_1265), .B1(n_1363), .B2(n_1364), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1785 ( .A(n_486), .B(n_1735), .Y(n_1785) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_490), .Y(n_594) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g834 ( .A(n_492), .Y(n_834) );
INVxp67_ASAP7_75t_SL g931 ( .A(n_492), .Y(n_931) );
INVx1_ASAP7_75t_L g1062 ( .A(n_492), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1855 ( .A1(n_492), .A2(n_1346), .B1(n_1856), .B2(n_1857), .Y(n_1855) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g596 ( .A(n_493), .Y(n_596) );
INVx1_ASAP7_75t_L g1011 ( .A(n_493), .Y(n_1011) );
INVx8_ASAP7_75t_L g554 ( .A(n_494), .Y(n_554) );
BUFx2_ASAP7_75t_L g803 ( .A(n_494), .Y(n_803) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g843 ( .A(n_497), .Y(n_843) );
OAI31xp33_ASAP7_75t_L g924 ( .A1(n_497), .A2(n_925), .A3(n_930), .B(n_932), .Y(n_924) );
OAI31xp33_ASAP7_75t_L g1050 ( .A1(n_497), .A2(n_1051), .A3(n_1052), .B(n_1060), .Y(n_1050) );
OAI31xp33_ASAP7_75t_L g1194 ( .A1(n_497), .A2(n_1195), .A3(n_1202), .B(n_1203), .Y(n_1194) );
OAI31xp33_ASAP7_75t_SL g1427 ( .A1(n_497), .A2(n_1428), .A3(n_1429), .B(n_1432), .Y(n_1427) );
OAI31xp33_ASAP7_75t_L g1460 ( .A1(n_497), .A2(n_1461), .A3(n_1465), .B(n_1466), .Y(n_1460) );
OAI31xp33_ASAP7_75t_L g1494 ( .A1(n_497), .A2(n_1495), .A3(n_1499), .B(n_1500), .Y(n_1494) );
BUFx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx3_ASAP7_75t_L g597 ( .A(n_498), .Y(n_597) );
BUFx2_ASAP7_75t_SL g731 ( .A(n_498), .Y(n_731) );
INVx1_ASAP7_75t_L g1014 ( .A(n_498), .Y(n_1014) );
OAI31xp33_ASAP7_75t_L g1240 ( .A1(n_498), .A2(n_1241), .A3(n_1243), .B(n_1247), .Y(n_1240) );
OAI21xp5_ASAP7_75t_L g1340 ( .A1(n_498), .A2(n_1341), .B(n_1350), .Y(n_1340) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g1784 ( .A(n_500), .B(n_1785), .Y(n_1784) );
INVxp67_ASAP7_75t_L g1791 ( .A(n_500), .Y(n_1791) );
OAI31xp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_510), .A3(n_529), .B(n_536), .Y(n_501) );
INVx2_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_504), .A2(n_508), .B1(n_949), .B2(n_950), .Y(n_948) );
AOI22xp5_ASAP7_75t_L g1371 ( .A1(n_504), .A2(n_824), .B1(n_1357), .B2(n_1359), .Y(n_1371) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g648 ( .A(n_505), .Y(n_648) );
INVx1_ASAP7_75t_L g713 ( .A(n_505), .Y(n_713) );
INVx1_ASAP7_75t_L g740 ( .A(n_505), .Y(n_740) );
OR2x4_ASAP7_75t_L g535 ( .A(n_506), .B(n_509), .Y(n_535) );
BUFx3_ASAP7_75t_L g604 ( .A(n_506), .Y(n_604) );
BUFx3_ASAP7_75t_L g620 ( .A(n_506), .Y(n_620) );
INVx2_ASAP7_75t_L g668 ( .A(n_506), .Y(n_668) );
BUFx4f_ASAP7_75t_L g1042 ( .A(n_506), .Y(n_1042) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g741 ( .A(n_508), .Y(n_741) );
INVx1_ASAP7_75t_L g884 ( .A(n_508), .Y(n_884) );
INVx1_ASAP7_75t_L g1065 ( .A(n_508), .Y(n_1065) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_511), .Y(n_735) );
OAI22xp33_ASAP7_75t_L g766 ( .A1(n_511), .A2(n_666), .B1(n_746), .B2(n_754), .Y(n_766) );
OAI22xp33_ASAP7_75t_L g916 ( .A1(n_511), .A2(n_898), .B1(n_908), .B2(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g606 ( .A(n_512), .Y(n_606) );
INVx2_ASAP7_75t_L g650 ( .A(n_512), .Y(n_650) );
INVx1_ASAP7_75t_L g936 ( .A(n_512), .Y(n_936) );
INVx2_ASAP7_75t_L g1294 ( .A(n_512), .Y(n_1294) );
INVx4_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g778 ( .A(n_513), .Y(n_778) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_513), .Y(n_795) );
HB1xp67_ASAP7_75t_L g1095 ( .A(n_513), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1786 ( .A(n_513), .B(n_1776), .Y(n_1786) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx3_ASAP7_75t_L g623 ( .A(n_514), .Y(n_623) );
BUFx2_ASAP7_75t_L g672 ( .A(n_514), .Y(n_672) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
BUFx2_ASAP7_75t_L g527 ( .A(n_515), .Y(n_527) );
BUFx2_ASAP7_75t_L g524 ( .A(n_516), .Y(n_524) );
AND2x4_ASAP7_75t_L g974 ( .A(n_516), .B(n_975), .Y(n_974) );
INVx2_ASAP7_75t_L g1211 ( .A(n_516), .Y(n_1211) );
NAND3xp33_ASAP7_75t_L g1066 ( .A(n_517), .B(n_1067), .C(n_1068), .Y(n_1066) );
NAND3xp33_ASAP7_75t_L g1865 ( .A(n_517), .B(n_1866), .C(n_1867), .Y(n_1865) );
CKINVDCx8_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
CKINVDCx8_ASAP7_75t_R g715 ( .A(n_518), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_518), .B(n_815), .Y(n_814) );
NOR3xp33_ASAP7_75t_L g951 ( .A(n_518), .B(n_952), .C(n_956), .Y(n_951) );
NOR3xp33_ASAP7_75t_L g1292 ( .A(n_518), .B(n_1293), .C(n_1297), .Y(n_1292) );
NOR3xp33_ASAP7_75t_L g1372 ( .A(n_518), .B(n_1373), .C(n_1376), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_520), .A2(n_525), .B1(n_589), .B2(n_652), .Y(n_651) );
AOI222xp33_ASAP7_75t_L g1866 ( .A1(n_520), .A2(n_526), .B1(n_821), .B2(n_1859), .C1(n_1860), .C2(n_1861), .Y(n_1866) );
BUFx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx3_ASAP7_75t_L g887 ( .A(n_521), .Y(n_887) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_524), .Y(n_521) );
AND2x4_ASAP7_75t_L g526 ( .A(n_522), .B(n_527), .Y(n_526) );
AND2x4_ASAP7_75t_L g717 ( .A(n_522), .B(n_524), .Y(n_717) );
AND2x4_ASAP7_75t_L g818 ( .A(n_522), .B(n_524), .Y(n_818) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_522), .B(n_527), .Y(n_1212) );
INVx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_523), .B(n_1209), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_525), .A2(n_879), .B1(n_887), .B2(n_888), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_525), .A2(n_887), .B1(n_1105), .B2(n_1116), .Y(n_1115) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g716 ( .A1(n_526), .A2(n_706), .B1(n_717), .B2(n_718), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_526), .A2(n_717), .B1(n_728), .B2(n_737), .Y(n_736) );
AOI222xp33_ASAP7_75t_L g816 ( .A1(n_526), .A2(n_817), .B1(n_818), .B2(n_819), .C1(n_820), .C2(n_821), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_526), .A2(n_717), .B1(n_928), .B2(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g958 ( .A(n_526), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_526), .A2(n_717), .B1(n_1054), .B2(n_1059), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_526), .A2(n_717), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g655 ( .A(n_532), .Y(n_655) );
BUFx3_ASAP7_75t_L g940 ( .A(n_532), .Y(n_940) );
INVx2_ASAP7_75t_L g955 ( .A(n_532), .Y(n_955) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_534), .A2(n_713), .B1(n_827), .B2(n_828), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g1867 ( .A1(n_534), .A2(n_955), .B1(n_1856), .B2(n_1857), .Y(n_1867) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g720 ( .A(n_535), .Y(n_720) );
BUFx2_ASAP7_75t_L g953 ( .A(n_535), .Y(n_953) );
BUFx2_ASAP7_75t_L g1111 ( .A(n_535), .Y(n_1111) );
OAI31xp33_ASAP7_75t_L g645 ( .A1(n_536), .A2(n_646), .A3(n_649), .B(n_653), .Y(n_645) );
BUFx2_ASAP7_75t_L g890 ( .A(n_536), .Y(n_890) );
AOI21xp5_ASAP7_75t_L g1290 ( .A1(n_536), .A2(n_1291), .B(n_1300), .Y(n_1290) );
AND2x2_ASAP7_75t_SL g536 ( .A(n_537), .B(n_539), .Y(n_536) );
AND2x2_ASAP7_75t_L g721 ( .A(n_537), .B(n_539), .Y(n_721) );
AND2x4_ASAP7_75t_L g830 ( .A(n_537), .B(n_539), .Y(n_830) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_537), .B(n_539), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_537), .B(n_539), .Y(n_1216) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OA33x2_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_548), .A3(n_555), .B1(n_562), .B2(n_570), .B3(n_574), .Y(n_541) );
OAI33xp33_ASAP7_75t_L g693 ( .A1(n_542), .A2(n_644), .A3(n_694), .B1(n_695), .B2(n_699), .B3(n_701), .Y(n_693) );
OAI33xp33_ASAP7_75t_L g743 ( .A1(n_542), .A2(n_574), .A3(n_744), .B1(n_747), .B2(n_750), .B3(n_755), .Y(n_743) );
INVx1_ASAP7_75t_L g984 ( .A(n_542), .Y(n_984) );
OAI33xp33_ASAP7_75t_L g1080 ( .A1(n_542), .A2(n_644), .A3(n_1081), .B1(n_1084), .B2(n_1087), .B3(n_1090), .Y(n_1080) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OAI33xp33_ASAP7_75t_L g625 ( .A1(n_543), .A2(n_626), .A3(n_632), .B1(n_635), .B2(n_639), .B3(n_644), .Y(n_625) );
OAI33xp33_ASAP7_75t_L g1235 ( .A1(n_543), .A2(n_1193), .A3(n_1236), .B1(n_1237), .B2(n_1238), .B3(n_1239), .Y(n_1235) );
OAI33xp33_ASAP7_75t_L g1476 ( .A1(n_543), .A2(n_808), .A3(n_1477), .B1(n_1480), .B2(n_1483), .B3(n_1486), .Y(n_1476) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g801 ( .A(n_544), .Y(n_801) );
INVx2_ASAP7_75t_L g851 ( .A(n_544), .Y(n_851) );
INVx2_ASAP7_75t_L g1184 ( .A(n_544), .Y(n_1184) );
AND2x4_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .Y(n_544) );
OR2x6_ASAP7_75t_L g791 ( .A(n_545), .B(n_792), .Y(n_791) );
OR2x2_ASAP7_75t_L g1182 ( .A(n_545), .B(n_792), .Y(n_1182) );
INVx1_ASAP7_75t_L g1289 ( .A(n_545), .Y(n_1289) );
BUFx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g962 ( .A(n_546), .Y(n_962) );
OAI22xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B1(n_551), .B2(n_552), .Y(n_548) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_550), .A2(n_552), .B1(n_665), .B2(n_691), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_550), .A2(n_552), .B1(n_745), .B2(n_746), .Y(n_744) );
OAI22xp33_ASAP7_75t_L g802 ( .A1(n_550), .A2(n_776), .B1(n_794), .B2(n_803), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_550), .A2(n_785), .B1(n_790), .B2(n_811), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g1273 ( .A1(n_550), .A2(n_552), .B1(n_1274), .B2(n_1275), .Y(n_1273) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_552), .A2(n_676), .B1(n_686), .B2(n_702), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_552), .A2(n_702), .B1(n_756), .B2(n_757), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g1139 ( .A1(n_552), .A2(n_899), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_552), .A2(n_1149), .B1(n_1151), .B2(n_1152), .Y(n_1148) );
INVx5_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx6_ASAP7_75t_L g573 ( .A(n_553), .Y(n_573) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g631 ( .A(n_554), .Y(n_631) );
INVx1_ASAP7_75t_L g643 ( .A(n_554), .Y(n_643) );
INVx2_ASAP7_75t_SL g811 ( .A(n_554), .Y(n_811) );
INVx2_ASAP7_75t_L g912 ( .A(n_554), .Y(n_912) );
INVx2_ASAP7_75t_L g1034 ( .A(n_554), .Y(n_1034) );
INVx4_ASAP7_75t_L g1186 ( .A(n_554), .Y(n_1186) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_556), .A2(n_608), .B1(n_612), .B2(n_633), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g858 ( .A1(n_556), .A2(n_561), .B1(n_859), .B2(n_860), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_556), .A2(n_633), .B1(n_1085), .B2(n_1086), .Y(n_1084) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx4_ASAP7_75t_L g696 ( .A(n_557), .Y(n_696) );
INVx2_ASAP7_75t_L g903 ( .A(n_557), .Y(n_903) );
INVx4_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g565 ( .A(n_559), .Y(n_565) );
BUFx3_ASAP7_75t_L g752 ( .A(n_559), .Y(n_752) );
BUFx2_ASAP7_75t_L g805 ( .A(n_559), .Y(n_805) );
INVx1_ASAP7_75t_L g907 ( .A(n_559), .Y(n_907) );
AND2x2_ASAP7_75t_L g988 ( .A(n_560), .B(n_989), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_561), .A2(n_636), .B1(n_1088), .B2(n_1089), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_566), .B1(n_567), .B2(n_569), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_563), .A2(n_779), .B1(n_796), .B2(n_806), .Y(n_807) );
OAI221xp5_ASAP7_75t_L g1276 ( .A1(n_563), .A2(n_576), .B1(n_806), .B2(n_1277), .C(n_1278), .Y(n_1276) );
INVx4_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g638 ( .A(n_565), .Y(n_638) );
INVx2_ASAP7_75t_L g1457 ( .A(n_565), .Y(n_1457) );
OAI22xp5_ASAP7_75t_L g1329 ( .A1(n_567), .A2(n_752), .B1(n_1318), .B2(n_1321), .Y(n_1329) );
BUFx4f_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx4_ASAP7_75t_L g698 ( .A(n_568), .Y(n_698) );
BUFx4f_ASAP7_75t_L g700 ( .A(n_568), .Y(n_700) );
BUFx4f_ASAP7_75t_L g877 ( .A(n_568), .Y(n_877) );
BUFx6f_ASAP7_75t_L g1023 ( .A(n_568), .Y(n_1023) );
BUFx4f_ASAP7_75t_L g1038 ( .A(n_568), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_571), .A2(n_573), .B1(n_862), .B2(n_863), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_571), .A2(n_911), .B1(n_912), .B2(n_913), .Y(n_910) );
OAI22xp33_ASAP7_75t_L g1081 ( .A1(n_571), .A2(n_573), .B1(n_1082), .B2(n_1083), .Y(n_1081) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_571), .A2(n_642), .B1(n_1091), .B2(n_1092), .Y(n_1090) );
BUFx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx3_ASAP7_75t_L g1032 ( .A(n_572), .Y(n_1032) );
INVx2_ASAP7_75t_SL g1150 ( .A(n_572), .Y(n_1150) );
BUFx6f_ASAP7_75t_L g1332 ( .A(n_572), .Y(n_1332) );
OAI22xp5_ASAP7_75t_SL g852 ( .A1(n_573), .A2(n_629), .B1(n_853), .B2(n_854), .Y(n_852) );
OAI33xp33_ASAP7_75t_L g896 ( .A1(n_574), .A2(n_801), .A3(n_897), .B1(n_901), .B2(n_905), .B3(n_910), .Y(n_896) );
OAI33xp33_ASAP7_75t_L g1138 ( .A1(n_574), .A2(n_851), .A3(n_1139), .B1(n_1142), .B2(n_1145), .B3(n_1148), .Y(n_1138) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g644 ( .A(n_575), .Y(n_644) );
AOI33xp33_ASAP7_75t_L g983 ( .A1(n_575), .A2(n_984), .A3(n_985), .B1(n_993), .B2(n_1001), .B3(n_1002), .Y(n_983) );
AND2x4_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx4_ASAP7_75t_L g1762 ( .A(n_576), .Y(n_1762) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND3x1_ASAP7_75t_L g580 ( .A(n_581), .B(n_598), .C(n_645), .Y(n_580) );
OAI31xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .A3(n_593), .B(n_597), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_589), .B1(n_590), .B2(n_592), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_587), .A2(n_838), .B1(n_879), .B2(n_880), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_587), .A2(n_1055), .B1(n_1105), .B2(n_1106), .Y(n_1104) );
BUFx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_588), .A2(n_590), .B1(n_706), .B2(n_707), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_588), .A2(n_817), .B1(n_820), .B2(n_838), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_588), .A2(n_590), .B1(n_928), .B2(n_929), .Y(n_927) );
INVx1_ASAP7_75t_L g1013 ( .A(n_588), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g1244 ( .A1(n_588), .A2(n_1055), .B1(n_1245), .B2(n_1246), .Y(n_1244) );
AOI222xp33_ASAP7_75t_L g1858 ( .A1(n_588), .A2(n_1055), .B1(n_1058), .B2(n_1859), .C1(n_1860), .C2(n_1861), .Y(n_1858) );
AOI22xp5_ASAP7_75t_L g1462 ( .A1(n_590), .A2(n_1265), .B1(n_1463), .B2(n_1464), .Y(n_1462) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OAI31xp33_ASAP7_75t_SL g703 ( .A1(n_597), .A2(n_704), .A3(n_708), .B(n_709), .Y(n_703) );
OAI31xp33_ASAP7_75t_L g871 ( .A1(n_597), .A2(n_872), .A3(n_874), .B(n_881), .Y(n_871) );
OAI31xp33_ASAP7_75t_L g1102 ( .A1(n_597), .A2(n_1103), .A3(n_1107), .B(n_1108), .Y(n_1102) );
NOR2xp33_ASAP7_75t_SL g598 ( .A(n_599), .B(n_625), .Y(n_598) );
OAI22xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_605), .B2(n_606), .Y(n_600) );
OAI22xp33_ASAP7_75t_L g626 ( .A1(n_601), .A2(n_621), .B1(n_627), .B2(n_631), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g865 ( .A1(n_602), .A2(n_853), .B1(n_859), .B2(n_866), .Y(n_865) );
OAI22xp33_ASAP7_75t_L g870 ( .A1(n_602), .A2(n_760), .B1(n_854), .B2(n_860), .Y(n_870) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVxp67_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g918 ( .A(n_604), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_605), .A2(n_624), .B1(n_633), .B2(n_636), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g1224 ( .A1(n_609), .A2(n_1225), .B1(n_1226), .B2(n_1227), .Y(n_1224) );
OAI22xp5_ASAP7_75t_L g1443 ( .A1(n_609), .A2(n_1227), .B1(n_1444), .B2(n_1445), .Y(n_1443) );
OAI22xp5_ASAP7_75t_L g1491 ( .A1(n_609), .A2(n_1227), .B1(n_1481), .B2(n_1487), .Y(n_1491) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_610), .A2(n_617), .B1(n_640), .B2(n_642), .Y(n_639) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g681 ( .A(n_614), .Y(n_681) );
INVx8_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_615), .A2(n_683), .B1(n_749), .B2(n_757), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_615), .A2(n_683), .B1(n_856), .B2(n_862), .Y(n_868) );
OAI22xp33_ASAP7_75t_SL g1043 ( .A1(n_615), .A2(n_1020), .B1(n_1031), .B2(n_1044), .Y(n_1043) );
INVx5_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx3_ASAP7_75t_L g675 ( .A(n_616), .Y(n_675) );
INVx2_ASAP7_75t_SL g763 ( .A(n_616), .Y(n_763) );
INVx2_ASAP7_75t_SL g1391 ( .A(n_616), .Y(n_1391) );
HB1xp67_ASAP7_75t_L g1805 ( .A(n_616), .Y(n_1805) );
OAI33xp33_ASAP7_75t_L g864 ( .A1(n_618), .A2(n_663), .A3(n_865), .B1(n_868), .B2(n_869), .B3(n_870), .Y(n_864) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_622), .B2(n_624), .Y(n_619) );
OAI22xp33_ASAP7_75t_L g793 ( .A1(n_620), .A2(n_794), .B1(n_795), .B2(n_796), .Y(n_793) );
OAI22xp33_ASAP7_75t_L g1094 ( .A1(n_620), .A2(n_1082), .B1(n_1088), .B2(n_1095), .Y(n_1094) );
OAI22xp33_ASAP7_75t_L g1101 ( .A1(n_620), .A2(n_670), .B1(n_1083), .B2(n_1089), .Y(n_1101) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g867 ( .A(n_623), .Y(n_867) );
OAI22xp33_ASAP7_75t_L g1049 ( .A1(n_623), .A2(n_1027), .B1(n_1039), .B2(n_1042), .Y(n_1049) );
OAI22xp33_ASAP7_75t_L g1179 ( .A1(n_623), .A2(n_1042), .B1(n_1180), .B2(n_1181), .Y(n_1179) );
OAI22xp5_ASAP7_75t_L g1232 ( .A1(n_623), .A2(n_1042), .B1(n_1233), .B2(n_1234), .Y(n_1232) );
OAI22xp33_ASAP7_75t_L g1409 ( .A1(n_623), .A2(n_1042), .B1(n_1410), .B2(n_1411), .Y(n_1409) );
OAI22xp33_ASAP7_75t_L g1450 ( .A1(n_623), .A2(n_1451), .B1(n_1452), .B2(n_1453), .Y(n_1450) );
OAI22xp33_ASAP7_75t_L g1493 ( .A1(n_623), .A2(n_1451), .B1(n_1479), .B2(n_1485), .Y(n_1493) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
INVx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_630), .Y(n_641) );
INVx4_ASAP7_75t_L g1026 ( .A(n_630), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_633), .A2(n_696), .B1(n_748), .B2(n_749), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_633), .A2(n_906), .B1(n_908), .B2(n_909), .Y(n_905) );
OAI22xp5_ASAP7_75t_L g1142 ( .A1(n_633), .A2(n_906), .B1(n_1143), .B2(n_1144), .Y(n_1142) );
INVx5_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g702 ( .A(n_641), .Y(n_702) );
INVx3_ASAP7_75t_L g899 ( .A(n_641), .Y(n_899) );
BUFx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI22xp33_ASAP7_75t_L g1024 ( .A1(n_643), .A2(n_1025), .B1(n_1026), .B2(n_1027), .Y(n_1024) );
OAI22xp33_ASAP7_75t_L g1416 ( .A1(n_643), .A2(n_1026), .B1(n_1407), .B2(n_1410), .Y(n_1416) );
OAI33xp33_ASAP7_75t_L g850 ( .A1(n_644), .A2(n_851), .A3(n_852), .B1(n_855), .B2(n_858), .B3(n_861), .Y(n_850) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI22xp33_ASAP7_75t_L g690 ( .A1(n_650), .A2(n_666), .B1(n_691), .B2(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_655), .A2(n_823), .B1(n_824), .B2(n_825), .Y(n_822) );
XNOR2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_769), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_722), .B1(n_767), .B2(n_768), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g768 ( .A(n_659), .Y(n_768) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_703), .C(n_710), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_693), .Y(n_661) );
OAI33xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .A3(n_673), .B1(n_680), .B2(n_687), .B3(n_690), .Y(n_662) );
OAI33xp33_ASAP7_75t_L g758 ( .A1(n_663), .A2(n_759), .A3(n_762), .B1(n_764), .B2(n_765), .B3(n_766), .Y(n_758) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_669), .B2(n_670), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_666), .A2(n_745), .B1(n_753), .B2(n_760), .Y(n_759) );
BUFx4f_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
OAI22xp33_ASAP7_75t_L g775 ( .A1(n_667), .A2(n_776), .B1(n_777), .B2(n_779), .Y(n_775) );
INVx3_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_SL g1451 ( .A(n_668), .Y(n_1451) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_669), .A2(n_692), .B1(n_696), .B2(n_700), .Y(n_699) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g761 ( .A(n_672), .Y(n_761) );
INVx1_ASAP7_75t_L g1114 ( .A(n_672), .Y(n_1114) );
OAI22xp33_ASAP7_75t_SL g673 ( .A1(n_674), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_674), .A2(n_682), .B1(n_696), .B2(n_697), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_675), .A2(n_783), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
OAI22xp5_ASAP7_75t_L g1403 ( .A1(n_675), .A2(n_1231), .B1(n_1404), .B2(n_1405), .Y(n_1403) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_677), .A2(n_748), .B1(n_756), .B2(n_763), .Y(n_762) );
INVx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
BUFx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g1044 ( .A(n_679), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B1(n_683), .B2(n_686), .Y(n_680) );
OAI22xp33_ASAP7_75t_SL g920 ( .A1(n_683), .A2(n_904), .B1(n_913), .B2(n_921), .Y(n_920) );
OAI221xp5_ASAP7_75t_L g1306 ( .A1(n_683), .A2(n_1275), .B1(n_1280), .B2(n_1307), .C(n_1308), .Y(n_1306) );
CKINVDCx8_ASAP7_75t_R g683 ( .A(n_684), .Y(n_683) );
INVx3_ASAP7_75t_L g1227 ( .A(n_684), .Y(n_1227) );
INVx3_ASAP7_75t_L g1231 ( .A(n_684), .Y(n_1231) );
INVx3_ASAP7_75t_L g1322 ( .A(n_684), .Y(n_1322) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g784 ( .A(n_685), .Y(n_784) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
BUFx2_ASAP7_75t_L g1809 ( .A(n_689), .Y(n_1809) );
BUFx2_ASAP7_75t_L g1851 ( .A(n_689), .Y(n_1851) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g806 ( .A(n_698), .Y(n_806) );
INVx2_ASAP7_75t_L g926 ( .A(n_698), .Y(n_926) );
INVx2_ASAP7_75t_L g1188 ( .A(n_698), .Y(n_1188) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_700), .A2(n_751), .B1(n_753), .B2(n_754), .Y(n_750) );
OAI211xp5_ASAP7_75t_SL g1279 ( .A1(n_700), .A2(n_1280), .B(n_1281), .C(n_1286), .Y(n_1279) );
OAI31xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_714), .A3(n_719), .B(n_721), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g957 ( .A(n_717), .Y(n_957) );
OAI31xp33_ASAP7_75t_L g732 ( .A1(n_721), .A2(n_733), .A3(n_734), .B(n_738), .Y(n_732) );
OAI31xp33_ASAP7_75t_L g933 ( .A1(n_721), .A2(n_934), .A3(n_935), .B(n_939), .Y(n_933) );
INVx2_ASAP7_75t_L g767 ( .A(n_722), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_732), .C(n_742), .Y(n_723) );
OAI31xp33_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .A3(n_730), .B(n_731), .Y(n_724) );
OAI31xp33_ASAP7_75t_L g1130 ( .A1(n_731), .A2(n_1131), .A3(n_1135), .B(n_1136), .Y(n_1130) );
OAI21xp5_ASAP7_75t_L g1853 ( .A1(n_731), .A2(n_1854), .B(n_1862), .Y(n_1853) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI22xp33_ASAP7_75t_SL g1298 ( .A1(n_740), .A2(n_824), .B1(n_1267), .B2(n_1299), .Y(n_1298) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_758), .Y(n_742) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_752), .A2(n_1037), .B1(n_1038), .B2(n_1039), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1238 ( .A1(n_752), .A2(n_926), .B1(n_1223), .B2(n_1234), .Y(n_1238) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g1228 ( .A1(n_763), .A2(n_1229), .B1(n_1230), .B2(n_1231), .Y(n_1228) );
OAI22xp5_ASAP7_75t_L g1412 ( .A1(n_763), .A2(n_1044), .B1(n_1413), .B2(n_1414), .Y(n_1412) );
OAI22xp5_ASAP7_75t_L g1492 ( .A1(n_763), .A2(n_1322), .B1(n_1482), .B2(n_1488), .Y(n_1492) );
INVx1_ASAP7_75t_L g982 ( .A(n_765), .Y(n_982) );
OAI33xp33_ASAP7_75t_L g1093 ( .A1(n_765), .A2(n_774), .A3(n_1094), .B1(n_1096), .B2(n_1099), .B3(n_1101), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g1300 ( .A1(n_765), .A2(n_774), .B1(n_1301), .B2(n_1306), .Y(n_1300) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVxp67_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NOR4xp25_ASAP7_75t_L g844 ( .A(n_773), .B(n_798), .C(n_813), .D(n_831), .Y(n_844) );
OAI33xp33_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_775), .A3(n_780), .B1(n_786), .B2(n_791), .B3(n_793), .Y(n_773) );
OAI33xp33_ASAP7_75t_L g1040 ( .A1(n_774), .A2(n_791), .A3(n_1041), .B1(n_1043), .B2(n_1045), .B3(n_1049), .Y(n_1040) );
OAI33xp33_ASAP7_75t_L g1313 ( .A1(n_774), .A2(n_791), .A3(n_1314), .B1(n_1317), .B2(n_1320), .B3(n_1324), .Y(n_1313) );
OAI22xp33_ASAP7_75t_L g1041 ( .A1(n_777), .A2(n_1025), .B1(n_1037), .B2(n_1042), .Y(n_1041) );
OAI22xp5_ASAP7_75t_L g1221 ( .A1(n_777), .A2(n_1042), .B1(n_1222), .B2(n_1223), .Y(n_1221) );
OAI22xp5_ASAP7_75t_SL g1406 ( .A1(n_777), .A2(n_1042), .B1(n_1407), .B2(n_1408), .Y(n_1406) );
OAI22xp5_ASAP7_75t_L g1440 ( .A1(n_777), .A2(n_1042), .B1(n_1441), .B2(n_1442), .Y(n_1440) );
INVx3_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g923 ( .A(n_778), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_782), .B1(n_783), .B2(n_785), .Y(n_780) );
INVx2_ASAP7_75t_L g971 ( .A(n_781), .Y(n_971) );
OAI22xp5_ASAP7_75t_SL g804 ( .A1(n_782), .A2(n_789), .B1(n_805), .B2(n_806), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_783), .A2(n_787), .B1(n_789), .B2(n_790), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g1317 ( .A1(n_783), .A2(n_1307), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
BUFx3_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g1048 ( .A(n_784), .Y(n_1048) );
OR2x2_ASAP7_75t_L g1775 ( .A(n_784), .B(n_1776), .Y(n_1775) );
INVx3_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx3_ASAP7_75t_L g1046 ( .A(n_788), .Y(n_1046) );
INVx2_ASAP7_75t_SL g1174 ( .A(n_788), .Y(n_1174) );
AND2x4_ASAP7_75t_L g1817 ( .A(n_788), .B(n_1818), .Y(n_1817) );
INVx1_ASAP7_75t_L g1394 ( .A(n_791), .Y(n_1394) );
INVx1_ASAP7_75t_L g1125 ( .A(n_795), .Y(n_1125) );
OAI22xp33_ASAP7_75t_L g1158 ( .A1(n_795), .A2(n_917), .B1(n_1141), .B2(n_1147), .Y(n_1158) );
OAI22xp33_ASAP7_75t_L g1169 ( .A1(n_795), .A2(n_1042), .B1(n_1170), .B2(n_1171), .Y(n_1169) );
OAI22xp33_ASAP7_75t_L g1324 ( .A1(n_795), .A2(n_1042), .B1(n_1325), .B2(n_1326), .Y(n_1324) );
OAI22xp33_ASAP7_75t_L g1490 ( .A1(n_795), .A2(n_1451), .B1(n_1478), .B2(n_1484), .Y(n_1490) );
INVxp67_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OAI33xp33_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_802), .A3(n_804), .B1(n_807), .B2(n_808), .B3(n_810), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_SL g1029 ( .A(n_801), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1417 ( .A1(n_805), .A2(n_1038), .B1(n_1404), .B2(n_1413), .Y(n_1417) );
OAI33xp33_ASAP7_75t_L g1018 ( .A1(n_808), .A2(n_1019), .A3(n_1024), .B1(n_1028), .B2(n_1030), .B3(n_1036), .Y(n_1018) );
OAI33xp33_ASAP7_75t_L g1454 ( .A1(n_808), .A2(n_1184), .A3(n_1455), .B1(n_1456), .B2(n_1458), .B3(n_1459), .Y(n_1454) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g1193 ( .A(n_809), .Y(n_1193) );
AOI33xp33_ASAP7_75t_L g1378 ( .A1(n_809), .A2(n_1029), .A3(n_1379), .B1(n_1380), .B2(n_1384), .B3(n_1385), .Y(n_1378) );
NAND3xp33_ASAP7_75t_L g1839 ( .A(n_809), .B(n_1840), .C(n_1842), .Y(n_1839) );
OAI22xp33_ASAP7_75t_L g897 ( .A1(n_811), .A2(n_898), .B1(n_899), .B2(n_900), .Y(n_897) );
OAI22xp5_ASAP7_75t_L g1477 ( .A1(n_811), .A2(n_1026), .B1(n_1478), .B2(n_1479), .Y(n_1477) );
HB1xp67_ASAP7_75t_L g1757 ( .A(n_811), .Y(n_1757) );
INVxp67_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
AOI31xp33_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_822), .A3(n_826), .B(n_829), .Y(n_813) );
INVxp67_ASAP7_75t_SL g815 ( .A(n_816), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g1253 ( .A1(n_818), .A2(n_1208), .B1(n_1245), .B2(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_L g1295 ( .A(n_818), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_818), .B(n_1363), .Y(n_1375) );
AOI22xp33_ASAP7_75t_SL g1423 ( .A1(n_818), .A2(n_1212), .B1(n_1424), .B2(n_1425), .Y(n_1423) );
AOI22xp33_ASAP7_75t_SL g1470 ( .A1(n_818), .A2(n_1212), .B1(n_1463), .B2(n_1471), .Y(n_1470) );
AOI22xp33_ASAP7_75t_SL g1504 ( .A1(n_818), .A2(n_1212), .B1(n_1497), .B2(n_1505), .Y(n_1504) );
INVx2_ASAP7_75t_L g1215 ( .A(n_824), .Y(n_1215) );
AO21x1_ASAP7_75t_L g947 ( .A1(n_829), .A2(n_948), .B(n_951), .Y(n_947) );
CKINVDCx14_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
OAI31xp33_ASAP7_75t_L g1121 ( .A1(n_830), .A2(n_1122), .A3(n_1123), .B(n_1129), .Y(n_1121) );
AOI31xp67_ASAP7_75t_SL g831 ( .A1(n_832), .A2(n_835), .A3(n_840), .B(n_843), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
NAND3xp33_ASAP7_75t_L g1052 ( .A(n_836), .B(n_1053), .C(n_1057), .Y(n_1052) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g1134 ( .A(n_839), .Y(n_1134) );
INVxp67_ASAP7_75t_SL g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g1358 ( .A(n_842), .Y(n_1358) );
INVx1_ASAP7_75t_L g941 ( .A(n_845), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_847), .B1(n_891), .B2(n_892), .Y(n_845) );
INVx2_ASAP7_75t_SL g846 ( .A(n_847), .Y(n_846) );
NAND3xp33_ASAP7_75t_L g848 ( .A(n_849), .B(n_871), .C(n_882), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_850), .B(n_864), .Y(n_849) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_877), .A2(n_902), .B1(n_903), .B2(n_904), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g1145 ( .A1(n_877), .A2(n_906), .B1(n_1146), .B2(n_1147), .Y(n_1145) );
OAI211xp5_ASAP7_75t_L g1747 ( .A1(n_877), .A2(n_1748), .B(n_1749), .C(n_1753), .Y(n_1747) );
OAI31xp33_ASAP7_75t_L g882 ( .A1(n_883), .A2(n_885), .A3(n_889), .B(n_890), .Y(n_882) );
OAI31xp33_ASAP7_75t_L g1109 ( .A1(n_890), .A2(n_1110), .A3(n_1112), .B(n_1117), .Y(n_1109) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
NAND3xp33_ASAP7_75t_L g894 ( .A(n_895), .B(n_924), .C(n_933), .Y(n_894) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_896), .B(n_914), .Y(n_895) );
OAI22xp33_ASAP7_75t_L g922 ( .A1(n_900), .A2(n_909), .B1(n_917), .B2(n_923), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g1330 ( .A1(n_906), .A2(n_1023), .B1(n_1316), .B2(n_1326), .Y(n_1330) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx2_ASAP7_75t_L g1021 ( .A(n_907), .Y(n_1021) );
OAI22xp33_ASAP7_75t_L g1154 ( .A1(n_917), .A2(n_1140), .B1(n_1146), .B2(n_1155), .Y(n_1154) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
OAI22xp33_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_1161), .B1(n_1162), .B2(n_1508), .Y(n_942) );
INVx1_ASAP7_75t_L g1508 ( .A(n_943), .Y(n_1508) );
XNOR2x1_ASAP7_75t_L g943 ( .A(n_944), .B(n_1075), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_1015), .B1(n_1073), .B2(n_1074), .Y(n_944) );
INVx1_ASAP7_75t_L g1074 ( .A(n_945), .Y(n_1074) );
NAND4xp25_ASAP7_75t_SL g946 ( .A(n_947), .B(n_959), .C(n_983), .D(n_1006), .Y(n_946) );
INVx2_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
AOI33xp33_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_963), .A3(n_970), .B1(n_976), .B2(n_979), .B3(n_982), .Y(n_959) );
BUFx3_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g1398 ( .A(n_961), .Y(n_1398) );
AOI33xp33_ASAP7_75t_L g1802 ( .A1(n_961), .A2(n_1803), .A3(n_1804), .B1(n_1807), .B2(n_1809), .B3(n_1810), .Y(n_1802) );
NAND3xp33_ASAP7_75t_L g1843 ( .A(n_961), .B(n_1844), .C(n_1846), .Y(n_1843) );
INVx1_ASAP7_75t_L g1771 ( .A(n_962), .Y(n_1771) );
BUFx2_ASAP7_75t_SL g964 ( .A(n_965), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx2_ASAP7_75t_SL g966 ( .A(n_967), .Y(n_966) );
INVx2_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g1811 ( .A(n_969), .Y(n_1811) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx2_ASAP7_75t_L g981 ( .A(n_973), .Y(n_981) );
INVx2_ASAP7_75t_R g1806 ( .A(n_973), .Y(n_1806) );
INVx5_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
BUFx2_ASAP7_75t_L g1305 ( .A(n_974), .Y(n_1305) );
BUFx12f_ASAP7_75t_L g1392 ( .A(n_974), .Y(n_1392) );
BUFx3_ASAP7_75t_L g1808 ( .A(n_974), .Y(n_1808) );
BUFx3_ASAP7_75t_L g1845 ( .A(n_974), .Y(n_1845) );
INVx1_ASAP7_75t_L g1209 ( .A(n_975), .Y(n_1209) );
BUFx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
AND2x4_ASAP7_75t_L g1821 ( .A(n_978), .B(n_1797), .Y(n_1821) );
INVx1_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
INVx2_ASAP7_75t_SL g1003 ( .A(n_987), .Y(n_1003) );
INVx2_ASAP7_75t_L g1287 ( .A(n_987), .Y(n_1287) );
INVx1_ASAP7_75t_L g1386 ( .A(n_987), .Y(n_1386) );
INVx3_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
BUFx6f_ASAP7_75t_L g1347 ( .A(n_988), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_988), .B(n_1732), .Y(n_1739) );
NAND2xp5_ASAP7_75t_L g1780 ( .A(n_988), .B(n_1735), .Y(n_1780) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
BUFx3_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
INVx2_ASAP7_75t_L g1005 ( .A(n_992), .Y(n_1005) );
BUFx6f_ASAP7_75t_L g1387 ( .A(n_992), .Y(n_1387) );
INVx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx2_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g1761 ( .A(n_996), .Y(n_1761) );
INVx2_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1367 ( .A(n_999), .Y(n_1367) );
INVx2_ASAP7_75t_L g1383 ( .A(n_999), .Y(n_1383) );
BUFx2_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1000), .Y(n_1198) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
AO21x1_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1008), .B(n_1014), .Y(n_1006) );
INVx2_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
NAND2xp5_ASAP7_75t_SL g1270 ( .A(n_1011), .B(n_1271), .Y(n_1270) );
AO21x1_ASAP7_75t_L g1355 ( .A1(n_1014), .A2(n_1356), .B(n_1360), .Y(n_1355) );
INVx3_ASAP7_75t_SL g1073 ( .A(n_1015), .Y(n_1073) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1016), .Y(n_1072) );
NAND3xp33_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1050), .C(n_1063), .Y(n_1016) );
NOR2xp33_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1040), .Y(n_1017) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_1020), .A2(n_1021), .B1(n_1022), .B2(n_1023), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_1021), .A2(n_1173), .B1(n_1177), .B2(n_1188), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_1021), .A2(n_1171), .B1(n_1181), .B2(n_1188), .Y(n_1189) );
OAI22xp5_ASAP7_75t_L g1237 ( .A1(n_1021), .A2(n_1038), .B1(n_1225), .B2(n_1229), .Y(n_1237) );
OAI22xp5_ASAP7_75t_L g1418 ( .A1(n_1021), .A2(n_1188), .B1(n_1408), .B2(n_1411), .Y(n_1418) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_1022), .A2(n_1035), .B1(n_1046), .B2(n_1047), .Y(n_1045) );
OAI22xp5_ASAP7_75t_L g1483 ( .A1(n_1023), .A2(n_1457), .B1(n_1484), .B2(n_1485), .Y(n_1483) );
OAI22xp5_ASAP7_75t_L g1185 ( .A1(n_1026), .A2(n_1170), .B1(n_1180), .B2(n_1186), .Y(n_1185) );
OAI22xp5_ASAP7_75t_L g1419 ( .A1(n_1026), .A2(n_1186), .B1(n_1405), .B2(n_1414), .Y(n_1419) );
OAI22xp5_ASAP7_75t_L g1455 ( .A1(n_1026), .A2(n_1033), .B1(n_1441), .B2(n_1452), .Y(n_1455) );
OAI22xp5_ASAP7_75t_L g1459 ( .A1(n_1026), .A2(n_1186), .B1(n_1445), .B2(n_1449), .Y(n_1459) );
OAI22xp5_ASAP7_75t_L g1486 ( .A1(n_1026), .A2(n_1033), .B1(n_1487), .B2(n_1488), .Y(n_1486) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
NAND3xp33_ASAP7_75t_L g1832 ( .A(n_1029), .B(n_1833), .C(n_1837), .Y(n_1832) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_1031), .A2(n_1032), .B1(n_1033), .B2(n_1035), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_1032), .A2(n_1033), .B1(n_1222), .B2(n_1233), .Y(n_1236) );
OAI22xp5_ASAP7_75t_L g1239 ( .A1(n_1032), .A2(n_1186), .B1(n_1226), .B2(n_1230), .Y(n_1239) );
OAI22xp5_ASAP7_75t_L g1328 ( .A1(n_1032), .A2(n_1186), .B1(n_1315), .B2(n_1325), .Y(n_1328) );
OAI22xp5_ASAP7_75t_L g1331 ( .A1(n_1033), .A2(n_1319), .B1(n_1323), .B2(n_1332), .Y(n_1331) );
BUFx6f_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
OAI22xp33_ASAP7_75t_L g1314 ( .A1(n_1042), .A2(n_1294), .B1(n_1315), .B2(n_1316), .Y(n_1314) );
OAI22xp5_ASAP7_75t_L g1172 ( .A1(n_1044), .A2(n_1173), .B1(n_1174), .B2(n_1175), .Y(n_1172) );
OAI22xp5_ASAP7_75t_L g1446 ( .A1(n_1044), .A2(n_1447), .B1(n_1448), .B2(n_1449), .Y(n_1446) );
OAI22xp5_ASAP7_75t_L g1320 ( .A1(n_1046), .A2(n_1321), .B1(n_1322), .B2(n_1323), .Y(n_1320) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
AOI22xp5_ASAP7_75t_L g1496 ( .A1(n_1055), .A2(n_1265), .B1(n_1497), .B2(n_1498), .Y(n_1496) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1059), .Y(n_1057) );
OAI31xp33_ASAP7_75t_L g1063 ( .A1(n_1064), .A2(n_1066), .A3(n_1069), .B(n_1070), .Y(n_1063) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1070), .Y(n_1377) );
OA22x2_ASAP7_75t_L g1075 ( .A1(n_1076), .A2(n_1077), .B1(n_1118), .B2(n_1119), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
NAND3xp33_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1102), .C(n_1109), .Y(n_1078) );
NOR2xp33_ASAP7_75t_SL g1079 ( .A(n_1080), .B(n_1093), .Y(n_1079) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVxp67_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1114), .Y(n_1155) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1120), .Y(n_1159) );
NAND3xp33_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1130), .C(n_1137), .Y(n_1120) );
INVx2_ASAP7_75t_SL g1124 ( .A(n_1125), .Y(n_1124) );
NOR2xp33_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1153), .Y(n_1137) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
XOR2x2_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1351), .Y(n_1162) );
XNOR2xp5_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1255), .Y(n_1163) );
XNOR2xp5_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1217), .Y(n_1164) );
NAND3xp33_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1194), .C(n_1204), .Y(n_1166) );
NOR2xp33_ASAP7_75t_SL g1167 ( .A(n_1168), .B(n_1183), .Y(n_1167) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_1175), .A2(n_1178), .B1(n_1186), .B2(n_1191), .Y(n_1190) );
OAI33xp33_ASAP7_75t_L g1183 ( .A1(n_1184), .A2(n_1185), .A3(n_1187), .B1(n_1189), .B2(n_1190), .B3(n_1193), .Y(n_1183) );
OAI33xp33_ASAP7_75t_L g1327 ( .A1(n_1184), .A2(n_1193), .A3(n_1328), .B1(n_1329), .B2(n_1330), .B3(n_1331), .Y(n_1327) );
OAI33xp33_ASAP7_75t_L g1415 ( .A1(n_1184), .A2(n_1193), .A3(n_1416), .B1(n_1417), .B2(n_1418), .B3(n_1419), .Y(n_1415) );
OAI22xp5_ASAP7_75t_L g1456 ( .A1(n_1188), .A2(n_1444), .B1(n_1447), .B2(n_1457), .Y(n_1456) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
NAND3xp33_ASAP7_75t_SL g1341 ( .A(n_1196), .B(n_1342), .C(n_1344), .Y(n_1341) );
NAND3xp33_ASAP7_75t_L g1854 ( .A(n_1196), .B(n_1855), .C(n_1858), .Y(n_1854) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
INVx2_ASAP7_75t_L g1365 ( .A(n_1197), .Y(n_1365) );
AOI32xp33_ASAP7_75t_L g1207 ( .A1(n_1201), .A2(n_1208), .A3(n_1210), .B1(n_1212), .B2(n_1213), .Y(n_1207) );
OAI31xp33_ASAP7_75t_SL g1204 ( .A1(n_1205), .A2(n_1206), .A3(n_1214), .B(n_1216), .Y(n_1204) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1209), .Y(n_1801) );
AND2x2_ASAP7_75t_L g1796 ( .A(n_1210), .B(n_1797), .Y(n_1796) );
INVx3_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVxp67_ASAP7_75t_L g1252 ( .A(n_1212), .Y(n_1252) );
INVxp67_ASAP7_75t_L g1296 ( .A(n_1212), .Y(n_1296) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1212), .Y(n_1374) );
OAI31xp33_ASAP7_75t_SL g1248 ( .A1(n_1216), .A2(n_1249), .A3(n_1250), .B(n_1251), .Y(n_1248) );
OAI21xp5_ASAP7_75t_L g1333 ( .A1(n_1216), .A2(n_1334), .B(n_1339), .Y(n_1333) );
OAI31xp33_ASAP7_75t_L g1420 ( .A1(n_1216), .A2(n_1421), .A3(n_1422), .B(n_1426), .Y(n_1420) );
OAI31xp33_ASAP7_75t_SL g1467 ( .A1(n_1216), .A2(n_1468), .A3(n_1469), .B(n_1472), .Y(n_1467) );
OAI31xp33_ASAP7_75t_SL g1501 ( .A1(n_1216), .A2(n_1502), .A3(n_1503), .B(n_1506), .Y(n_1501) );
OAI21xp5_ASAP7_75t_L g1863 ( .A1(n_1216), .A2(n_1864), .B(n_1865), .Y(n_1863) );
NAND3xp33_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1240), .C(n_1248), .Y(n_1218) );
NOR2xp33_ASAP7_75t_SL g1219 ( .A(n_1220), .B(n_1235), .Y(n_1219) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1242), .Y(n_1349) );
XOR2xp5_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1310), .Y(n_1255) );
OAI21xp5_ASAP7_75t_L g1257 ( .A1(n_1258), .A2(n_1288), .B(n_1290), .Y(n_1257) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
OAI21xp5_ASAP7_75t_L g1272 ( .A1(n_1273), .A2(n_1276), .B(n_1279), .Y(n_1272) );
BUFx6f_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx2_ASAP7_75t_L g1382 ( .A(n_1283), .Y(n_1382) );
AND2x4_ASAP7_75t_L g1731 ( .A(n_1283), .B(n_1732), .Y(n_1731) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
INVx3_ASAP7_75t_L g1754 ( .A(n_1285), .Y(n_1754) );
BUFx2_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
NAND2xp5_ASAP7_75t_SL g1291 ( .A(n_1292), .B(n_1298), .Y(n_1291) );
NAND3xp33_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1333), .C(n_1340), .Y(n_1311) );
NOR2xp33_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1327), .Y(n_1312) );
OAI221xp5_ASAP7_75t_L g1755 ( .A1(n_1332), .A2(n_1756), .B1(n_1757), .B2(n_1758), .C(n_1759), .Y(n_1755) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_1345), .A2(n_1346), .B1(n_1348), .B2(n_1349), .Y(n_1344) );
INVx3_ASAP7_75t_L g1751 ( .A(n_1347), .Y(n_1751) );
BUFx6f_ASAP7_75t_L g1841 ( .A(n_1347), .Y(n_1841) );
AOI22xp5_ASAP7_75t_L g1351 ( .A1(n_1352), .A2(n_1433), .B1(n_1434), .B2(n_1507), .Y(n_1351) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1352), .Y(n_1507) );
XNOR2x1_ASAP7_75t_SL g1352 ( .A(n_1353), .B(n_1399), .Y(n_1352) );
NAND4xp75_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1370), .C(n_1378), .D(n_1388), .Y(n_1354) );
NOR2xp33_ASAP7_75t_L g1360 ( .A(n_1361), .B(n_1369), .Y(n_1360) );
NAND3xp33_ASAP7_75t_L g1361 ( .A(n_1362), .B(n_1365), .C(n_1366), .Y(n_1361) );
NAND2xp5_ASAP7_75t_L g1366 ( .A(n_1367), .B(n_1368), .Y(n_1366) );
AO21x1_ASAP7_75t_L g1370 ( .A1(n_1371), .A2(n_1372), .B(n_1377), .Y(n_1370) );
INVx2_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
AND2x4_ASAP7_75t_L g1741 ( .A(n_1387), .B(n_1732), .Y(n_1741) );
BUFx2_ASAP7_75t_L g1752 ( .A(n_1387), .Y(n_1752) );
AOI32xp33_ASAP7_75t_L g1388 ( .A1(n_1389), .A2(n_1393), .A3(n_1394), .B1(n_1395), .B2(n_1396), .Y(n_1388) );
INVx2_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
AND3x1_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1420), .C(n_1427), .Y(n_1400) );
NOR2xp33_ASAP7_75t_L g1401 ( .A(n_1402), .B(n_1415), .Y(n_1401) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
XNOR2x1_ASAP7_75t_L g1434 ( .A(n_1435), .B(n_1473), .Y(n_1434) );
XNOR2xp5_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1437), .Y(n_1435) );
AND3x1_ASAP7_75t_L g1437 ( .A(n_1438), .B(n_1460), .C(n_1467), .Y(n_1437) );
NOR2xp33_ASAP7_75t_SL g1438 ( .A(n_1439), .B(n_1454), .Y(n_1438) );
OR2x2_ASAP7_75t_L g1813 ( .A(n_1451), .B(n_1814), .Y(n_1813) );
AND3x1_ASAP7_75t_L g1474 ( .A(n_1475), .B(n_1494), .C(n_1501), .Y(n_1474) );
NOR2xp33_ASAP7_75t_L g1475 ( .A(n_1476), .B(n_1489), .Y(n_1475) );
OAI221xp5_ASAP7_75t_L g1509 ( .A1(n_1510), .A2(n_1723), .B1(n_1725), .B2(n_1822), .C(n_1826), .Y(n_1509) );
AOI21xp5_ASAP7_75t_L g1510 ( .A1(n_1511), .A2(n_1634), .B(n_1693), .Y(n_1510) );
NAND5xp2_ASAP7_75t_L g1511 ( .A(n_1512), .B(n_1577), .C(n_1597), .D(n_1610), .E(n_1620), .Y(n_1511) );
O2A1O1Ixp33_ASAP7_75t_L g1512 ( .A1(n_1513), .A2(n_1544), .B(n_1551), .C(n_1562), .Y(n_1512) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1513), .Y(n_1581) );
AND2x2_ASAP7_75t_L g1513 ( .A(n_1514), .B(n_1534), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1570 ( .A(n_1514), .B(n_1541), .Y(n_1570) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1514), .B(n_1536), .Y(n_1609) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1514), .B(n_1535), .Y(n_1638) );
NAND2xp5_ASAP7_75t_L g1646 ( .A(n_1514), .B(n_1647), .Y(n_1646) );
NAND2xp5_ASAP7_75t_L g1682 ( .A(n_1514), .B(n_1548), .Y(n_1682) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1514), .Y(n_1705) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1515), .B(n_1530), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_1515), .B(n_1576), .Y(n_1575) );
NAND2xp5_ASAP7_75t_L g1588 ( .A(n_1515), .B(n_1535), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1515), .B(n_1531), .Y(n_1596) );
AND3x1_ASAP7_75t_L g1670 ( .A(n_1515), .B(n_1531), .C(n_1535), .Y(n_1670) );
OR2x2_ASAP7_75t_L g1711 ( .A(n_1515), .B(n_1576), .Y(n_1711) );
INVx2_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_1516), .B(n_1530), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1516), .B(n_1531), .Y(n_1601) );
OR2x2_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1524), .Y(n_1516) );
INVx2_ASAP7_75t_L g1631 ( .A(n_1518), .Y(n_1631) );
AND2x6_ASAP7_75t_L g1518 ( .A(n_1519), .B(n_1520), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1522 ( .A(n_1519), .B(n_1523), .Y(n_1522) );
AND2x4_ASAP7_75t_L g1525 ( .A(n_1519), .B(n_1526), .Y(n_1525) );
AND2x6_ASAP7_75t_L g1528 ( .A(n_1519), .B(n_1529), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1519), .B(n_1523), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1560 ( .A(n_1519), .B(n_1523), .Y(n_1560) );
OAI21xp5_ASAP7_75t_L g1870 ( .A1(n_1520), .A2(n_1871), .B(n_1872), .Y(n_1870) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1521), .B(n_1527), .Y(n_1526) );
INVxp67_ASAP7_75t_L g1633 ( .A(n_1522), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_1530), .B(n_1576), .Y(n_1673) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
OR2x2_ASAP7_75t_L g1606 ( .A(n_1531), .B(n_1576), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1667 ( .A(n_1531), .B(n_1576), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_1532), .B(n_1533), .Y(n_1531) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1534), .B(n_1596), .Y(n_1595) );
NAND2xp5_ASAP7_75t_L g1681 ( .A(n_1534), .B(n_1601), .Y(n_1681) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1534), .Y(n_1708) );
AND2x2_ASAP7_75t_L g1534 ( .A(n_1535), .B(n_1540), .Y(n_1534) );
AND2x2_ASAP7_75t_L g1616 ( .A(n_1535), .B(n_1550), .Y(n_1616) );
OR2x2_ASAP7_75t_L g1618 ( .A(n_1535), .B(n_1619), .Y(n_1618) );
INVx2_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1536), .B(n_1550), .Y(n_1549) );
OAI322xp33_ASAP7_75t_L g1562 ( .A1(n_1536), .A2(n_1558), .A3(n_1563), .B1(n_1569), .B2(n_1571), .C1(n_1573), .C2(n_1574), .Y(n_1562) );
BUFx2_ASAP7_75t_L g1576 ( .A(n_1536), .Y(n_1576) );
OR2x2_ASAP7_75t_L g1599 ( .A(n_1536), .B(n_1600), .Y(n_1599) );
AOI321xp33_ASAP7_75t_L g1620 ( .A1(n_1536), .A2(n_1621), .A3(n_1622), .B1(n_1623), .B2(n_1625), .C(n_1627), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1658 ( .A(n_1536), .B(n_1601), .Y(n_1658) );
OR2x2_ASAP7_75t_L g1719 ( .A(n_1536), .B(n_1653), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1536 ( .A(n_1537), .B(n_1538), .Y(n_1536) );
NAND2xp5_ASAP7_75t_L g1615 ( .A(n_1540), .B(n_1552), .Y(n_1615) );
NAND2xp5_ASAP7_75t_L g1619 ( .A(n_1540), .B(n_1601), .Y(n_1619) );
NOR2xp33_ASAP7_75t_L g1625 ( .A(n_1540), .B(n_1626), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1668 ( .A(n_1540), .B(n_1592), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g1692 ( .A(n_1540), .B(n_1550), .Y(n_1692) );
OAI21xp33_ASAP7_75t_L g1713 ( .A1(n_1540), .A2(n_1692), .B(n_1714), .Y(n_1713) );
INVx2_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1541), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_1541), .B(n_1554), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1541), .B(n_1558), .Y(n_1622) );
AND2x2_ASAP7_75t_L g1645 ( .A(n_1541), .B(n_1576), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1653 ( .A(n_1541), .B(n_1601), .Y(n_1653) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_1541), .B(n_1566), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1541 ( .A(n_1542), .B(n_1543), .Y(n_1541) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
NAND2xp5_ASAP7_75t_L g1545 ( .A(n_1546), .B(n_1549), .Y(n_1545) );
NAND2xp5_ASAP7_75t_L g1675 ( .A(n_1546), .B(n_1611), .Y(n_1675) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
NAND2xp5_ASAP7_75t_L g1563 ( .A(n_1547), .B(n_1564), .Y(n_1563) );
NOR2xp33_ASAP7_75t_L g1605 ( .A(n_1547), .B(n_1606), .Y(n_1605) );
NAND2xp5_ASAP7_75t_L g1637 ( .A(n_1547), .B(n_1638), .Y(n_1637) );
AND2x2_ASAP7_75t_L g1669 ( .A(n_1547), .B(n_1670), .Y(n_1669) );
AND2x2_ASAP7_75t_L g1677 ( .A(n_1547), .B(n_1616), .Y(n_1677) );
INVx2_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1647 ( .A(n_1548), .B(n_1564), .Y(n_1647) );
O2A1O1Ixp33_ASAP7_75t_L g1721 ( .A1(n_1548), .A2(n_1690), .B(n_1691), .C(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1549), .Y(n_1722) );
OR2x2_ASAP7_75t_L g1621 ( .A(n_1550), .B(n_1596), .Y(n_1621) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1550), .Y(n_1691) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1557), .Y(n_1551) );
NAND2xp5_ASAP7_75t_L g1624 ( .A(n_1552), .B(n_1558), .Y(n_1624) );
INVx2_ASAP7_75t_L g1642 ( .A(n_1552), .Y(n_1642) );
A2O1A1O1Ixp25_ASAP7_75t_L g1687 ( .A1(n_1552), .A2(n_1566), .B(n_1644), .C(n_1688), .D(n_1689), .Y(n_1687) );
OR2x2_ASAP7_75t_L g1702 ( .A(n_1552), .B(n_1703), .Y(n_1702) );
INVx2_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1572 ( .A(n_1553), .B(n_1557), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1553), .B(n_1566), .Y(n_1580) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
OR2x2_ASAP7_75t_L g1565 ( .A(n_1554), .B(n_1566), .Y(n_1565) );
AND2x2_ASAP7_75t_L g1592 ( .A(n_1554), .B(n_1593), .Y(n_1592) );
AND2x2_ASAP7_75t_L g1680 ( .A(n_1554), .B(n_1566), .Y(n_1680) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_1555), .B(n_1556), .Y(n_1554) );
NAND2xp5_ASAP7_75t_L g1573 ( .A(n_1557), .B(n_1564), .Y(n_1573) );
NOR2xp33_ASAP7_75t_L g1604 ( .A(n_1557), .B(n_1565), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1557), .B(n_1592), .Y(n_1639) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1557), .B(n_1566), .Y(n_1649) );
OR2x2_ASAP7_75t_L g1660 ( .A(n_1557), .B(n_1566), .Y(n_1660) );
CKINVDCx6p67_ASAP7_75t_R g1557 ( .A(n_1558), .Y(n_1557) );
OR2x2_ASAP7_75t_L g1603 ( .A(n_1558), .B(n_1566), .Y(n_1603) );
AND2x2_ASAP7_75t_L g1611 ( .A(n_1558), .B(n_1566), .Y(n_1611) );
NAND2xp5_ASAP7_75t_L g1684 ( .A(n_1558), .B(n_1685), .Y(n_1684) );
CKINVDCx5p33_ASAP7_75t_R g1706 ( .A(n_1558), .Y(n_1706) );
OR2x2_ASAP7_75t_L g1709 ( .A(n_1558), .B(n_1579), .Y(n_1709) );
OR2x6_ASAP7_75t_L g1558 ( .A(n_1559), .B(n_1561), .Y(n_1558) );
OR2x2_ASAP7_75t_L g1662 ( .A(n_1559), .B(n_1561), .Y(n_1662) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1563), .Y(n_1695) );
NAND2xp5_ASAP7_75t_L g1589 ( .A(n_1564), .B(n_1570), .Y(n_1589) );
INVx2_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
INVx3_ASAP7_75t_L g1584 ( .A(n_1566), .Y(n_1584) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1566), .Y(n_1593) );
AOI22xp5_ASAP7_75t_L g1610 ( .A1(n_1566), .A2(n_1611), .B1(n_1612), .B2(n_1617), .Y(n_1610) );
AND2x4_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1568), .Y(n_1566) );
INVxp67_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
NAND2xp5_ASAP7_75t_L g1608 ( .A(n_1572), .B(n_1609), .Y(n_1608) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1573), .Y(n_1720) );
CKINVDCx14_ASAP7_75t_R g1574 ( .A(n_1575), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1576), .B(n_1596), .Y(n_1650) );
NOR2xp33_ASAP7_75t_L g1577 ( .A(n_1578), .B(n_1590), .Y(n_1577) );
OAI211xp5_ASAP7_75t_L g1578 ( .A1(n_1579), .A2(n_1581), .B(n_1582), .C(n_1589), .Y(n_1578) );
AOI21xp33_ASAP7_75t_L g1651 ( .A1(n_1579), .A2(n_1652), .B(n_1653), .Y(n_1651) );
CKINVDCx6p67_ASAP7_75t_R g1579 ( .A(n_1580), .Y(n_1579) );
AOI21xp33_ASAP7_75t_L g1715 ( .A1(n_1581), .A2(n_1656), .B(n_1716), .Y(n_1715) );
NAND2xp5_ASAP7_75t_L g1582 ( .A(n_1583), .B(n_1585), .Y(n_1582) );
CKINVDCx14_ASAP7_75t_R g1583 ( .A(n_1584), .Y(n_1583) );
AOI221xp5_ASAP7_75t_L g1717 ( .A1(n_1585), .A2(n_1611), .B1(n_1718), .B2(n_1720), .C(n_1721), .Y(n_1717) );
NOR2xp33_ASAP7_75t_L g1585 ( .A(n_1586), .B(n_1588), .Y(n_1585) );
CKINVDCx14_ASAP7_75t_R g1586 ( .A(n_1587), .Y(n_1586) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1588), .Y(n_1685) );
NOR2xp33_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1594), .Y(n_1590) );
AOI21xp5_ASAP7_75t_L g1696 ( .A1(n_1591), .A2(n_1697), .B(n_1698), .Y(n_1696) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1596), .Y(n_1626) );
AOI221xp5_ASAP7_75t_L g1597 ( .A1(n_1598), .A2(n_1602), .B1(n_1604), .B2(n_1605), .C(n_1607), .Y(n_1597) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
NAND2xp5_ASAP7_75t_L g1671 ( .A(n_1599), .B(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1644 ( .A(n_1601), .B(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
NAND2xp5_ASAP7_75t_L g1652 ( .A(n_1603), .B(n_1609), .Y(n_1652) );
OAI221xp5_ASAP7_75t_L g1689 ( .A1(n_1603), .A2(n_1627), .B1(n_1690), .B2(n_1691), .C(n_1692), .Y(n_1689) );
AOI221xp5_ASAP7_75t_L g1699 ( .A1(n_1604), .A2(n_1638), .B1(n_1700), .B2(n_1706), .C(n_1707), .Y(n_1699) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
AOI222xp33_ASAP7_75t_L g1663 ( .A1(n_1611), .A2(n_1664), .B1(n_1668), .B2(n_1669), .C1(n_1671), .C2(n_1674), .Y(n_1663) );
NAND2xp5_ASAP7_75t_L g1690 ( .A(n_1611), .B(n_1642), .Y(n_1690) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
NOR2xp33_ASAP7_75t_L g1661 ( .A(n_1613), .B(n_1662), .Y(n_1661) );
NAND2xp5_ASAP7_75t_L g1613 ( .A(n_1614), .B(n_1616), .Y(n_1613) );
OAI21xp33_ASAP7_75t_L g1648 ( .A1(n_1614), .A2(n_1649), .B(n_1650), .Y(n_1648) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1616), .Y(n_1665) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
AOI211xp5_ASAP7_75t_SL g1707 ( .A1(n_1619), .A2(n_1708), .B(n_1709), .C(n_1710), .Y(n_1707) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
OAI22xp5_ASAP7_75t_L g1678 ( .A1(n_1624), .A2(n_1679), .B1(n_1681), .B2(n_1682), .Y(n_1678) );
INVx2_ASAP7_75t_SL g1627 ( .A(n_1628), .Y(n_1627) );
OAI22xp5_ASAP7_75t_SL g1629 ( .A1(n_1630), .A2(n_1631), .B1(n_1632), .B2(n_1633), .Y(n_1629) );
CKINVDCx20_ASAP7_75t_R g1724 ( .A(n_1631), .Y(n_1724) );
NAND5xp2_ASAP7_75t_L g1634 ( .A(n_1635), .B(n_1654), .C(n_1663), .D(n_1676), .E(n_1687), .Y(n_1634) );
AOI211xp5_ASAP7_75t_L g1635 ( .A1(n_1636), .A2(n_1639), .B(n_1640), .C(n_1651), .Y(n_1635) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
AOI221xp5_ASAP7_75t_L g1712 ( .A1(n_1639), .A2(n_1669), .B1(n_1680), .B2(n_1713), .C(n_1715), .Y(n_1712) );
OAI211xp5_ASAP7_75t_L g1640 ( .A1(n_1641), .A2(n_1643), .B(n_1646), .C(n_1648), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1656 ( .A(n_1641), .B(n_1657), .Y(n_1656) );
INVx2_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1645), .Y(n_1704) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1647), .Y(n_1686) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1649), .Y(n_1716) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1650), .Y(n_1714) );
INVxp67_ASAP7_75t_SL g1688 ( .A(n_1652), .Y(n_1688) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1653), .Y(n_1657) );
O2A1O1Ixp33_ASAP7_75t_SL g1654 ( .A1(n_1655), .A2(n_1658), .B(n_1659), .C(n_1661), .Y(n_1654) );
INVxp67_ASAP7_75t_SL g1655 ( .A(n_1656), .Y(n_1655) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1658), .Y(n_1698) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
AOI211xp5_ASAP7_75t_L g1676 ( .A1(n_1662), .A2(n_1677), .B(n_1678), .C(n_1683), .Y(n_1676) );
A2O1A1Ixp33_ASAP7_75t_L g1694 ( .A1(n_1662), .A2(n_1667), .B(n_1695), .C(n_1696), .Y(n_1694) );
NAND2xp5_ASAP7_75t_SL g1664 ( .A(n_1665), .B(n_1666), .Y(n_1664) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
AOI21xp33_ASAP7_75t_L g1683 ( .A1(n_1672), .A2(n_1684), .B(n_1686), .Y(n_1683) );
OAI21xp33_ASAP7_75t_L g1700 ( .A1(n_1672), .A2(n_1701), .B(n_1702), .Y(n_1700) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1673), .Y(n_1672) );
INVxp67_ASAP7_75t_SL g1674 ( .A(n_1675), .Y(n_1674) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1677), .Y(n_1697) );
INVx2_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
NAND4xp25_ASAP7_75t_L g1693 ( .A(n_1694), .B(n_1699), .C(n_1712), .D(n_1717), .Y(n_1693) );
OR2x2_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1705), .Y(n_1703) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
CKINVDCx20_ASAP7_75t_R g1723 ( .A(n_1724), .Y(n_1723) );
NAND3xp33_ASAP7_75t_L g1726 ( .A(n_1727), .B(n_1772), .C(n_1792), .Y(n_1726) );
OAI31xp33_ASAP7_75t_L g1727 ( .A1(n_1728), .A2(n_1742), .A3(n_1763), .B(n_1768), .Y(n_1727) );
NAND2xp5_ASAP7_75t_L g1728 ( .A(n_1729), .B(n_1736), .Y(n_1728) );
AOI21xp5_ASAP7_75t_L g1729 ( .A1(n_1730), .A2(n_1733), .B(n_1734), .Y(n_1729) );
BUFx6f_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1735), .Y(n_1746) );
AOI22xp33_ASAP7_75t_L g1736 ( .A1(n_1737), .A2(n_1738), .B1(n_1740), .B2(n_1741), .Y(n_1736) );
BUFx6f_ASAP7_75t_L g1738 ( .A(n_1739), .Y(n_1738) );
INVx2_ASAP7_75t_L g1743 ( .A(n_1744), .Y(n_1743) );
NOR2x1_ASAP7_75t_L g1744 ( .A(n_1745), .B(n_1746), .Y(n_1744) );
INVx2_ASAP7_75t_SL g1750 ( .A(n_1751), .Y(n_1750) );
INVx2_ASAP7_75t_L g1838 ( .A(n_1751), .Y(n_1838) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
INVx2_ASAP7_75t_L g1764 ( .A(n_1765), .Y(n_1764) );
INVx4_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
INVx2_ASAP7_75t_L g1766 ( .A(n_1767), .Y(n_1766) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
INVx1_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
BUFx2_ASAP7_75t_L g1770 ( .A(n_1771), .Y(n_1770) );
AOI21xp33_ASAP7_75t_SL g1772 ( .A1(n_1773), .A2(n_1781), .B(n_1782), .Y(n_1772) );
INVx8_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
AND2x4_ASAP7_75t_L g1774 ( .A(n_1775), .B(n_1778), .Y(n_1774) );
INVx1_ASAP7_75t_L g1815 ( .A(n_1776), .Y(n_1815) );
INVx1_ASAP7_75t_L g1818 ( .A(n_1776), .Y(n_1818) );
OR2x2_ASAP7_75t_L g1778 ( .A(n_1779), .B(n_1780), .Y(n_1778) );
AND2x4_ASAP7_75t_L g1797 ( .A(n_1779), .B(n_1789), .Y(n_1797) );
AND2x4_ASAP7_75t_L g1783 ( .A(n_1784), .B(n_1786), .Y(n_1783) );
OR2x2_ASAP7_75t_L g1787 ( .A(n_1788), .B(n_1791), .Y(n_1787) );
NOR3xp33_ASAP7_75t_L g1792 ( .A(n_1793), .B(n_1812), .C(n_1819), .Y(n_1792) );
NAND2xp5_ASAP7_75t_L g1793 ( .A(n_1794), .B(n_1802), .Y(n_1793) );
AOI22xp33_ASAP7_75t_L g1794 ( .A1(n_1795), .A2(n_1796), .B1(n_1798), .B2(n_1799), .Y(n_1794) );
AND2x4_ASAP7_75t_L g1799 ( .A(n_1797), .B(n_1800), .Y(n_1799) );
INVx2_ASAP7_75t_L g1800 ( .A(n_1801), .Y(n_1800) );
INVxp67_ASAP7_75t_L g1814 ( .A(n_1815), .Y(n_1814) );
INVx2_ASAP7_75t_L g1816 ( .A(n_1817), .Y(n_1816) );
INVx1_ASAP7_75t_L g1819 ( .A(n_1820), .Y(n_1819) );
INVx3_ASAP7_75t_L g1820 ( .A(n_1821), .Y(n_1820) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1823), .Y(n_1822) );
BUFx3_ASAP7_75t_L g1823 ( .A(n_1824), .Y(n_1823) );
INVxp33_ASAP7_75t_SL g1827 ( .A(n_1828), .Y(n_1827) );
HB1xp67_ASAP7_75t_L g1829 ( .A(n_1830), .Y(n_1829) );
NAND3xp33_ASAP7_75t_L g1830 ( .A(n_1831), .B(n_1853), .C(n_1863), .Y(n_1830) );
AND4x1_ASAP7_75t_L g1831 ( .A(n_1832), .B(n_1839), .C(n_1843), .D(n_1849), .Y(n_1831) );
INVx1_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
INVx1_ASAP7_75t_L g1835 ( .A(n_1836), .Y(n_1835) );
INVx1_ASAP7_75t_L g1847 ( .A(n_1848), .Y(n_1847) );
NAND3xp33_ASAP7_75t_L g1849 ( .A(n_1850), .B(n_1851), .C(n_1852), .Y(n_1849) );
BUFx3_ASAP7_75t_L g1868 ( .A(n_1869), .Y(n_1868) );
INVx1_ASAP7_75t_L g1872 ( .A(n_1873), .Y(n_1872) );
endmodule