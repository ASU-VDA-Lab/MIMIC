module fake_jpeg_17684_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx11_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_0),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_21),
.A2(n_17),
.B1(n_11),
.B2(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_16),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_15),
.B(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_11),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_24),
.B1(n_22),
.B2(n_19),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_33),
.B1(n_10),
.B2(n_13),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_33),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_18),
.B1(n_12),
.B2(n_9),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_18),
.B1(n_9),
.B2(n_15),
.Y(n_41)
);

AO22x1_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_12),
.B1(n_13),
.B2(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_5),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_42),
.B1(n_36),
.B2(n_12),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_48),
.B(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_2),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_43),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_2),
.B(n_3),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_3),
.B(n_4),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_6),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_59),
.B(n_61),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_52),
.B(n_3),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_60),
.B1(n_48),
.B2(n_62),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_47),
.B(n_4),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_57),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_51),
.B(n_54),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_66),
.C(n_6),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_8),
.Y(n_71)
);


endmodule