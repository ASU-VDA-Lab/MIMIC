module fake_ariane_3362_n_1272 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_269, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_274, n_115, n_272, n_133, n_66, n_205, n_236, n_265, n_71, n_267, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_281, n_209, n_49, n_262, n_20, n_174, n_275, n_100, n_17, n_283, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_271, n_46, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_278, n_122, n_268, n_257, n_266, n_198, n_282, n_148, n_232, n_164, n_52, n_277, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_276, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_279, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_270, n_194, n_97, n_154, n_280, n_215, n_252, n_142, n_251, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_273, n_54, n_25, n_1272);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_269;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_274;
input n_115;
input n_272;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_267;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_281;
input n_209;
input n_49;
input n_262;
input n_20;
input n_174;
input n_275;
input n_100;
input n_17;
input n_283;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_271;
input n_46;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_278;
input n_122;
input n_268;
input n_257;
input n_266;
input n_198;
input n_282;
input n_148;
input n_232;
input n_164;
input n_52;
input n_277;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_276;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_279;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_270;
input n_194;
input n_97;
input n_154;
input n_280;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_273;
input n_54;
input n_25;

output n_1272;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1018;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_461;
wire n_1121;
wire n_490;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_1178;
wire n_1026;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_967;
wire n_1083;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_1015;
wire n_545;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_321;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_888;
wire n_845;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1266;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_1072;
wire n_695;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_617;
wire n_543;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_774;
wire n_933;
wire n_954;
wire n_596;
wire n_1168;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_203),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_243),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_200),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_182),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_90),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_109),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_2),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_152),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_145),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_13),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_271),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_102),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_222),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_259),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_262),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_223),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_193),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_16),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_214),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_167),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_111),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_184),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_246),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_149),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_88),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_177),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_235),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_57),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_8),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_128),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_194),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_27),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_75),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_62),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_142),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_114),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_266),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_96),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_121),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_212),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_36),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_198),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_175),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_218),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_8),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_34),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_147),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_199),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_183),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_7),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_71),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_164),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_207),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_260),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_70),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_155),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_89),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_132),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_2),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_170),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_49),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_44),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_112),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_75),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_248),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_161),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_279),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_92),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_40),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_54),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_126),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_80),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_270),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_174),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_245),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_261),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_168),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_190),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_71),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_61),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_18),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_125),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_202),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_51),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_263),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_159),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_73),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_46),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_116),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_216),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_41),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_156),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_141),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_181),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_80),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_242),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_81),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_11),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_255),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_256),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_187),
.Y(n_386)
);

BUFx2_ASAP7_75t_SL g387 ( 
.A(n_47),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_63),
.Y(n_388)
);

BUFx2_ASAP7_75t_SL g389 ( 
.A(n_25),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_213),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_211),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_144),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_26),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_27),
.Y(n_394)
);

BUFx10_ASAP7_75t_L g395 ( 
.A(n_120),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_12),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_47),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_231),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_232),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_74),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_237),
.Y(n_401)
);

BUFx10_ASAP7_75t_L g402 ( 
.A(n_153),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_79),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_138),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_250),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_133),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_278),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_146),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_56),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_252),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_206),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_179),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_54),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_189),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_229),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_221),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_143),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_99),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_118),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_276),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_4),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_178),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_60),
.Y(n_423)
);

BUFx10_ASAP7_75t_L g424 ( 
.A(n_38),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_241),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_195),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_13),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_244),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_5),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_91),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_137),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_165),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_21),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_32),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_257),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_104),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_131),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_254),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_40),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_129),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_93),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_95),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_124),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_64),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_283),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_53),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_108),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_173),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_247),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_267),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_30),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_139),
.Y(n_452)
);

BUFx5_ASAP7_75t_L g453 ( 
.A(n_269),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_61),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_38),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_134),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_220),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_277),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_123),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_172),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_39),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_204),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_23),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_106),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_264),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_197),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_192),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_275),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_113),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_226),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_157),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_176),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_86),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_274),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_135),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_140),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_127),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_272),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_282),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_296),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_299),
.B(n_0),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_355),
.B(n_0),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_355),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_290),
.B(n_1),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_326),
.B(n_349),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_296),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_401),
.B(n_1),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_314),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_344),
.B(n_3),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_386),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_290),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_296),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_316),
.B(n_3),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_289),
.B(n_4),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_433),
.B(n_5),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_306),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_357),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_306),
.Y(n_499)
);

BUFx8_ASAP7_75t_L g500 ( 
.A(n_298),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_386),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_357),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_436),
.B(n_6),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_395),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_319),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_331),
.Y(n_506)
);

BUFx12f_ASAP7_75t_L g507 ( 
.A(n_395),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_395),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_291),
.B(n_7),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_306),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_357),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_302),
.B(n_9),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_402),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_357),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_346),
.B(n_9),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_308),
.B(n_10),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_382),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_433),
.B(n_10),
.Y(n_518)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_354),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_402),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_402),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_461),
.Y(n_522)
);

BUFx12f_ASAP7_75t_L g523 ( 
.A(n_471),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_307),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_436),
.B(n_309),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_373),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_310),
.B(n_11),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_293),
.B(n_424),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_328),
.B(n_14),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_376),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_307),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_471),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_293),
.B(n_15),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_471),
.Y(n_534)
);

INVx5_ASAP7_75t_L g535 ( 
.A(n_307),
.Y(n_535)
);

BUFx12f_ASAP7_75t_L g536 ( 
.A(n_293),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_312),
.B(n_15),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_320),
.B(n_16),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_385),
.B(n_17),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_323),
.B(n_17),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_424),
.B(n_18),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_324),
.B(n_19),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_328),
.B(n_19),
.Y(n_543)
);

BUFx12f_ASAP7_75t_L g544 ( 
.A(n_424),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_307),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_380),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_374),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_382),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_374),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_383),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_381),
.Y(n_551)
);

BUFx8_ASAP7_75t_SL g552 ( 
.A(n_439),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_327),
.B(n_20),
.Y(n_553)
);

BUFx8_ASAP7_75t_L g554 ( 
.A(n_378),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_329),
.B(n_20),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_381),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_371),
.B(n_21),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_381),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_397),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_333),
.B(n_22),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_381),
.Y(n_561)
);

BUFx12f_ASAP7_75t_L g562 ( 
.A(n_301),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_371),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_377),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_403),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_427),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_454),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_315),
.B(n_22),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_473),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_377),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_438),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_334),
.B(n_23),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_313),
.Y(n_573)
);

BUFx8_ASAP7_75t_SL g574 ( 
.A(n_337),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_438),
.B(n_24),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_445),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_387),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_288),
.Y(n_578)
);

INVx6_ASAP7_75t_L g579 ( 
.A(n_457),
.Y(n_579)
);

CKINVDCx6p67_ASAP7_75t_R g580 ( 
.A(n_337),
.Y(n_580)
);

INVx6_ASAP7_75t_L g581 ( 
.A(n_453),
.Y(n_581)
);

BUFx12f_ASAP7_75t_L g582 ( 
.A(n_317),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_343),
.B(n_345),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_288),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_353),
.B(n_25),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_367),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_375),
.B(n_26),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_303),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_379),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_384),
.B(n_28),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_284),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_390),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_391),
.B(n_29),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_303),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_398),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_332),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_432),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_389),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_318),
.Y(n_599)
);

CKINVDCx11_ASAP7_75t_R g600 ( 
.A(n_399),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_407),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_409),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_408),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_414),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_416),
.B(n_417),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_430),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_472),
.B(n_29),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_440),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_472),
.B(n_31),
.Y(n_609)
);

NOR2x1_ASAP7_75t_L g610 ( 
.A(n_450),
.B(n_87),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_418),
.B(n_31),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_456),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_460),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_464),
.B(n_32),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_465),
.B(n_33),
.Y(n_615)
);

BUFx8_ASAP7_75t_SL g616 ( 
.A(n_410),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_468),
.B(n_33),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_SL g618 ( 
.A1(n_522),
.A2(n_411),
.B1(n_449),
.B2(n_410),
.Y(n_618)
);

AO22x2_ASAP7_75t_L g619 ( 
.A1(n_539),
.A2(n_489),
.B1(n_515),
.B2(n_568),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_611),
.A2(n_459),
.B1(n_419),
.B2(n_418),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_539),
.A2(n_419),
.B1(n_330),
.B2(n_336),
.Y(n_621)
);

AO22x2_ASAP7_75t_L g622 ( 
.A1(n_533),
.A2(n_352),
.B1(n_359),
.B2(n_304),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_528),
.A2(n_340),
.B1(n_347),
.B2(n_335),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_511),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_483),
.B(n_364),
.Y(n_625)
);

AO22x2_ASAP7_75t_L g626 ( 
.A1(n_541),
.A2(n_443),
.B1(n_475),
.B2(n_474),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_576),
.B(n_365),
.Y(n_627)
);

AND2x4_ASAP7_75t_SL g628 ( 
.A(n_580),
.B(n_476),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_576),
.B(n_366),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_490),
.B(n_285),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_521),
.B(n_369),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_578),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_511),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_490),
.B(n_491),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_579),
.A2(n_388),
.B1(n_393),
.B2(n_372),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_490),
.B(n_394),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_548),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_579),
.A2(n_400),
.B1(n_413),
.B2(n_396),
.Y(n_638)
);

OA22x2_ASAP7_75t_L g639 ( 
.A1(n_485),
.A2(n_423),
.B1(n_429),
.B2(n_421),
.Y(n_639)
);

OAI22xp33_ASAP7_75t_SL g640 ( 
.A1(n_481),
.A2(n_444),
.B1(n_446),
.B2(n_434),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_481),
.A2(n_455),
.B1(n_463),
.B2(n_451),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_491),
.B(n_286),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_491),
.B(n_287),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_501),
.B(n_292),
.Y(n_644)
);

AO22x2_ASAP7_75t_L g645 ( 
.A1(n_607),
.A2(n_609),
.B1(n_529),
.B2(n_557),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_571),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_L g647 ( 
.A1(n_487),
.A2(n_295),
.B1(n_297),
.B2(n_294),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_548),
.Y(n_648)
);

OAI22xp33_ASAP7_75t_L g649 ( 
.A1(n_487),
.A2(n_305),
.B1(n_311),
.B2(n_300),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_498),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_578),
.Y(n_651)
);

OAI22xp33_ASAP7_75t_L g652 ( 
.A1(n_494),
.A2(n_322),
.B1(n_325),
.B2(n_321),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_578),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_616),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_584),
.Y(n_655)
);

OA22x2_ASAP7_75t_L g656 ( 
.A1(n_602),
.A2(n_339),
.B1(n_341),
.B2(n_338),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_501),
.B(n_342),
.Y(n_657)
);

AO22x2_ASAP7_75t_L g658 ( 
.A1(n_607),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_658)
);

OA22x2_ASAP7_75t_L g659 ( 
.A1(n_546),
.A2(n_598),
.B1(n_577),
.B2(n_492),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_502),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_584),
.Y(n_661)
);

OR2x6_ASAP7_75t_L g662 ( 
.A(n_536),
.B(n_544),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_529),
.A2(n_350),
.B1(n_351),
.B2(n_348),
.Y(n_663)
);

OR2x6_ASAP7_75t_L g664 ( 
.A(n_504),
.B(n_35),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_514),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_584),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_591),
.B(n_356),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_501),
.B(n_358),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_543),
.A2(n_361),
.B1(n_362),
.B2(n_360),
.Y(n_669)
);

OAI22xp33_ASAP7_75t_SL g670 ( 
.A1(n_583),
.A2(n_479),
.B1(n_478),
.B2(n_477),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_SL g671 ( 
.A1(n_519),
.A2(n_470),
.B1(n_469),
.B2(n_467),
.Y(n_671)
);

OA22x2_ASAP7_75t_L g672 ( 
.A1(n_546),
.A2(n_466),
.B1(n_462),
.B2(n_458),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_488),
.Y(n_673)
);

INVx8_ASAP7_75t_L g674 ( 
.A(n_507),
.Y(n_674)
);

AO22x2_ASAP7_75t_L g675 ( 
.A1(n_609),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_517),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_543),
.A2(n_406),
.B1(n_452),
.B2(n_448),
.Y(n_677)
);

AO22x2_ASAP7_75t_L g678 ( 
.A1(n_557),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_SL g679 ( 
.A1(n_523),
.A2(n_363),
.B1(n_368),
.B2(n_370),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_508),
.A2(n_520),
.B1(n_532),
.B2(n_513),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_508),
.A2(n_520),
.B1(n_532),
.B2(n_513),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_SL g682 ( 
.A1(n_583),
.A2(n_530),
.B1(n_495),
.B2(n_512),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_480),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_505),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_480),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_506),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_508),
.B(n_392),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_513),
.B(n_520),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_SL g689 ( 
.A1(n_509),
.A2(n_404),
.B1(n_405),
.B2(n_412),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_480),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_594),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_L g692 ( 
.A1(n_532),
.A2(n_415),
.B1(n_420),
.B2(n_422),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_591),
.B(n_425),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_600),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_534),
.B(n_426),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_575),
.A2(n_428),
.B1(n_431),
.B2(n_435),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_534),
.B(n_437),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_575),
.A2(n_447),
.B1(n_442),
.B2(n_441),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_534),
.B(n_453),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_594),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_614),
.A2(n_617),
.B1(n_615),
.B2(n_599),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_592),
.B(n_453),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_614),
.B(n_453),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_673),
.Y(n_704)
);

OR2x6_ASAP7_75t_L g705 ( 
.A(n_674),
.B(n_562),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_SL g706 ( 
.A(n_674),
.B(n_582),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_682),
.B(n_573),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_684),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_618),
.B(n_574),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_686),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_631),
.B(n_603),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_624),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_633),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_637),
.Y(n_714)
);

INVxp67_ASAP7_75t_SL g715 ( 
.A(n_648),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_632),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_632),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_651),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_651),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_653),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_646),
.B(n_482),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_655),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_655),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_627),
.B(n_525),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_661),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_661),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_666),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_645),
.B(n_605),
.Y(n_728)
);

AND2x2_ASAP7_75t_SL g729 ( 
.A(n_621),
.B(n_615),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_634),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_666),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_645),
.B(n_702),
.Y(n_732)
);

XNOR2xp5_ASAP7_75t_L g733 ( 
.A(n_694),
.B(n_552),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_691),
.Y(n_734)
);

OAI21xp5_ASAP7_75t_L g735 ( 
.A1(n_703),
.A2(n_516),
.B(n_512),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_691),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_700),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_700),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_650),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_660),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_636),
.B(n_606),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_665),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_676),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_625),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_679),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_685),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_690),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_629),
.B(n_667),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_634),
.B(n_482),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_699),
.Y(n_750)
);

XOR2xp5_ASAP7_75t_L g751 ( 
.A(n_654),
.B(n_620),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_659),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_683),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_701),
.B(n_484),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_683),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_683),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_688),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_663),
.A2(n_527),
.B(n_516),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_643),
.B(n_605),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_644),
.Y(n_760)
);

BUFx6f_ASAP7_75t_SL g761 ( 
.A(n_662),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_693),
.B(n_696),
.Y(n_762)
);

XNOR2x2_ASAP7_75t_L g763 ( 
.A(n_622),
.B(n_537),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_657),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_668),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_695),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_623),
.B(n_586),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_697),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_656),
.Y(n_769)
);

BUFx8_ASAP7_75t_L g770 ( 
.A(n_678),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_639),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_669),
.B(n_500),
.Y(n_772)
);

BUFx12f_ASAP7_75t_L g773 ( 
.A(n_662),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_672),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_677),
.B(n_500),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_698),
.B(n_554),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_SL g777 ( 
.A(n_671),
.B(n_484),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_628),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_630),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_642),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_687),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_647),
.B(n_617),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_716),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_738),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_711),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_717),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_754),
.B(n_664),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_724),
.B(n_619),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_753),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_718),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_754),
.B(n_619),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_719),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_767),
.B(n_658),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_759),
.B(n_658),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_720),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_759),
.B(n_758),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_748),
.B(n_762),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_722),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_704),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_723),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_758),
.B(n_675),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_728),
.B(n_675),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_725),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_726),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_779),
.B(n_635),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_780),
.B(n_638),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_735),
.A2(n_610),
.B(n_538),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_777),
.B(n_670),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_727),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_728),
.B(n_678),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_732),
.B(n_664),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_781),
.B(n_626),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_708),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_731),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_749),
.B(n_641),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_729),
.B(n_622),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_764),
.B(n_649),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_710),
.Y(n_818)
);

AND2x2_ASAP7_75t_SL g819 ( 
.A(n_729),
.B(n_496),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_734),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_721),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_765),
.B(n_652),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_741),
.B(n_496),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_736),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_737),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_715),
.B(n_554),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_744),
.B(n_707),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_739),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_740),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_743),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_742),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_735),
.B(n_760),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_742),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_766),
.B(n_518),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_705),
.B(n_752),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_707),
.B(n_589),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_768),
.B(n_692),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_712),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_713),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_750),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_730),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_755),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_778),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_782),
.B(n_527),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_714),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_732),
.B(n_595),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_769),
.B(n_601),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_774),
.B(n_550),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_771),
.B(n_526),
.Y(n_849)
);

BUFx4f_ASAP7_75t_L g850 ( 
.A(n_757),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_782),
.A2(n_503),
.B1(n_542),
.B2(n_537),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_705),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_772),
.B(n_550),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_746),
.Y(n_854)
);

INVxp33_ASAP7_75t_L g855 ( 
.A(n_751),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_756),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_772),
.B(n_565),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_775),
.B(n_565),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_775),
.B(n_567),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_747),
.A2(n_503),
.B(n_540),
.Y(n_860)
);

AND2x2_ASAP7_75t_SL g861 ( 
.A(n_776),
.B(n_553),
.Y(n_861)
);

BUFx12f_ASAP7_75t_L g862 ( 
.A(n_773),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_733),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_814),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_798),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_862),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_798),
.Y(n_867)
);

AND2x6_ASAP7_75t_L g868 ( 
.A(n_801),
.B(n_770),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_791),
.B(n_745),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_791),
.B(n_559),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_797),
.B(n_709),
.Y(n_871)
);

INVx5_ASAP7_75t_L g872 ( 
.A(n_814),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_785),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_862),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_814),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_821),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_798),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_788),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_783),
.Y(n_879)
);

OR2x6_ASAP7_75t_L g880 ( 
.A(n_787),
.B(n_761),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_783),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_SL g882 ( 
.A(n_819),
.B(n_706),
.Y(n_882)
);

INVxp67_ASAP7_75t_SL g883 ( 
.A(n_831),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_804),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_790),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_787),
.B(n_566),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_805),
.Y(n_887)
);

OR2x6_ASAP7_75t_L g888 ( 
.A(n_787),
.B(n_761),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_794),
.B(n_567),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_804),
.Y(n_890)
);

AND2x2_ASAP7_75t_SL g891 ( 
.A(n_819),
.B(n_763),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_796),
.B(n_604),
.Y(n_892)
);

AND2x2_ASAP7_75t_SL g893 ( 
.A(n_819),
.B(n_553),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_852),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_804),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_796),
.B(n_608),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_793),
.B(n_680),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_841),
.B(n_569),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_814),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_790),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_SL g901 ( 
.A(n_861),
.B(n_681),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_792),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_820),
.Y(n_903)
);

BUFx12f_ASAP7_75t_L g904 ( 
.A(n_835),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_799),
.B(n_813),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_863),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_792),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_814),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_789),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_827),
.B(n_563),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_789),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_844),
.B(n_689),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_832),
.B(n_594),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_833),
.B(n_597),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_815),
.Y(n_915)
);

CKINVDCx6p67_ASAP7_75t_R g916 ( 
.A(n_843),
.Y(n_916)
);

BUFx4f_ASAP7_75t_L g917 ( 
.A(n_835),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_855),
.B(n_555),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_784),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_789),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_841),
.B(n_849),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_795),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_811),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_841),
.B(n_612),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_799),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_789),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_921),
.B(n_923),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_879),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_916),
.Y(n_929)
);

NAND2x1p5_ASAP7_75t_L g930 ( 
.A(n_872),
.B(n_799),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_918),
.Y(n_931)
);

BUFx12f_ASAP7_75t_L g932 ( 
.A(n_866),
.Y(n_932)
);

INVx6_ASAP7_75t_SL g933 ( 
.A(n_880),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_874),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_874),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_894),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_872),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_875),
.Y(n_938)
);

INVx1_ASAP7_75t_SL g939 ( 
.A(n_894),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_919),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_872),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_866),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_887),
.B(n_915),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_875),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_925),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_872),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_881),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_875),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_885),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_904),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_865),
.Y(n_951)
);

BUFx8_ASAP7_75t_L g952 ( 
.A(n_886),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_905),
.Y(n_953)
);

INVx3_ASAP7_75t_SL g954 ( 
.A(n_906),
.Y(n_954)
);

INVx5_ASAP7_75t_L g955 ( 
.A(n_925),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_917),
.Y(n_956)
);

INVx5_ASAP7_75t_L g957 ( 
.A(n_926),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_869),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_900),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_905),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_891),
.A2(n_816),
.B1(n_808),
.B2(n_810),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_867),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_926),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_909),
.Y(n_964)
);

CKINVDCx11_ASAP7_75t_R g965 ( 
.A(n_880),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_902),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_886),
.B(n_853),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_907),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_926),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_871),
.A2(n_806),
.B1(n_811),
.B2(n_857),
.Y(n_970)
);

INVx8_ASAP7_75t_L g971 ( 
.A(n_888),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_893),
.B(n_857),
.Y(n_972)
);

BUFx2_ASAP7_75t_SL g973 ( 
.A(n_870),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_917),
.Y(n_974)
);

INVx8_ASAP7_75t_L g975 ( 
.A(n_888),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_893),
.B(n_858),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_909),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_878),
.B(n_813),
.Y(n_978)
);

BUFx12f_ASAP7_75t_L g979 ( 
.A(n_906),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_877),
.Y(n_980)
);

INVx6_ASAP7_75t_L g981 ( 
.A(n_924),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_922),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_926),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_864),
.B(n_813),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_958),
.A2(n_891),
.B1(n_816),
.B2(n_882),
.Y(n_985)
);

CKINVDCx8_ASAP7_75t_R g986 ( 
.A(n_973),
.Y(n_986)
);

INVx6_ASAP7_75t_L g987 ( 
.A(n_952),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_928),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_947),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_946),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_951),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_949),
.Y(n_992)
);

CKINVDCx11_ASAP7_75t_R g993 ( 
.A(n_936),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_931),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_951),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_972),
.B(n_883),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_957),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_959),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_966),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_962),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_968),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_962),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_976),
.A2(n_901),
.B1(n_812),
.B2(n_859),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_961),
.A2(n_859),
.B1(n_858),
.B2(n_811),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_961),
.A2(n_811),
.B1(n_818),
.B2(n_868),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_SL g1006 ( 
.A1(n_952),
.A2(n_802),
.B1(n_868),
.B2(n_912),
.Y(n_1006)
);

CKINVDCx11_ASAP7_75t_R g1007 ( 
.A(n_936),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_SL g1008 ( 
.A1(n_952),
.A2(n_868),
.B1(n_912),
.B2(n_640),
.Y(n_1008)
);

BUFx4f_ASAP7_75t_L g1009 ( 
.A(n_932),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_943),
.B(n_873),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_934),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_967),
.A2(n_818),
.B1(n_868),
.B2(n_898),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_980),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_982),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_957),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_978),
.B(n_883),
.Y(n_1016)
);

INVx6_ASAP7_75t_L g1017 ( 
.A(n_971),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_942),
.Y(n_1018)
);

INVx6_ASAP7_75t_L g1019 ( 
.A(n_971),
.Y(n_1019)
);

CKINVDCx11_ASAP7_75t_R g1020 ( 
.A(n_942),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_940),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_970),
.A2(n_851),
.B1(n_896),
.B2(n_892),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_934),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_SL g1024 ( 
.A1(n_939),
.A2(n_851),
.B(n_560),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_971),
.B(n_975),
.Y(n_1025)
);

INVx5_ASAP7_75t_SL g1026 ( 
.A(n_927),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_940),
.Y(n_1027)
);

OAI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_954),
.A2(n_850),
.B1(n_896),
.B2(n_892),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_978),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_946),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_965),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_927),
.Y(n_1032)
);

INVx6_ASAP7_75t_L g1033 ( 
.A(n_975),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_927),
.Y(n_1034)
);

OAI22xp33_ASAP7_75t_R g1035 ( 
.A1(n_979),
.A2(n_560),
.B1(n_572),
.B2(n_542),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_981),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_979),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_960),
.B(n_884),
.Y(n_1038)
);

OAI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_932),
.A2(n_850),
.B1(n_876),
.B2(n_826),
.Y(n_1039)
);

INVx6_ASAP7_75t_L g1040 ( 
.A(n_975),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_981),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_960),
.B(n_890),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_1035),
.A2(n_836),
.B1(n_828),
.B2(n_910),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_988),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_1022),
.A2(n_840),
.B1(n_800),
.B2(n_824),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_1011),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1029),
.B(n_807),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_1032),
.B(n_1034),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1022),
.A2(n_840),
.B1(n_803),
.B2(n_825),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_1023),
.Y(n_1050)
);

BUFx4f_ASAP7_75t_SL g1051 ( 
.A(n_1018),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_1016),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_991),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_997),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_989),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_1028),
.B(n_955),
.Y(n_1056)
);

OAI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_1024),
.A2(n_585),
.B(n_572),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_1008),
.A2(n_830),
.B1(n_839),
.B2(n_829),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_985),
.A2(n_829),
.B1(n_786),
.B2(n_846),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_997),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_993),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_992),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1016),
.B(n_807),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_1007),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_995),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_1025),
.Y(n_1066)
);

CKINVDCx6p67_ASAP7_75t_R g1067 ( 
.A(n_1020),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_996),
.A2(n_1003),
.B1(n_1004),
.B2(n_1026),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_998),
.B(n_889),
.Y(n_1069)
);

BUFx4f_ASAP7_75t_SL g1070 ( 
.A(n_1031),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_999),
.B(n_964),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_1025),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_1039),
.B(n_955),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_SL g1074 ( 
.A1(n_987),
.A2(n_974),
.B1(n_817),
.B2(n_822),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1026),
.A2(n_840),
.B1(n_824),
.B2(n_825),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1000),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_1005),
.A2(n_1006),
.B1(n_1012),
.B2(n_994),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1002),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1001),
.B(n_964),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_SL g1080 ( 
.A1(n_1026),
.A2(n_950),
.B1(n_956),
.B2(n_929),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1010),
.B(n_935),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_1025),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_986),
.A2(n_809),
.B1(n_945),
.B2(n_955),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1013),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_SL g1085 ( 
.A1(n_1037),
.A2(n_935),
.B1(n_837),
.B2(n_950),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_SL g1086 ( 
.A1(n_1017),
.A2(n_953),
.B1(n_823),
.B2(n_590),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1027),
.A2(n_838),
.B1(n_903),
.B2(n_895),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1014),
.B(n_1021),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1009),
.A2(n_809),
.B1(n_984),
.B2(n_899),
.Y(n_1089)
);

AOI222xp33_ASAP7_75t_L g1090 ( 
.A1(n_1057),
.A2(n_587),
.B1(n_593),
.B2(n_834),
.C1(n_845),
.C2(n_860),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1052),
.B(n_1041),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1085),
.A2(n_1019),
.B1(n_1033),
.B2(n_1017),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_1058),
.A2(n_784),
.B1(n_854),
.B2(n_933),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1068),
.A2(n_933),
.B1(n_845),
.B2(n_1036),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1043),
.A2(n_933),
.B1(n_1042),
.B2(n_1038),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1059),
.A2(n_564),
.B1(n_570),
.B2(n_612),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1063),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1063),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1077),
.A2(n_564),
.B1(n_570),
.B2(n_612),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1086),
.A2(n_984),
.B1(n_864),
.B2(n_908),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1074),
.A2(n_570),
.B1(n_613),
.B2(n_833),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1069),
.B(n_990),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1044),
.Y(n_1103)
);

OAI22x1_ASAP7_75t_L g1104 ( 
.A1(n_1055),
.A2(n_849),
.B1(n_930),
.B2(n_948),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1088),
.B(n_1030),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1045),
.A2(n_1040),
.B1(n_930),
.B2(n_809),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1049),
.A2(n_1015),
.B1(n_948),
.B2(n_946),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1088),
.B(n_977),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1048),
.A2(n_1053),
.B1(n_1076),
.B2(n_1065),
.Y(n_1109)
);

OAI22x1_ASAP7_75t_L g1110 ( 
.A1(n_1062),
.A2(n_849),
.B1(n_1015),
.B2(n_897),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1071),
.B(n_977),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1048),
.A2(n_1053),
.B1(n_1076),
.B2(n_1065),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1078),
.A2(n_914),
.B1(n_913),
.B2(n_789),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1075),
.A2(n_937),
.B1(n_941),
.B2(n_957),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1056),
.B(n_983),
.Y(n_1115)
);

OA21x2_ASAP7_75t_L g1116 ( 
.A1(n_1056),
.A2(n_913),
.B(n_847),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1078),
.A2(n_849),
.B1(n_847),
.B2(n_596),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1081),
.A2(n_944),
.B1(n_938),
.B2(n_963),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1080),
.A2(n_944),
.B1(n_938),
.B2(n_963),
.Y(n_1119)
);

OAI222xp33_ASAP7_75t_L g1120 ( 
.A1(n_1073),
.A2(n_588),
.B1(n_848),
.B2(n_842),
.C1(n_856),
.C2(n_558),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1084),
.A2(n_842),
.B1(n_856),
.B2(n_920),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1087),
.A2(n_909),
.B1(n_911),
.B2(n_920),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1071),
.B(n_938),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1073),
.A2(n_911),
.B1(n_944),
.B2(n_963),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_1079),
.A2(n_911),
.B1(n_969),
.B2(n_963),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_SL g1126 ( 
.A1(n_1066),
.A2(n_983),
.B1(n_969),
.B2(n_453),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1047),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1066),
.A2(n_983),
.B1(n_969),
.B2(n_581),
.Y(n_1128)
);

OAI222xp33_ASAP7_75t_L g1129 ( 
.A1(n_1089),
.A2(n_510),
.B1(n_551),
.B2(n_46),
.C1(n_48),
.C2(n_50),
.Y(n_1129)
);

AOI221xp5_ASAP7_75t_L g1130 ( 
.A1(n_1046),
.A2(n_486),
.B1(n_493),
.B2(n_497),
.C(n_499),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_SL g1131 ( 
.A1(n_1083),
.A2(n_45),
.B(n_51),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1054),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1066),
.A2(n_486),
.B1(n_556),
.B2(n_549),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1051),
.A2(n_1067),
.B1(n_1061),
.B2(n_1064),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1072),
.A2(n_497),
.B1(n_556),
.B2(n_549),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1046),
.B(n_45),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1097),
.B(n_1050),
.Y(n_1137)
);

AOI221xp5_ASAP7_75t_L g1138 ( 
.A1(n_1129),
.A2(n_1050),
.B1(n_1064),
.B2(n_497),
.C(n_531),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_SL g1139 ( 
.A1(n_1116),
.A2(n_1082),
.B1(n_1072),
.B2(n_1070),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1131),
.A2(n_1060),
.B1(n_1054),
.B2(n_1082),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1103),
.B(n_1105),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_L g1142 ( 
.A(n_1090),
.B(n_1060),
.C(n_1072),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1102),
.B(n_52),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1108),
.B(n_52),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1091),
.B(n_55),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1098),
.B(n_58),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_SL g1147 ( 
.A1(n_1134),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1127),
.B(n_59),
.Y(n_1148)
);

NOR3xp33_ASAP7_75t_SL g1149 ( 
.A(n_1136),
.B(n_63),
.C(n_64),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1115),
.B(n_524),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1111),
.B(n_65),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1123),
.B(n_66),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_1132),
.B(n_561),
.C(n_545),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_L g1154 ( 
.A1(n_1110),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.C(n_69),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_R g1155 ( 
.A(n_1124),
.B(n_69),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1092),
.B(n_561),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1118),
.B(n_72),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1125),
.B(n_74),
.Y(n_1158)
);

AOI221xp5_ASAP7_75t_L g1159 ( 
.A1(n_1110),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.C(n_79),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1109),
.B(n_78),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1119),
.B(n_561),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1112),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1116),
.B(n_81),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1094),
.B(n_82),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1095),
.B(n_82),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1104),
.B(n_83),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1106),
.B(n_535),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1104),
.B(n_84),
.Y(n_1168)
);

AOI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_1099),
.A2(n_1101),
.B1(n_1100),
.B2(n_1093),
.C(n_1117),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1120),
.A2(n_85),
.B(n_86),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1162),
.A2(n_1096),
.B1(n_1122),
.B2(n_1113),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1141),
.B(n_1107),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1137),
.B(n_1114),
.Y(n_1173)
);

NAND4xp75_ASAP7_75t_L g1174 ( 
.A(n_1149),
.B(n_1130),
.C(n_1126),
.D(n_1128),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1145),
.B(n_1121),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1163),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1146),
.B(n_1133),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1139),
.B(n_1135),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1148),
.B(n_94),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_1143),
.B(n_97),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1166),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1168),
.Y(n_1182)
);

AND2x2_ASAP7_75t_SL g1183 ( 
.A(n_1154),
.B(n_98),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1152),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1150),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1144),
.B(n_1151),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1150),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_1160),
.B(n_100),
.Y(n_1188)
);

NAND4xp75_ASAP7_75t_L g1189 ( 
.A(n_1138),
.B(n_101),
.C(n_103),
.D(n_105),
.Y(n_1189)
);

NOR3xp33_ASAP7_75t_L g1190 ( 
.A(n_1147),
.B(n_107),
.C(n_110),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1142),
.B(n_115),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1170),
.A2(n_547),
.B1(n_119),
.B2(n_122),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1140),
.B(n_117),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1167),
.B(n_130),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_1182),
.Y(n_1195)
);

NAND4xp75_ASAP7_75t_L g1196 ( 
.A(n_1183),
.B(n_1159),
.C(n_1164),
.D(n_1156),
.Y(n_1196)
);

NAND4xp75_ASAP7_75t_L g1197 ( 
.A(n_1183),
.B(n_1158),
.C(n_1165),
.D(n_1157),
.Y(n_1197)
);

NAND4xp75_ASAP7_75t_L g1198 ( 
.A(n_1192),
.B(n_1161),
.C(n_1169),
.D(n_1155),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1176),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1181),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_1182),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1181),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1172),
.B(n_1173),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1172),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1184),
.B(n_1153),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_1179),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1185),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1201),
.A2(n_1186),
.B1(n_1175),
.B2(n_1193),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1201),
.Y(n_1209)
);

INVxp67_ASAP7_75t_L g1210 ( 
.A(n_1195),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1202),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1200),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1204),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1200),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1203),
.Y(n_1215)
);

XOR2x2_ASAP7_75t_L g1216 ( 
.A(n_1197),
.B(n_1190),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1206),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1206),
.B(n_1180),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1207),
.Y(n_1219)
);

XOR2x2_ASAP7_75t_L g1220 ( 
.A(n_1198),
.B(n_1191),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1199),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1199),
.Y(n_1222)
);

NOR2x1_ASAP7_75t_L g1223 ( 
.A(n_1206),
.B(n_1205),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1213),
.Y(n_1224)
);

INVxp67_ASAP7_75t_L g1225 ( 
.A(n_1218),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1215),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1223),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1215),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1209),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1211),
.Y(n_1230)
);

AOI22x1_ASAP7_75t_L g1231 ( 
.A1(n_1208),
.A2(n_1188),
.B1(n_1194),
.B2(n_1196),
.Y(n_1231)
);

AOI22x1_ASAP7_75t_L g1232 ( 
.A1(n_1217),
.A2(n_1216),
.B1(n_1210),
.B2(n_1220),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1219),
.Y(n_1233)
);

AOI22x1_ASAP7_75t_L g1234 ( 
.A1(n_1210),
.A2(n_1194),
.B1(n_1196),
.B2(n_1177),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1224),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_SL g1236 ( 
.A(n_1229),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1230),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1233),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1234),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1226),
.Y(n_1240)
);

OAI322xp33_ASAP7_75t_L g1241 ( 
.A1(n_1232),
.A2(n_1222),
.A3(n_1221),
.B1(n_1214),
.B2(n_1212),
.C1(n_1187),
.C2(n_1178),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1228),
.Y(n_1242)
);

OA22x2_ASAP7_75t_SL g1243 ( 
.A1(n_1239),
.A2(n_1234),
.B1(n_1232),
.B2(n_1231),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1236),
.A2(n_1225),
.B1(n_1227),
.B2(n_1222),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1235),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1237),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1242),
.A2(n_1174),
.B1(n_1189),
.B2(n_1171),
.Y(n_1247)
);

AOI32xp33_ASAP7_75t_L g1248 ( 
.A1(n_1243),
.A2(n_1242),
.A3(n_1241),
.B1(n_1240),
.B2(n_1238),
.Y(n_1248)
);

AO22x2_ASAP7_75t_L g1249 ( 
.A1(n_1244),
.A2(n_136),
.B1(n_148),
.B2(n_150),
.Y(n_1249)
);

NOR4xp25_ASAP7_75t_L g1250 ( 
.A(n_1245),
.B(n_151),
.C(n_154),
.D(n_158),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_SL g1251 ( 
.A1(n_1246),
.A2(n_160),
.B(n_162),
.C(n_163),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1247),
.A2(n_166),
.B1(n_169),
.B2(n_171),
.Y(n_1252)
);

NOR4xp25_ASAP7_75t_L g1253 ( 
.A(n_1248),
.B(n_180),
.C(n_185),
.D(n_186),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1252),
.A2(n_188),
.B1(n_191),
.B2(n_196),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1250),
.A2(n_1249),
.B1(n_1251),
.B2(n_201),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1253),
.B(n_205),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1255),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1256),
.A2(n_1254),
.B1(n_208),
.B2(n_209),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1258),
.Y(n_1259)
);

OR3x2_ASAP7_75t_L g1260 ( 
.A(n_1258),
.B(n_1257),
.C(n_210),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1260),
.A2(n_215),
.B1(n_217),
.B2(n_219),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1259),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1261),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1262),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1263),
.A2(n_281),
.B1(n_228),
.B2(n_230),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1264),
.A2(n_233),
.B1(n_234),
.B2(n_236),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1266),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1265),
.Y(n_1268)
);

AO22x2_ASAP7_75t_L g1269 ( 
.A1(n_1267),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1269),
.Y(n_1270)
);

AOI221xp5_ASAP7_75t_L g1271 ( 
.A1(n_1270),
.A2(n_1268),
.B1(n_249),
.B2(n_251),
.C(n_253),
.Y(n_1271)
);

AOI211xp5_ASAP7_75t_L g1272 ( 
.A1(n_1271),
.A2(n_258),
.B(n_273),
.C(n_280),
.Y(n_1272)
);


endmodule