module real_aes_11860_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_0), .Y(n_545) );
INVx1_ASAP7_75t_L g137 ( .A(n_1), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_2), .Y(n_607) );
AND2x2_ASAP7_75t_L g561 ( .A(n_3), .B(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_3), .Y(n_589) );
INVx1_ASAP7_75t_L g601 ( .A(n_3), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_3), .B(n_62), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_4), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_5), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_6), .B(n_157), .Y(n_230) );
INVx2_ASAP7_75t_L g491 ( .A(n_7), .Y(n_491) );
OR2x2_ASAP7_75t_L g642 ( .A(n_7), .B(n_542), .Y(n_642) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_8), .Y(n_670) );
BUFx2_ASAP7_75t_L g493 ( .A(n_9), .Y(n_493) );
BUFx2_ASAP7_75t_L g529 ( .A(n_9), .Y(n_529) );
INVx1_ASAP7_75t_L g544 ( .A(n_9), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_10), .A2(n_37), .B1(n_508), .B2(n_514), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g581 ( .A1(n_10), .A2(n_37), .B1(n_582), .B2(n_585), .C(n_588), .Y(n_581) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_11), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_12), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_13), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_14), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_15), .A2(n_75), .B1(n_525), .B2(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g559 ( .A(n_15), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_16), .B(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_17), .B(n_122), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_18), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_19), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_20), .B(n_115), .Y(n_200) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_21), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_22), .B(n_117), .Y(n_116) );
AO221x1_ASAP7_75t_L g594 ( .A1(n_23), .A2(n_28), .B1(n_595), .B2(n_597), .C(n_598), .Y(n_594) );
INVx1_ASAP7_75t_L g643 ( .A(n_23), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_24), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_25), .B(n_122), .Y(n_229) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_26), .Y(n_90) );
OAI21xp33_ASAP7_75t_L g179 ( .A1(n_27), .A2(n_92), .B(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g651 ( .A(n_28), .Y(n_651) );
INVx1_ASAP7_75t_L g490 ( .A(n_29), .Y(n_490) );
INVx1_ASAP7_75t_L g542 ( .A(n_29), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_30), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_31), .B(n_115), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_32), .Y(n_166) );
XNOR2xp5_ASAP7_75t_L g480 ( .A(n_33), .B(n_481), .Y(n_480) );
OAI21x1_ASAP7_75t_L g110 ( .A1(n_34), .A2(n_56), .B(n_111), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_35), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_36), .B(n_115), .Y(n_114) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_36), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_38), .Y(n_244) );
AND2x6_ASAP7_75t_L g83 ( .A(n_39), .B(n_84), .Y(n_83) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_39), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_39), .B(n_660), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_40), .A2(n_66), .B1(n_157), .B2(n_182), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_41), .A2(n_57), .B1(n_518), .B2(n_521), .Y(n_517) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_41), .A2(n_594), .B1(n_602), .B2(n_611), .C(n_614), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_42), .A2(n_65), .B1(n_495), .B2(n_500), .Y(n_494) );
AOI22xp33_ASAP7_75t_SL g578 ( .A1(n_42), .A2(n_65), .B1(n_579), .B2(n_580), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_43), .B(n_170), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_44), .Y(n_159) );
INVx1_ASAP7_75t_L g84 ( .A(n_45), .Y(n_84) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_45), .Y(n_660) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_46), .Y(n_208) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_47), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_48), .B(n_182), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_49), .B(n_182), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_50), .B(n_128), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_51), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_52), .B(n_170), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_53), .B(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g148 ( .A(n_54), .Y(n_148) );
INVx2_ASAP7_75t_L g568 ( .A(n_55), .Y(n_568) );
INVx1_ASAP7_75t_L g591 ( .A(n_57), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g124 ( .A(n_58), .B(n_123), .Y(n_124) );
INVx1_ASAP7_75t_L g141 ( .A(n_59), .Y(n_141) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_59), .Y(n_696) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_60), .Y(n_252) );
BUFx10_ASAP7_75t_L g691 ( .A(n_61), .Y(n_691) );
INVx2_ASAP7_75t_L g562 ( .A(n_62), .Y(n_562) );
INVx1_ASAP7_75t_L g246 ( .A(n_63), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_64), .B(n_123), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_67), .B(n_170), .Y(n_202) );
INVx1_ASAP7_75t_L g150 ( .A(n_68), .Y(n_150) );
INVx2_ASAP7_75t_L g111 ( .A(n_69), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_70), .Y(n_678) );
NOR2xp67_ASAP7_75t_L g176 ( .A(n_71), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g565 ( .A(n_72), .Y(n_565) );
BUFx3_ASAP7_75t_L g499 ( .A(n_73), .Y(n_499) );
INVx1_ASAP7_75t_L g506 ( .A(n_73), .Y(n_506) );
INVx1_ASAP7_75t_L g498 ( .A(n_74), .Y(n_498) );
BUFx3_ASAP7_75t_L g505 ( .A(n_74), .Y(n_505) );
INVx1_ASAP7_75t_L g569 ( .A(n_75), .Y(n_569) );
NAND2xp33_ASAP7_75t_L g204 ( .A(n_76), .B(n_170), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_94), .B(n_479), .Y(n_77) );
BUFx2_ASAP7_75t_SL g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_85), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx2_ASAP7_75t_SL g126 ( .A(n_82), .Y(n_126) );
INVx8_ASAP7_75t_L g183 ( .A(n_82), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_82), .A2(n_128), .B(n_254), .Y(n_253) );
INVx8_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
AOI21xp33_ASAP7_75t_L g151 ( .A1(n_83), .A2(n_129), .B(n_149), .Y(n_151) );
INVx1_ASAP7_75t_L g163 ( .A(n_83), .Y(n_163) );
INVx1_ASAP7_75t_L g215 ( .A(n_83), .Y(n_215) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
AO21x1_ASAP7_75t_L g706 ( .A1(n_86), .A2(n_707), .B(n_708), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_87), .B(n_91), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx2_ASAP7_75t_L g146 ( .A(n_89), .Y(n_146) );
INVx2_ASAP7_75t_L g178 ( .A(n_89), .Y(n_178) );
INVx2_ASAP7_75t_L g180 ( .A(n_89), .Y(n_180) );
INVx2_ASAP7_75t_L g182 ( .A(n_89), .Y(n_182) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_90), .Y(n_118) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_90), .Y(n_123) );
INVx2_ASAP7_75t_L g158 ( .A(n_90), .Y(n_158) );
INVx1_ASAP7_75t_L g243 ( .A(n_90), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_91), .A2(n_144), .B(n_149), .Y(n_143) );
AO21x1_ASAP7_75t_L g239 ( .A1(n_91), .A2(n_240), .B(n_245), .Y(n_239) );
AOI21x1_ASAP7_75t_L g247 ( .A1(n_91), .A2(n_248), .B(n_250), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_92), .Y(n_91) );
BUFx2_ASAP7_75t_L g142 ( .A(n_92), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_92), .B(n_165), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_92), .A2(n_176), .B1(n_179), .B2(n_181), .Y(n_175) );
INVx3_ASAP7_75t_L g227 ( .A(n_92), .Y(n_227) );
BUFx12f_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx5_ASAP7_75t_L g119 ( .A(n_93), .Y(n_119) );
INVx5_ASAP7_75t_L g155 ( .A(n_93), .Y(n_155) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx3_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
NAND4xp75_ASAP7_75t_L g98 ( .A(n_99), .B(n_338), .C(n_393), .D(n_440), .Y(n_98) );
NOR2x1_ASAP7_75t_L g99 ( .A(n_100), .B(n_288), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g100 ( .A(n_101), .B(n_267), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_187), .B1(n_233), .B2(n_255), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_130), .Y(n_103) );
AND2x2_ASAP7_75t_L g273 ( .A(n_104), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g313 ( .A(n_104), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g327 ( .A(n_104), .B(n_260), .Y(n_327) );
INVx2_ASAP7_75t_L g344 ( .A(n_104), .Y(n_344) );
INVx2_ASAP7_75t_L g404 ( .A(n_104), .Y(n_404) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g258 ( .A(n_105), .B(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g266 ( .A(n_105), .B(n_173), .Y(n_266) );
BUFx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g325 ( .A(n_106), .Y(n_325) );
OAI21x1_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_112), .B(n_127), .Y(n_106) );
OAI21x1_ASAP7_75t_SL g221 ( .A1(n_107), .A2(n_222), .B(n_232), .Y(n_221) );
BUFx4f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_108), .B(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g192 ( .A(n_108), .Y(n_192) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g129 ( .A(n_109), .Y(n_129) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g171 ( .A(n_110), .Y(n_171) );
OAI21x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_120), .B(n_126), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_116), .B(n_119), .Y(n_113) );
INVx2_ASAP7_75t_L g139 ( .A(n_115), .Y(n_139) );
INVx2_ASAP7_75t_L g226 ( .A(n_115), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_117), .B(n_141), .Y(n_140) );
INVxp67_ASAP7_75t_L g211 ( .A(n_117), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_117), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
INVx2_ASAP7_75t_SL g125 ( .A(n_119), .Y(n_125) );
CKINVDCx6p67_ASAP7_75t_R g198 ( .A(n_119), .Y(n_198) );
INVx2_ASAP7_75t_SL g213 ( .A(n_119), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_124), .B(n_125), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g144 ( .A1(n_122), .A2(n_145), .B1(n_147), .B2(n_148), .Y(n_144) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_122), .A2(n_157), .B1(n_207), .B2(n_208), .Y(n_206) );
INVx5_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g248 ( .A(n_123), .B(n_249), .Y(n_248) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_129), .B(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_129), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_152), .Y(n_130) );
INVx1_ASAP7_75t_L g275 ( .A(n_131), .Y(n_275) );
INVxp67_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g370 ( .A(n_132), .B(n_259), .Y(n_370) );
AND2x2_ASAP7_75t_L g384 ( .A(n_132), .B(n_153), .Y(n_384) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g261 ( .A(n_133), .B(n_153), .Y(n_261) );
AND2x2_ASAP7_75t_L g357 ( .A(n_133), .B(n_153), .Y(n_357) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g282 ( .A(n_134), .Y(n_282) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_143), .B(n_151), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_140), .B(n_142), .Y(n_135) );
NOR2x1_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_139), .A2(n_241), .B1(n_242), .B2(n_244), .Y(n_240) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g704 ( .A(n_147), .Y(n_704) );
AND2x2_ASAP7_75t_L g274 ( .A(n_152), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g314 ( .A(n_152), .Y(n_314) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_172), .Y(n_152) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_153), .Y(n_264) );
INVx2_ASAP7_75t_SL g299 ( .A(n_153), .Y(n_299) );
INVx1_ASAP7_75t_L g308 ( .A(n_153), .Y(n_308) );
AND2x2_ASAP7_75t_L g469 ( .A(n_153), .B(n_325), .Y(n_469) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_164), .B(n_169), .Y(n_153) );
OAI21xp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_162), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_155), .A2(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_L g231 ( .A(n_155), .Y(n_231) );
OAI22xp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B1(n_160), .B2(n_161), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g167 ( .A(n_158), .Y(n_167) );
INVx2_ASAP7_75t_L g196 ( .A(n_158), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_160), .A2(n_166), .B1(n_167), .B2(n_168), .Y(n_165) );
INVx2_ASAP7_75t_L g174 ( .A(n_170), .Y(n_174) );
NOR2x1p5_ASAP7_75t_SL g214 ( .A(n_170), .B(n_215), .Y(n_214) );
BUFx5_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g186 ( .A(n_171), .Y(n_186) );
INVx1_ASAP7_75t_L g342 ( .A(n_172), .Y(n_342) );
INVx2_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g259 ( .A(n_173), .Y(n_259) );
AND2x2_ASAP7_75t_L g307 ( .A(n_173), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g324 ( .A(n_173), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g397 ( .A(n_173), .Y(n_397) );
AO31x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .A3(n_183), .B(n_184), .Y(n_173) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g193 ( .A1(n_183), .A2(n_194), .B(n_199), .Y(n_193) );
OAI21x1_ASAP7_75t_SL g222 ( .A1(n_183), .A2(n_223), .B(n_228), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_216), .Y(n_187) );
OR2x2_ASAP7_75t_L g475 ( .A(n_188), .B(n_436), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_203), .Y(n_188) );
INVx2_ASAP7_75t_L g234 ( .A(n_189), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_189), .B(n_220), .Y(n_305) );
AND2x2_ASAP7_75t_L g329 ( .A(n_189), .B(n_272), .Y(n_329) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g270 ( .A(n_190), .Y(n_270) );
OAI21x1_ASAP7_75t_SL g190 ( .A1(n_191), .A2(n_193), .B(n_202), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_197), .B(n_198), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_198), .A2(n_206), .B(n_209), .C(n_214), .Y(n_205) );
INVx1_ASAP7_75t_L g219 ( .A(n_203), .Y(n_219) );
INVx1_ASAP7_75t_L g236 ( .A(n_203), .Y(n_236) );
INVx2_ASAP7_75t_L g294 ( .A(n_203), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_203), .B(n_237), .Y(n_303) );
AND2x2_ASAP7_75t_L g335 ( .A(n_203), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g347 ( .A(n_203), .B(n_220), .Y(n_347) );
INVx1_ASAP7_75t_L g425 ( .A(n_203), .Y(n_425) );
AND2x4_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_212), .C(n_213), .Y(n_209) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g277 ( .A(n_218), .Y(n_277) );
AND2x2_ASAP7_75t_L g371 ( .A(n_218), .B(n_285), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_218), .B(n_352), .Y(n_373) );
AND2x4_ASAP7_75t_L g432 ( .A(n_218), .B(n_387), .Y(n_432) );
AND2x4_ASAP7_75t_L g447 ( .A(n_218), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
INVx1_ASAP7_75t_L g419 ( .A(n_220), .Y(n_419) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
BUFx3_ASAP7_75t_L g272 ( .A(n_221), .Y(n_272) );
AOI21x1_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_227), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .Y(n_228) );
AND2x4_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
AND2x2_ASAP7_75t_L g364 ( .A(n_234), .B(n_302), .Y(n_364) );
INVx1_ASAP7_75t_L g399 ( .A(n_234), .Y(n_399) );
INVx2_ASAP7_75t_L g448 ( .A(n_234), .Y(n_448) );
AND2x2_ASAP7_75t_L g466 ( .A(n_234), .B(n_347), .Y(n_466) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_235), .Y(n_350) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx1_ASAP7_75t_L g362 ( .A(n_237), .Y(n_362) );
AND2x2_ASAP7_75t_L g390 ( .A(n_237), .B(n_272), .Y(n_390) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
BUFx3_ASAP7_75t_L g287 ( .A(n_238), .Y(n_287) );
INVx1_ASAP7_75t_L g337 ( .A(n_238), .Y(n_337) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_247), .B(n_253), .Y(n_238) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVxp67_ASAP7_75t_L g254 ( .A(n_245), .Y(n_254) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_262), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
AND2x4_ASAP7_75t_SL g365 ( .A(n_258), .B(n_298), .Y(n_365) );
AND2x4_ASAP7_75t_L g415 ( .A(n_260), .B(n_266), .Y(n_415) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g401 ( .A(n_261), .B(n_285), .Y(n_401) );
INVx1_ASAP7_75t_L g405 ( .A(n_261), .Y(n_405) );
OAI222xp33_ASAP7_75t_L g470 ( .A1(n_262), .A2(n_471), .B1(n_473), .B2(n_475), .C1(n_476), .C2(n_478), .Y(n_470) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g322 ( .A(n_264), .Y(n_322) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_266), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g296 ( .A(n_266), .Y(n_296) );
AND2x2_ASAP7_75t_L g332 ( .A(n_266), .B(n_322), .Y(n_332) );
AND2x2_ASAP7_75t_L g383 ( .A(n_266), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g421 ( .A(n_266), .B(n_356), .Y(n_421) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_273), .B(n_276), .C(n_283), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx1_ASAP7_75t_L g311 ( .A(n_269), .Y(n_311) );
AND2x4_ASAP7_75t_L g320 ( .A(n_269), .B(n_272), .Y(n_320) );
BUFx2_ASAP7_75t_L g387 ( .A(n_269), .Y(n_387) );
AND2x2_ASAP7_75t_L g412 ( .A(n_269), .B(n_294), .Y(n_412) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g352 ( .A(n_270), .B(n_287), .Y(n_352) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g293 ( .A(n_272), .B(n_294), .Y(n_293) );
BUFx2_ASAP7_75t_L g411 ( .A(n_272), .Y(n_411) );
INVx2_ASAP7_75t_SL g439 ( .A(n_274), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_280), .B(n_324), .Y(n_450) );
AND2x2_ASAP7_75t_L g459 ( .A(n_280), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g341 ( .A(n_281), .B(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_281), .B(n_342), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_281), .B(n_325), .Y(n_456) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g298 ( .A(n_282), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g464 ( .A(n_282), .B(n_325), .Y(n_464) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g292 ( .A(n_285), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g377 ( .A(n_285), .B(n_363), .Y(n_377) );
AND2x2_ASAP7_75t_L g431 ( .A(n_285), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g438 ( .A(n_285), .B(n_320), .Y(n_438) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_315), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI221xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_295), .B1(n_300), .B2(n_306), .C(n_309), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g310 ( .A(n_293), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g452 ( .A(n_293), .Y(n_452) );
INVx1_ASAP7_75t_L g388 ( .A(n_294), .Y(n_388) );
OR2x6_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_297), .A2(n_349), .B1(n_351), .B2(n_353), .Y(n_348) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g343 ( .A(n_298), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g369 ( .A(n_299), .B(n_325), .Y(n_369) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_302), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g318 ( .A(n_303), .Y(n_318) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g463 ( .A(n_307), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g460 ( .A(n_308), .B(n_397), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_311), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_313), .A2(n_331), .B(n_333), .Y(n_330) );
OR2x2_ASAP7_75t_L g374 ( .A(n_314), .B(n_375), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_330), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_321), .B1(n_326), .B2(n_328), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g334 ( .A(n_320), .B(n_335), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_320), .A2(n_327), .B1(n_368), .B2(n_371), .C(n_372), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_320), .B(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g406 ( .A(n_324), .B(n_357), .Y(n_406) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_325), .Y(n_355) );
INVx1_ASAP7_75t_L g376 ( .A(n_325), .Y(n_376) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_329), .B(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_L g422 ( .A(n_329), .Y(n_422) );
AND2x2_ASAP7_75t_L g435 ( .A(n_329), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVxp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g382 ( .A(n_335), .Y(n_382) );
INVx2_ASAP7_75t_L g436 ( .A(n_336), .Y(n_436) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_337), .Y(n_409) );
NOR2x1_ASAP7_75t_L g338 ( .A(n_339), .B(n_366), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_340), .B(n_358), .Y(n_339) );
O2A1O1Ixp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B(n_345), .C(n_348), .Y(n_340) );
AND2x2_ASAP7_75t_L g427 ( .A(n_344), .B(n_384), .Y(n_427) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_344), .Y(n_444) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g363 ( .A(n_347), .Y(n_363) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g430 ( .A(n_356), .Y(n_430) );
BUFx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_357), .B(n_375), .Y(n_378) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_364), .B(n_365), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_359), .A2(n_403), .B1(n_406), .B2(n_407), .Y(n_402) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g467 ( .A(n_361), .Y(n_467) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_362), .B(n_419), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_379), .Y(n_366) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_369), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_SL g468 ( .A(n_370), .B(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g472 ( .A(n_370), .B(n_375), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_370), .B(n_469), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B1(n_377), .B2(n_378), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OA22x2_ASAP7_75t_L g449 ( .A1(n_377), .A2(n_450), .B1(n_451), .B2(n_454), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B(n_385), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
AOI21xp33_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_389), .B(n_391), .Y(n_385) );
NAND2xp33_ASAP7_75t_SL g416 ( .A(n_386), .B(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2x1_ASAP7_75t_L g393 ( .A(n_394), .B(n_413), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_398), .B(n_402), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g455 ( .A(n_396), .Y(n_455) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OA21x2_ASAP7_75t_L g442 ( .A1(n_401), .A2(n_443), .B(n_445), .Y(n_442) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
AND2x2_ASAP7_75t_L g429 ( .A(n_404), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g445 ( .A(n_406), .Y(n_445) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g420 ( .A(n_408), .Y(n_420) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g461 ( .A(n_410), .Y(n_461) );
AND2x4_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_428), .Y(n_413) );
AOI222xp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_421), .B2(n_422), .C1(n_423), .C2(n_427), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g457 ( .A1(n_424), .A2(n_458), .B1(n_461), .B2(n_462), .C(n_465), .Y(n_457) );
OR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_426), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B(n_433), .Y(n_428) );
AOI21xp5_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_437), .B(n_439), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g453 ( .A(n_436), .Y(n_453) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR3x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_457), .C(n_470), .Y(n_440) );
OAI21x1_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_446), .B(n_449), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x6_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g477 ( .A(n_452), .Y(n_477) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_468), .Y(n_465) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI221xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_658), .B2(n_663), .C(n_700), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_481), .A2(n_701), .B1(n_704), .B2(n_705), .Y(n_700) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND4xp75_ASAP7_75t_L g483 ( .A(n_484), .B(n_556), .C(n_636), .D(n_649), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_532), .Y(n_484) );
AOI33xp33_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_494), .A3(n_507), .B1(n_517), .B2(n_524), .B3(n_528), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_492), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g687 ( .A(n_489), .Y(n_687) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AND2x4_ASAP7_75t_L g530 ( .A(n_490), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_491), .Y(n_531) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g635 ( .A(n_493), .Y(n_635) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g525 ( .A(n_496), .Y(n_525) );
INVx2_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g657 ( .A(n_498), .Y(n_657) );
INVx2_ASAP7_75t_L g512 ( .A(n_499), .Y(n_512) );
AND2x2_ASAP7_75t_L g516 ( .A(n_499), .B(n_505), .Y(n_516) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_504), .Y(n_527) );
INVx1_ASAP7_75t_L g646 ( .A(n_504), .Y(n_646) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx2_ASAP7_75t_L g513 ( .A(n_505), .Y(n_513) );
INVx1_ASAP7_75t_L g656 ( .A(n_506), .Y(n_656) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_SL g520 ( .A(n_510), .Y(n_520) );
INVx6_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g639 ( .A(n_511), .Y(n_639) );
AND2x2_ASAP7_75t_L g648 ( .A(n_511), .B(n_540), .Y(n_648) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g550 ( .A(n_512), .Y(n_550) );
INVx1_ASAP7_75t_L g537 ( .A(n_513), .Y(n_537) );
BUFx4f_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_516), .Y(n_523) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g554 ( .A(n_523), .Y(n_554) );
AND2x2_ASAP7_75t_L g650 ( .A(n_525), .B(n_640), .Y(n_650) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
AND2x4_ASAP7_75t_L g647 ( .A(n_529), .B(n_648), .Y(n_647) );
AND2x4_ASAP7_75t_L g540 ( .A(n_531), .B(n_541), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_545), .B1(n_546), .B2(n_551), .C(n_552), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
INVx1_ASAP7_75t_L g689 ( .A(n_535), .Y(n_689) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g695 ( .A(n_536), .Y(n_695) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
OR2x6_ASAP7_75t_L g547 ( .A(n_539), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g555 ( .A(n_539), .Y(n_555) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .Y(n_539) );
AND2x4_ASAP7_75t_L g694 ( .A(n_540), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g641 ( .A(n_544), .B(n_642), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_545), .A2(n_551), .B1(n_624), .B2(n_627), .Y(n_623) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_593), .B(n_633), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_577), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B1(n_569), .B2(n_570), .Y(n_558) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
INVx2_ASAP7_75t_L g572 ( .A(n_561), .Y(n_572) );
AND2x4_ASAP7_75t_L g592 ( .A(n_561), .B(n_583), .Y(n_592) );
INVx1_ASAP7_75t_L g590 ( .A(n_562), .Y(n_590) );
INVx1_ASAP7_75t_L g600 ( .A(n_562), .Y(n_600) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_563), .Y(n_579) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_564), .B(n_568), .Y(n_610) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x4_ASAP7_75t_L g575 ( .A(n_565), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g584 ( .A(n_565), .B(n_568), .Y(n_584) );
INVx1_ASAP7_75t_L g587 ( .A(n_565), .Y(n_587) );
INVx1_ASAP7_75t_L g622 ( .A(n_565), .Y(n_622) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g576 ( .A(n_568), .Y(n_576) );
INVx1_ASAP7_75t_L g621 ( .A(n_568), .Y(n_621) );
INVx1_ASAP7_75t_L g626 ( .A(n_568), .Y(n_626) );
AND2x4_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
AND2x4_ASAP7_75t_L g612 ( .A(n_571), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_575), .Y(n_580) );
INVx3_ASAP7_75t_L g606 ( .A(n_575), .Y(n_606) );
AND2x4_ASAP7_75t_L g586 ( .A(n_576), .B(n_587), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B1(n_591), .B2(n_592), .Y(n_577) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g617 ( .A(n_583), .Y(n_617) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx3_ASAP7_75t_L g596 ( .A(n_584), .Y(n_596) );
BUFx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_586), .Y(n_597) );
BUFx3_ASAP7_75t_L g613 ( .A(n_586), .Y(n_613) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2x1p5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B1(n_607), .B2(n_608), .Y(n_602) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_603), .A2(n_615), .B1(n_637), .B2(n_643), .C1(n_644), .C2(n_647), .Y(n_636) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_607), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_649) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx8_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .B(n_618), .C(n_629), .Y(n_614) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_623), .Y(n_618) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g628 ( .A(n_622), .Y(n_628) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx8_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x6_ASAP7_75t_L g645 ( .A(n_641), .B(n_646), .Y(n_645) );
OR2x6_ASAP7_75t_L g653 ( .A(n_641), .B(n_654), .Y(n_653) );
CKINVDCx6p67_ASAP7_75t_R g644 ( .A(n_645), .Y(n_644) );
CKINVDCx6p67_ASAP7_75t_R g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
BUFx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_660), .B(n_662), .Y(n_683) );
INVx1_ASAP7_75t_SL g707 ( .A(n_660), .Y(n_707) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_679), .B1(n_696), .B2(n_697), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_664), .A2(n_696), .B1(n_702), .B2(n_703), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_673), .B2(n_674), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_669), .B2(n_672), .Y(n_666) );
CKINVDCx5p33_ASAP7_75t_R g672 ( .A(n_667), .Y(n_672) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
XOR2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_677), .B2(n_678), .Y(n_674) );
CKINVDCx5p33_ASAP7_75t_R g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx8_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx8_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
CKINVDCx20_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
BUFx4f_ASAP7_75t_L g702 ( .A(n_682), .Y(n_702) );
OR2x6_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
OR2x4_ASAP7_75t_L g699 ( .A(n_683), .B(n_685), .Y(n_699) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI31xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .A3(n_690), .B(n_692), .Y(n_685) );
BUFx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx6_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g703 ( .A(n_698), .Y(n_703) );
INVx8_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
BUFx2_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
endmodule