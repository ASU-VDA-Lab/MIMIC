module real_jpeg_33146_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_687, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_687;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_679;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_666;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_578;
wire n_328;
wire n_366;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_525;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_338;
wire n_175;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_650;
wire n_250;
wire n_254;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_586;
wire n_405;
wire n_412;
wire n_572;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_642;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_667;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_675;
wire n_179;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_268;
wire n_42;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_0),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_0),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_0),
.Y(n_379)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_0),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_1),
.A2(n_313),
.B1(n_314),
.B2(n_316),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_1),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_1),
.A2(n_313),
.B1(n_369),
.B2(n_371),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_1),
.A2(n_313),
.B1(n_511),
.B2(n_515),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_1),
.A2(n_313),
.B1(n_579),
.B2(n_581),
.Y(n_578)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_2),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

OAI22x1_ASAP7_75t_L g228 ( 
.A1(n_2),
.A2(n_95),
.B1(n_229),
.B2(n_232),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_2),
.A2(n_95),
.B1(n_287),
.B2(n_292),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_2),
.A2(n_95),
.B1(n_386),
.B2(n_390),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_3),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_4),
.A2(n_65),
.B1(n_67),
.B2(n_69),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_4),
.A2(n_69),
.B1(n_126),
.B2(n_130),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_4),
.A2(n_69),
.B1(n_148),
.B2(n_152),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_4),
.A2(n_69),
.B1(n_250),
.B2(n_253),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_5),
.A2(n_97),
.B1(n_338),
.B2(n_341),
.Y(n_337)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_5),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_5),
.A2(n_341),
.B1(n_420),
.B2(n_422),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_5),
.A2(n_341),
.B1(n_571),
.B2(n_573),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_5),
.A2(n_341),
.B1(n_642),
.B2(n_645),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_6),
.A2(n_58),
.B1(n_83),
.B2(n_89),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_6),
.A2(n_89),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_6),
.A2(n_89),
.B1(n_256),
.B2(n_260),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_6),
.A2(n_89),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_7),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_8),
.Y(n_143)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_8),
.Y(n_160)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_9),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_10),
.A2(n_361),
.B1(n_364),
.B2(n_367),
.Y(n_360)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_10),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_10),
.A2(n_334),
.B1(n_338),
.B2(n_367),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_10),
.A2(n_367),
.B1(n_551),
.B2(n_554),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_10),
.A2(n_367),
.B1(n_630),
.B2(n_633),
.Y(n_629)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_11),
.Y(n_105)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_11),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_12),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_L g263 ( 
.A1(n_13),
.A2(n_264),
.B1(n_268),
.B2(n_269),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_13),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_13),
.A2(n_268),
.B1(n_352),
.B2(n_355),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_13),
.A2(n_268),
.B1(n_452),
.B2(n_457),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_13),
.A2(n_268),
.B1(n_305),
.B2(n_535),
.Y(n_534)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_14),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_14),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_14),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_14),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_15),
.A2(n_191),
.B1(n_192),
.B2(n_194),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_15),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_15),
.A2(n_191),
.B1(n_321),
.B2(n_324),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_15),
.A2(n_191),
.B1(n_428),
.B2(n_430),
.Y(n_427)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_16),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_16),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_21),
.B(n_24),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_18),
.A2(n_53),
.B1(n_57),
.B2(n_62),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_18),
.A2(n_62),
.B1(n_168),
.B2(n_171),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_18),
.A2(n_62),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_18),
.A2(n_62),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_19),
.A2(n_333),
.B(n_336),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_19),
.B(n_335),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_19),
.Y(n_440)
);

OAI32xp33_ASAP7_75t_L g519 ( 
.A1(n_19),
.A2(n_163),
.A3(n_520),
.B1(n_521),
.B2(n_525),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_19),
.A2(n_440),
.B1(n_559),
.B2(n_560),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_19),
.B(n_139),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_19),
.A2(n_246),
.B1(n_641),
.B2(n_650),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_72),
.B(n_680),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_70),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_27),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_27),
.B(n_75),
.Y(n_679)
);

CKINVDCx16_ASAP7_75t_R g683 ( 
.A(n_27),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_28),
.A2(n_63),
.B(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_28),
.A2(n_52),
.B1(n_63),
.B2(n_82),
.Y(n_173)
);

OAI22x1_ASAP7_75t_L g310 ( 
.A1(n_28),
.A2(n_63),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_28),
.A2(n_63),
.B1(n_332),
.B2(n_337),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_28),
.A2(n_63),
.B1(n_312),
.B2(n_448),
.Y(n_472)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_29),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_29),
.A2(n_80),
.B1(n_190),
.B2(n_263),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_41),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_30)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_31),
.Y(n_325)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_32),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_33),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_33),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g424 ( 
.A(n_33),
.Y(n_424)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_34),
.Y(n_404)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_39),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_40),
.Y(n_164)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_40),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_40),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_47),
.B2(n_50),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_43),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_44),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_44),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_44),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_60),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_63),
.B(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_68),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_71),
.B(n_683),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_326),
.B(n_673),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_177),
.C(n_204),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_74),
.A2(n_674),
.B(n_679),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_173),
.C(n_174),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_76),
.A2(n_77),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_98),
.C(n_135),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_79),
.B(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_90),
.B2(n_91),
.Y(n_79)
);

AO22x1_ASAP7_75t_L g188 ( 
.A1(n_80),
.A2(n_91),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

AOI22x1_ASAP7_75t_L g446 ( 
.A1(n_80),
.A2(n_189),
.B1(n_447),
.B2(n_449),
.Y(n_446)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_86),
.Y(n_193)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_99),
.B(n_187),
.C(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_100),
.A2(n_136),
.B1(n_137),
.B2(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_100),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_100),
.A2(n_186),
.B1(n_199),
.B2(n_211),
.Y(n_210)
);

AO21x2_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_124),
.B(n_125),
.Y(n_100)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_101),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_101),
.A2(n_124),
.B1(n_219),
.B2(n_255),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_101),
.A2(n_124),
.B1(n_255),
.B2(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_101),
.A2(n_124),
.B1(n_344),
.B2(n_351),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_101),
.A2(n_124),
.B1(n_286),
.B2(n_344),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_101),
.A2(n_124),
.B1(n_351),
.B2(n_509),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_101),
.A2(n_124),
.B1(n_550),
.B2(n_569),
.Y(n_568)
);

AO21x2_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_110),
.B(n_115),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_108),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_109),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_110),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_112),
.Y(n_347)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_112),
.Y(n_516)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

OAI22x1_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_118),
.B1(n_121),
.B2(n_123),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_118),
.Y(n_253)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_120),
.Y(n_252)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_120),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_120),
.Y(n_609)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_121),
.Y(n_247)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_121),
.Y(n_304)
);

BUFx2_ASAP7_75t_SL g660 ( 
.A(n_121),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_122),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_122),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_124),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_124),
.B(n_440),
.Y(n_647)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_125),
.Y(n_216)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_128),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_129),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_129),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_133),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_134),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_134),
.Y(n_354)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_134),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_134),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_147),
.B1(n_156),
.B2(n_167),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_138),
.A2(n_156),
.B1(n_167),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_138),
.A2(n_156),
.B1(n_360),
.B2(n_368),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_138),
.A2(n_156),
.B1(n_360),
.B2(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_138),
.A2(n_156),
.B1(n_368),
.B2(n_451),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_138),
.A2(n_156),
.B1(n_320),
.B2(n_451),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_138),
.A2(n_156),
.B1(n_419),
.B2(n_558),
.Y(n_557)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_139),
.A2(n_175),
.B1(n_201),
.B2(n_228),
.Y(n_227)
);

AOI22x1_ASAP7_75t_L g318 ( 
.A1(n_139),
.A2(n_175),
.B1(n_228),
.B2(n_319),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AO21x2_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_157),
.B(n_163),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_145),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_150),
.Y(n_363)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_150),
.Y(n_370)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_151),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_151),
.Y(n_421)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_152),
.Y(n_520)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

NAND2xp33_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_164),
.Y(n_559)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_174),
.Y(n_181)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g674 ( 
.A1(n_178),
.A2(n_675),
.B(n_678),
.Y(n_674)
);

NOR2x1_ASAP7_75t_R g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_179),
.B(n_182),
.Y(n_678)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.C(n_197),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_184),
.B(n_187),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_191),
.A2(n_345),
.B(n_348),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_191),
.B(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_197),
.B(n_271),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_272),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_206),
.A2(n_676),
.B(n_677),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_270),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_207),
.B(n_270),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.C(n_237),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_209),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_213),
.B(n_275),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_213),
.A2(n_214),
.B(n_227),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_227),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_215),
.A2(n_217),
.B1(n_510),
.B2(n_549),
.Y(n_548)
);

AOI22x1_ASAP7_75t_SL g594 ( 
.A1(n_215),
.A2(n_217),
.B1(n_570),
.B2(n_595),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_225),
.Y(n_603)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_226),
.Y(n_599)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx5_ASAP7_75t_L g560 ( 
.A(n_230),
.Y(n_560)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_240),
.B1(n_261),
.B2(n_687),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_279),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_254),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_262),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_240),
.B(n_254),
.Y(n_482)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_245),
.B(n_248),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_241),
.A2(n_384),
.B1(n_628),
.B2(n_636),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_243),
.A2(n_246),
.B1(n_303),
.B2(n_381),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g640 ( 
.A1(n_243),
.A2(n_246),
.B1(n_629),
.B2(n_641),
.Y(n_640)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_243),
.Y(n_657)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_247),
.Y(n_246)
);

INVx8_ASAP7_75t_L g436 ( 
.A(n_244),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_245),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_246),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_246),
.A2(n_578),
.B1(n_585),
.B2(n_586),
.Y(n_577)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_249),
.A2(n_296),
.B(n_301),
.Y(n_295)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_251),
.Y(n_382)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_252),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_259),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_265),
.Y(n_335)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_273),
.B(n_276),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.C(n_282),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_278),
.A2(n_280),
.B1(n_281),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_278),
.Y(n_494)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_283),
.B(n_493),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_309),
.C(n_317),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_284),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_295),
.Y(n_284)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_285),
.Y(n_478)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_294),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_295),
.B(n_478),
.Y(n_477)
);

INVx3_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_300),
.Y(n_585)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_307),
.Y(n_429)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_307),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx6_ASAP7_75t_L g389 ( 
.A(n_308),
.Y(n_389)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_308),
.Y(n_620)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_308),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_309),
.A2(n_310),
.B1(n_318),
.B2(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_318),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_323),
.Y(n_372)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_323),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

OA21x2_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_502),
.B(n_667),
.Y(n_326)
);

NAND4xp25_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_465),
.C(n_489),
.D(n_495),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_442),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_329),
.B(n_442),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_373),
.B(n_441),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_330),
.B(n_540),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_342),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g464 ( 
.A(n_331),
.B(n_343),
.C(n_359),
.Y(n_464)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_SL g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_337),
.Y(n_449)
);

INVx11_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx12f_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_359),
.Y(n_342)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_366),
.Y(n_458)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_371),
.Y(n_398)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_416),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_374),
.B(n_416),
.Y(n_441)
);

OA21x2_ASAP7_75t_SL g374 ( 
.A1(n_375),
.A2(n_394),
.B(n_415),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_376),
.A2(n_377),
.B1(n_394),
.B2(n_395),
.Y(n_541)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_396),
.Y(n_415)
);

AO22x1_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_380),
.B1(n_384),
.B2(n_385),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_384),
.A2(n_385),
.B1(n_427),
.B2(n_434),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_384),
.A2(n_427),
.B1(n_530),
.B2(n_534),
.Y(n_529)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_389),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_389),
.Y(n_635)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_389),
.Y(n_644)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx2_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

OAI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_397),
.A2(n_399),
.B1(n_405),
.B2(n_414),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_403),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_410),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

BUFx2_ASAP7_75t_SL g411 ( 
.A(n_412),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XOR2x2_ASAP7_75t_SL g443 ( 
.A(n_415),
.B(n_444),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_415),
.B(n_446),
.C(n_459),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_416),
.A2(n_417),
.B1(n_541),
.B2(n_542),
.Y(n_540)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_425),
.C(n_437),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_418),
.B(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_421),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_424),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_425),
.A2(n_426),
.B1(n_438),
.B2(n_439),
.Y(n_507)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_435),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_440),
.B(n_526),
.Y(n_525)
);

OAI21xp33_ASAP7_75t_SL g595 ( 
.A1(n_440),
.A2(n_596),
.B(n_600),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_440),
.B(n_601),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_440),
.B(n_656),
.Y(n_655)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_460),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_443),
.B(n_461),
.C(n_497),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_450),
.B2(n_459),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_450),
.Y(n_459)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_464),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_463),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_464),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_480),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_SL g668 ( 
.A(n_466),
.B(n_480),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_SL g671 ( 
.A1(n_466),
.A2(n_480),
.B1(n_490),
.B2(n_492),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_476),
.C(n_479),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_468),
.B(n_501),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_471),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_487),
.C(n_488),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_473),
.B1(n_474),
.B2(n_475),
.Y(n_471)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_472),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_473),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_474),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_475),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_477),
.Y(n_501)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_479),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_486),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_482),
.B(n_486),
.C(n_491),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_483),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_492),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_490),
.B(n_492),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_498),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_496),
.B(n_498),
.C(n_670),
.Y(n_669)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

AOI21x1_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_543),
.B(n_666),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_539),
.Y(n_503)
);

NOR2xp67_ASAP7_75t_SL g666 ( 
.A(n_504),
.B(n_539),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_508),
.C(n_517),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_505),
.A2(n_506),
.B1(n_562),
.B2(n_563),
.Y(n_561)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_508),
.A2(n_517),
.B1(n_518),
.B2(n_564),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_508),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_528),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_519),
.A2(n_528),
.B1(n_529),
.B2(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_519),
.Y(n_547)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_524),
.Y(n_555)
);

INVx4_ASAP7_75t_SL g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_533),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_534),
.Y(n_586)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_541),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_544),
.A2(n_565),
.B(n_665),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_561),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_545),
.B(n_561),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_548),
.C(n_556),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_546),
.B(n_588),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_548),
.A2(n_556),
.B1(n_557),
.B2(n_589),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_548),
.Y(n_589)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_552),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

AOI21x1_ASAP7_75t_L g565 ( 
.A1(n_566),
.A2(n_590),
.B(n_664),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_567),
.B(n_587),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_567),
.B(n_587),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_575),
.C(n_577),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_568),
.A2(n_575),
.B1(n_576),
.B2(n_624),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_568),
.Y(n_624)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_572),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_577),
.B(n_623),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_578),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_591),
.A2(n_625),
.B(n_663),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_592),
.B(n_622),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_592),
.B(n_622),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_593),
.B(n_604),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_593),
.A2(n_594),
.B1(n_604),
.B2(n_605),
.Y(n_637)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx5_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_600),
.Y(n_615)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_606),
.A2(n_615),
.B1(n_616),
.B2(n_621),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_607),
.B(n_610),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx6_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_626),
.A2(n_638),
.B(n_662),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_627),
.B(n_637),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g662 ( 
.A(n_627),
.B(n_637),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_634),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_SL g638 ( 
.A1(n_639),
.A2(n_648),
.B(n_661),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_640),
.B(n_647),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_640),
.B(n_647),
.Y(n_661)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_643),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_646),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_649),
.B(n_654),
.Y(n_648)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_651),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_652),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_653),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_655),
.B(n_658),
.Y(n_654)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_657),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_659),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_660),
.Y(n_659)
);

O2A1O1Ixp5_ASAP7_75t_L g667 ( 
.A1(n_668),
.A2(n_669),
.B(n_671),
.C(n_672),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_681),
.B(n_684),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_682),
.Y(n_681)
);

CKINVDCx11_ASAP7_75t_R g684 ( 
.A(n_685),
.Y(n_684)
);


endmodule