module fake_jpeg_5435_n_73 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_73);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_73;

wire n_61;
wire n_45;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_59;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_38;
wire n_56;
wire n_50;
wire n_67;
wire n_57;
wire n_53;
wire n_54;
wire n_69;
wire n_40;
wire n_71;
wire n_48;
wire n_35;
wire n_46;
wire n_44;
wire n_36;
wire n_62;
wire n_37;
wire n_43;
wire n_70;
wire n_66;

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_17),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_49),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_0),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_52),
.Y(n_57)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_43),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_1),
.B(n_7),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_34),
.B1(n_2),
.B2(n_4),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_9),
.B1(n_11),
.B2(n_16),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_SL g58 ( 
.A(n_51),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_32),
.B1(n_5),
.B2(n_6),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_62),
.B1(n_54),
.B2(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_59),
.B1(n_23),
.B2(n_24),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_66),
.C(n_25),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_68),
.A2(n_18),
.B(n_26),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_27),
.C(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_29),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);


endmodule