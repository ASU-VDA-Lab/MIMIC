module real_jpeg_10371_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_184;
wire n_48;
wire n_56;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_213;
wire n_167;
wire n_216;
wire n_179;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_41),
.B1(n_57),
.B2(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_41),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_47),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_4),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_4),
.A2(n_54),
.B(n_58),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_4),
.A2(n_52),
.B1(n_60),
.B2(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_4),
.B(n_64),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_4),
.A2(n_38),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_38),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_4),
.A2(n_81),
.B1(n_82),
.B2(n_200),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_7),
.A2(n_38),
.B(n_43),
.C(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_38),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_7),
.A2(n_27),
.B1(n_30),
.B2(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_SL g69 ( 
.A(n_8),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_10),
.A2(n_35),
.B1(n_52),
.B2(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_35),
.B1(n_57),
.B2(n_58),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_10),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_11),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_11),
.A2(n_29),
.B1(n_57),
.B2(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_11),
.A2(n_29),
.B1(n_38),
.B2(n_39),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_13),
.A2(n_52),
.B1(n_60),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_13),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_120),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_120),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_13),
.A2(n_27),
.B1(n_30),
.B2(n_120),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_52),
.B1(n_60),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_14),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_101),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_14),
.A2(n_27),
.B1(n_30),
.B2(n_101),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_101),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_15),
.A2(n_52),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_15),
.A2(n_27),
.B1(n_30),
.B2(n_61),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_61),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_130),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_19),
.B(n_105),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_89),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_77),
.B2(n_78),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_24),
.B(n_36),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_25),
.A2(n_82),
.B(n_127),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_26),
.B(n_32),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_27),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_191)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_30),
.B(n_45),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_30),
.B(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_31),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_31),
.A2(n_32),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_32),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_33),
.A2(n_81),
.B(n_184),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_34),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_37),
.A2(n_44),
.B(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_39),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_38),
.B(n_68),
.Y(n_228)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_39),
.A2(n_73),
.B1(n_223),
.B2(n_228),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_42),
.A2(n_46),
.B(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_42),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_42),
.A2(n_44),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_42),
.A2(n_44),
.B1(n_190),
.B2(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_42),
.A2(n_44),
.B1(n_213),
.B2(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_42),
.A2(n_221),
.B(n_244),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_43),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_44),
.B(n_124),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_44),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_65),
.B2(n_76),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_59),
.B(n_62),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_51),
.A2(n_56),
.B1(n_59),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_51),
.A2(n_56),
.B1(n_100),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_51),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B(n_55),
.C(n_56),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_52),
.A2(n_53),
.B(n_124),
.C(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_67),
.B(n_68),
.C(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_68),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g223 ( 
.A(n_58),
.B(n_124),
.CON(n_223),
.SN(n_223)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_64),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B(n_71),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_75),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_66),
.A2(n_114),
.B1(n_115),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_66),
.A2(n_114),
.B1(n_144),
.B2(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_66),
.B(n_124),
.Y(n_211)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_103),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_67),
.A2(n_72),
.B1(n_168),
.B2(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_72),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_88),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_83),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_81),
.A2(n_82),
.B1(n_92),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_81),
.A2(n_82),
.B1(n_182),
.B2(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_81),
.A2(n_83),
.B(n_93),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_82),
.B(n_124),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_86),
.A2(n_97),
.B(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.C(n_102),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.C(n_110),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_109),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_110),
.A2(n_111),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.C(n_121),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B(n_116),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_173),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_154),
.B(n_172),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_174),
.C(n_255),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_151),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_151),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.C(n_140),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_149),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_143),
.B1(n_149),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_150),
.B(n_245),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_152),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_155),
.B(n_157),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_163),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_158),
.B(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_161),
.A2(n_163),
.B1(n_164),
.B2(n_253),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_161),
.Y(n_253)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.C(n_170),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_165),
.A2(n_166),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_169),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_249),
.B(n_254),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_232),
.B(n_248),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_216),
.B(n_231),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_207),
.B(n_215),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_196),
.B(n_206),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_185),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_185),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_191),
.B2(n_195),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_195),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_189),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_201),
.B(n_205),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_198),
.B(n_199),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_208),
.B(n_209),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_210),
.B(n_217),
.Y(n_231)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.CI(n_214),
.CON(n_210),
.SN(n_210)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_226),
.B2(n_230),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_220),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_222),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_225),
.C(n_230),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_226),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_229),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_233),
.B(n_234),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_240),
.B2(n_241),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_243),
.C(n_246),
.Y(n_250)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_246),
.B2(n_247),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_242),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_243),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_250),
.B(n_251),
.Y(n_254)
);


endmodule