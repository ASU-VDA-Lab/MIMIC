module fake_jpeg_12345_n_20 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_20);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_20;

wire n_13;
wire n_10;
wire n_14;
wire n_19;
wire n_18;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx5_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_SL g12 ( 
.A1(n_10),
.A2(n_11),
.B(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

NAND3xp33_ASAP7_75t_L g14 ( 
.A(n_12),
.B(n_10),
.C(n_1),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_11),
.A2(n_9),
.B1(n_8),
.B2(n_0),
.Y(n_13)
);

A2O1A1O1Ixp25_ASAP7_75t_L g15 ( 
.A1(n_13),
.A2(n_0),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_14),
.A2(n_15),
.B1(n_1),
.B2(n_3),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_0),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_17),
.B(n_5),
.Y(n_18)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_18),
.B(n_16),
.CI(n_5),
.CON(n_19),
.SN(n_19)
);

AOI32xp33_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_6),
.A3(n_16),
.B1(n_14),
.B2(n_18),
.Y(n_20)
);


endmodule