module fake_netlist_5_2211_n_1855 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1855);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1855;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1699;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_48),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_21),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_136),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_99),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_53),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_107),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_60),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_169),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_80),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_82),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_101),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_77),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_27),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_76),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_94),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_168),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_43),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_122),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_91),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_23),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_139),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_93),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_7),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_152),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_57),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_0),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_25),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_28),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_7),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_132),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_113),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_52),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_14),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_38),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_48),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_64),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_121),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_34),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_165),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_154),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_137),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_92),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_36),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_45),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_51),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_103),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_71),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_140),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_151),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_0),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_105),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_109),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_108),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_161),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_42),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_174),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_142),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_42),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_51),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_86),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_134),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_155),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_78),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_124),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_27),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_29),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_100),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_102),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_14),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_176),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_33),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_13),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_13),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_10),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_123),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_17),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_58),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_79),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_62),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_47),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_158),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_66),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_114),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_1),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_37),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_37),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_67),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_90),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_34),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_4),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_81),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_112),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_73),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_128),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_24),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_18),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_172),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_49),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_150),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_175),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_162),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_117),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_3),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_75),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_173),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_146),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_49),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_26),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_126),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_141),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_8),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_145),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_171),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_22),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_69),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_50),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_9),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_104),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_4),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_157),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_44),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_35),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_96),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_56),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_18),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_12),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_17),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_22),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_72),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_21),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_147),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_15),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_44),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_68),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_19),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_85),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_19),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_35),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_59),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_23),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_8),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_52),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_144),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_160),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_163),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_148),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_65),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_127),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_70),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_83),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_63),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_54),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_115),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_43),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_143),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_149),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_55),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_32),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_41),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_97),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_36),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_31),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_120),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_41),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_12),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_88),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_116),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_38),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_5),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_61),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_30),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_6),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_187),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_318),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_283),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_R g357 ( 
.A(n_208),
.B(n_129),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_180),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_180),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_1),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_346),
.B(n_2),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_342),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_334),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_269),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_202),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_229),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_318),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_177),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_178),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_206),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_202),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_318),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_226),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_192),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_352),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_318),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_214),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_214),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_226),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_334),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_197),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_286),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_265),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_207),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_200),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_188),
.B(n_2),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_286),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_265),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_209),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_323),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_323),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_212),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_215),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_239),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_213),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_297),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_218),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_249),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_253),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_181),
.Y(n_401)
);

BUFx6f_ASAP7_75t_SL g402 ( 
.A(n_234),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_256),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_223),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_R g405 ( 
.A(n_326),
.B(n_170),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_260),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_326),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_230),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_194),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_224),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_329),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_329),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_335),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_270),
.Y(n_414)
);

INVxp33_ASAP7_75t_L g415 ( 
.A(n_278),
.Y(n_415)
);

INVxp33_ASAP7_75t_SL g416 ( 
.A(n_349),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_287),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_288),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_296),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_195),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_335),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_235),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_297),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_188),
.B(n_3),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_189),
.B(n_5),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_301),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_307),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_224),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_317),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_242),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_238),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_257),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_317),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_308),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_179),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_345),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_245),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_251),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_349),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_354),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_432),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_367),
.Y(n_444)
);

OA21x2_ASAP7_75t_L g445 ( 
.A1(n_432),
.A2(n_293),
.B(n_189),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_358),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_435),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_368),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_359),
.B(n_252),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_368),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_370),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_370),
.Y(n_454)
);

AND3x2_ASAP7_75t_L g455 ( 
.A(n_387),
.B(n_424),
.C(n_361),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_364),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_373),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_373),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_369),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_377),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_377),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_378),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_378),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_369),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_410),
.Y(n_467)
);

NOR2xp67_ASAP7_75t_L g468 ( 
.A(n_410),
.B(n_244),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_371),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_428),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_428),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_429),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_433),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_433),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_401),
.B(n_293),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_382),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_386),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_390),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_376),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_409),
.B(n_196),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_371),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_420),
.B(n_196),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_430),
.B(n_324),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_355),
.B(n_199),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_425),
.B(n_324),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_399),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_400),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_385),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_364),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_385),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_393),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_403),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_393),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_406),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_414),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_417),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_396),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_418),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_365),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_396),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_419),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_426),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_427),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_434),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_398),
.Y(n_509)
);

NAND2x1p5_ASAP7_75t_L g510 ( 
.A(n_360),
.B(n_261),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_436),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_437),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_372),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_356),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_398),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_363),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_381),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_455),
.B(n_353),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_478),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_441),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_488),
.B(n_405),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_443),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_488),
.A2(n_485),
.B1(n_476),
.B2(n_455),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_441),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_478),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_488),
.B(n_336),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_456),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_255),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_485),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_486),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_480),
.A2(n_366),
.B1(n_416),
.B2(n_440),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_486),
.Y(n_533)
);

OR2x6_ASAP7_75t_L g534 ( 
.A(n_487),
.B(n_203),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_489),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_514),
.B(n_284),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_441),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_476),
.B(n_375),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_488),
.B(n_476),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_450),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_482),
.B(n_416),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_442),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_481),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_487),
.B(n_203),
.Y(n_545)
);

BUFx4f_ASAP7_75t_L g546 ( 
.A(n_510),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_447),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_481),
.B(n_362),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_514),
.B(n_415),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_488),
.B(n_404),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_443),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_442),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_482),
.B(n_440),
.Y(n_553)
);

OAI22xp33_ASAP7_75t_L g554 ( 
.A1(n_480),
.A2(n_246),
.B1(n_225),
.B2(n_310),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_443),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_443),
.Y(n_556)
);

INVx6_ASAP7_75t_L g557 ( 
.A(n_443),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_489),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_443),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_490),
.Y(n_560)
);

INVxp67_ASAP7_75t_SL g561 ( 
.A(n_445),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_453),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_490),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_484),
.B(n_404),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_452),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_452),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_452),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_485),
.A2(n_510),
.B1(n_484),
.B2(n_445),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_495),
.B(n_336),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_454),
.Y(n_570)
);

AND3x2_ASAP7_75t_L g571 ( 
.A(n_456),
.B(n_423),
.C(n_397),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_485),
.B(n_261),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_450),
.A2(n_408),
.B1(n_431),
.B2(n_422),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_453),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_491),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_454),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_491),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_445),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_514),
.B(n_289),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_453),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_453),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_453),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_506),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_445),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_454),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_510),
.B(n_408),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_460),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_453),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_493),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_460),
.Y(n_590)
);

NOR2x1p5_ASAP7_75t_L g591 ( 
.A(n_448),
.B(n_422),
.Y(n_591)
);

INVxp67_ASAP7_75t_SL g592 ( 
.A(n_445),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_510),
.A2(n_439),
.B1(n_438),
.B2(n_431),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_453),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_460),
.Y(n_595)
);

INVx6_ASAP7_75t_L g596 ( 
.A(n_496),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_461),
.Y(n_597)
);

AO22x2_ASAP7_75t_L g598 ( 
.A1(n_449),
.A2(n_340),
.B1(n_331),
.B2(n_295),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_516),
.B(n_438),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_444),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_506),
.A2(n_357),
.B1(n_316),
.B2(n_261),
.Y(n_601)
);

INVx5_ASAP7_75t_L g602 ( 
.A(n_464),
.Y(n_602)
);

OR2x2_ASAP7_75t_SL g603 ( 
.A(n_497),
.B(n_380),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_516),
.B(n_303),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_496),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_511),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_449),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_444),
.B(n_439),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_457),
.B(n_198),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_446),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_511),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_457),
.B(n_182),
.Y(n_612)
);

OR2x6_ASAP7_75t_L g613 ( 
.A(n_495),
.B(n_509),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_458),
.B(n_183),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_496),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_516),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_451),
.B(n_459),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_517),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_497),
.A2(n_275),
.B1(n_266),
.B2(n_264),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_466),
.B(n_402),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_517),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_517),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_458),
.B(n_184),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_464),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_496),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_503),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_464),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_496),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_496),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_493),
.B(n_392),
.Y(n_630)
);

INVx6_ASAP7_75t_L g631 ( 
.A(n_496),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_463),
.B(n_234),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_461),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_469),
.B(n_402),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_483),
.B(n_402),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_461),
.B(n_185),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_509),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_498),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_498),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_498),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_504),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_498),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_498),
.B(n_261),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_492),
.B(n_412),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_498),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_463),
.B(n_234),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_465),
.B(n_304),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_461),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_465),
.B(n_311),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_498),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_508),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_508),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_494),
.B(n_413),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_501),
.B(n_374),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_464),
.Y(n_655)
);

BUFx4f_ASAP7_75t_L g656 ( 
.A(n_508),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_464),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_515),
.B(n_252),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_508),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_508),
.B(n_261),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_513),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_508),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_464),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_508),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_512),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_504),
.Y(n_666)
);

BUFx4f_ASAP7_75t_L g667 ( 
.A(n_512),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_512),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_477),
.B(n_254),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_512),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_666),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_529),
.B(n_512),
.Y(n_672)
);

NOR2xp67_ASAP7_75t_SL g673 ( 
.A(n_578),
.B(n_584),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_529),
.B(n_512),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_546),
.B(n_290),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_539),
.B(n_512),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_564),
.B(n_464),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_541),
.B(n_472),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_553),
.B(n_199),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_520),
.Y(n_680)
);

A2O1A1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_523),
.A2(n_468),
.B(n_325),
.C(n_327),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_568),
.B(n_472),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_538),
.B(n_586),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_550),
.B(n_518),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_608),
.B(n_350),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_521),
.B(n_472),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_549),
.B(n_383),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_521),
.B(n_472),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_519),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_538),
.B(n_350),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_520),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_525),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_561),
.B(n_472),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_593),
.B(n_186),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_599),
.B(n_276),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_599),
.B(n_291),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_546),
.B(n_290),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_534),
.B(n_294),
.Y(n_698)
);

NOR2x1p5_ASAP7_75t_L g699 ( 
.A(n_548),
.B(n_630),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_592),
.B(n_472),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_597),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_530),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_613),
.B(n_477),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_546),
.B(n_290),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_549),
.B(n_472),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_526),
.A2(n_468),
.B(n_505),
.C(n_502),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_601),
.A2(n_578),
.B1(n_584),
.B2(n_569),
.Y(n_707)
);

NOR2xp67_ASAP7_75t_L g708 ( 
.A(n_617),
.B(n_644),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_569),
.A2(n_388),
.B1(n_421),
.B2(n_411),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_534),
.B(n_299),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_637),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_533),
.B(n_477),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_535),
.B(n_257),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_632),
.B(n_190),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_597),
.Y(n_715)
);

AND2x2_ASAP7_75t_SL g716 ( 
.A(n_658),
.B(n_290),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_558),
.B(n_475),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_534),
.A2(n_339),
.B1(n_321),
.B2(n_315),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_534),
.A2(n_391),
.B1(n_407),
.B2(n_247),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_545),
.B(n_302),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_560),
.B(n_479),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_569),
.A2(n_241),
.B1(n_243),
.B2(n_347),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_563),
.B(n_475),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_545),
.B(n_305),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_575),
.B(n_475),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_524),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_577),
.B(n_475),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_545),
.A2(n_339),
.B1(n_321),
.B2(n_315),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_632),
.B(n_191),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_545),
.B(n_306),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_583),
.B(n_475),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_548),
.B(n_479),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_537),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_542),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_606),
.B(n_611),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_666),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_597),
.B(n_475),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_543),
.B(n_669),
.Y(n_738)
);

BUFx6f_ASAP7_75t_SL g739 ( 
.A(n_613),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_542),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_540),
.B(n_607),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_547),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_526),
.A2(n_646),
.B(n_528),
.C(n_579),
.Y(n_743)
);

NOR2xp67_ASAP7_75t_L g744 ( 
.A(n_653),
.B(n_479),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_633),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_669),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_572),
.A2(n_290),
.B1(n_316),
.B2(n_257),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_633),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_633),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_646),
.B(n_193),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_573),
.B(n_201),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_569),
.A2(n_612),
.B1(n_623),
.B2(n_614),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_648),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_619),
.B(n_312),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_L g755 ( 
.A(n_620),
.B(n_499),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_648),
.B(n_475),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_540),
.B(n_204),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_648),
.B(n_499),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_528),
.B(n_316),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_532),
.B(n_205),
.Y(n_760)
);

BUFx12f_ASAP7_75t_L g761 ( 
.A(n_547),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_556),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_528),
.B(n_499),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_641),
.B(n_500),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_572),
.A2(n_316),
.B1(n_272),
.B2(n_337),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_536),
.B(n_500),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_630),
.B(n_500),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_636),
.A2(n_233),
.B1(n_228),
.B2(n_227),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_544),
.Y(n_769)
);

OR2x6_ASAP7_75t_L g770 ( 
.A(n_613),
.B(n_502),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_544),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_536),
.B(n_502),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_637),
.B(n_505),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_536),
.A2(n_316),
.B1(n_272),
.B2(n_257),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_634),
.B(n_210),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_579),
.B(n_505),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_609),
.A2(n_232),
.B1(n_220),
.B2(n_219),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_589),
.B(n_507),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_579),
.B(n_507),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_552),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_522),
.B(n_668),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_600),
.B(n_507),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_635),
.B(n_313),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_600),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_554),
.B(n_320),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_647),
.A2(n_257),
.B1(n_272),
.B2(n_337),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_L g787 ( 
.A(n_647),
.B(n_338),
.C(n_348),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_656),
.A2(n_473),
.B(n_462),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_527),
.B(n_211),
.Y(n_789)
);

OAI221xp5_ASAP7_75t_L g790 ( 
.A1(n_649),
.A2(n_474),
.B1(n_467),
.B2(n_471),
.C(n_470),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_613),
.B(n_591),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_616),
.B(n_462),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_618),
.B(n_621),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_624),
.B(n_257),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_649),
.B(n_341),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_610),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_622),
.B(n_462),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_551),
.B(n_473),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_604),
.B(n_216),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_551),
.B(n_473),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_604),
.A2(n_222),
.B1(n_217),
.B2(n_343),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_571),
.Y(n_802)
);

NOR2xp67_ASAP7_75t_L g803 ( 
.A(n_654),
.B(n_467),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_604),
.A2(n_344),
.B1(n_471),
.B2(n_470),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_552),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_551),
.B(n_474),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_559),
.B(n_221),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_598),
.A2(n_337),
.B1(n_257),
.B2(n_272),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_559),
.B(n_231),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_559),
.B(n_236),
.Y(n_810)
);

NAND2x1_ASAP7_75t_L g811 ( 
.A(n_557),
.B(n_596),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_656),
.B(n_237),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_598),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_565),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_656),
.B(n_240),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_626),
.B(n_6),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_565),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_667),
.B(n_248),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_556),
.B(n_250),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_556),
.B(n_258),
.Y(n_820)
);

INVxp33_ASAP7_75t_SL g821 ( 
.A(n_661),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_603),
.B(n_259),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_603),
.B(n_262),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_598),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_566),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_598),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_566),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_624),
.B(n_272),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_556),
.B(n_263),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_627),
.B(n_272),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_639),
.B(n_659),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_625),
.A2(n_628),
.B1(n_640),
.B2(n_664),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_627),
.B(n_663),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_L g834 ( 
.A(n_643),
.B(n_292),
.C(n_333),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_531),
.B(n_332),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_642),
.A2(n_282),
.B1(n_330),
.B2(n_328),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_667),
.B(n_281),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_531),
.B(n_279),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_567),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_610),
.B(n_297),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_531),
.B(n_280),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_827),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_745),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_684),
.B(n_667),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_683),
.A2(n_643),
.B(n_660),
.C(n_570),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_682),
.A2(n_555),
.B(n_665),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_679),
.A2(n_645),
.B(n_662),
.C(n_650),
.Y(n_847)
);

CKINVDCx10_ASAP7_75t_R g848 ( 
.A(n_739),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_827),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_684),
.B(n_679),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_707),
.A2(n_557),
.B1(n_660),
.B2(n_659),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_716),
.A2(n_557),
.B1(n_567),
.B2(n_576),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_681),
.A2(n_690),
.B(n_804),
.C(n_743),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_685),
.B(n_639),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_711),
.Y(n_855)
);

BUFx12f_ASAP7_75t_L g856 ( 
.A(n_761),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_676),
.A2(n_555),
.B(n_665),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_742),
.Y(n_858)
);

NOR2x1p5_ASAP7_75t_L g859 ( 
.A(n_741),
.B(n_267),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_716),
.A2(n_808),
.B1(n_774),
.B2(n_813),
.Y(n_860)
);

NOR2x1_ASAP7_75t_L g861 ( 
.A(n_708),
.B(n_651),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_685),
.B(n_581),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_687),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_693),
.A2(n_652),
.B(n_663),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_700),
.A2(n_555),
.B(n_665),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_701),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_705),
.A2(n_615),
.B(n_605),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_745),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_752),
.A2(n_557),
.B1(n_596),
.B2(n_631),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_821),
.B(n_671),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_678),
.B(n_581),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_784),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_701),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_695),
.B(n_581),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_715),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_686),
.A2(n_688),
.B(n_677),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_675),
.A2(n_576),
.B(n_585),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_672),
.A2(n_615),
.B(n_605),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_715),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_674),
.A2(n_615),
.B(n_605),
.Y(n_880)
);

OAI321xp33_ASAP7_75t_L g881 ( 
.A1(n_808),
.A2(n_322),
.A3(n_570),
.B1(n_585),
.B2(n_587),
.C(n_590),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_804),
.A2(n_587),
.B(n_590),
.C(n_595),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_748),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_675),
.A2(n_595),
.B(n_655),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_781),
.A2(n_638),
.B(n_629),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_763),
.A2(n_638),
.B(n_629),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_695),
.B(n_582),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_790),
.A2(n_655),
.B(n_582),
.C(n_273),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_766),
.A2(n_776),
.B(n_772),
.Y(n_889)
);

INVx4_ASAP7_75t_L g890 ( 
.A(n_745),
.Y(n_890)
);

AOI21x1_ASAP7_75t_L g891 ( 
.A1(n_833),
.A2(n_631),
.B(n_596),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_736),
.B(n_629),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_745),
.Y(n_893)
);

BUFx4f_ASAP7_75t_L g894 ( 
.A(n_791),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_696),
.B(n_582),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_803),
.B(n_670),
.Y(n_896)
);

AO22x1_ASAP7_75t_L g897 ( 
.A1(n_785),
.A2(n_300),
.B1(n_271),
.B2(n_274),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_767),
.Y(n_898)
);

AND2x2_ASAP7_75t_SL g899 ( 
.A(n_840),
.B(n_322),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_779),
.A2(n_638),
.B(n_562),
.Y(n_900)
);

OAI21x1_ASAP7_75t_L g901 ( 
.A1(n_737),
.A2(n_655),
.B(n_631),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_809),
.A2(n_562),
.B(n_574),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_831),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_696),
.B(n_562),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_810),
.A2(n_574),
.B(n_588),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_795),
.B(n_574),
.Y(n_906)
);

NAND3xp33_ASAP7_75t_L g907 ( 
.A(n_754),
.B(n_319),
.C(n_277),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_795),
.B(n_588),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_732),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_738),
.B(n_588),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_744),
.B(n_670),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_838),
.A2(n_670),
.B(n_657),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_738),
.B(n_670),
.Y(n_913)
);

OAI21x1_ASAP7_75t_L g914 ( 
.A1(n_756),
.A2(n_631),
.B(n_596),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_749),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_746),
.B(n_314),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_689),
.B(n_309),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_774),
.A2(n_298),
.B1(n_285),
.B2(n_268),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_783),
.B(n_322),
.Y(n_919)
);

AOI21x1_ASAP7_75t_L g920 ( 
.A1(n_697),
.A2(n_657),
.B(n_602),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_692),
.B(n_337),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_694),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_783),
.B(n_11),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_697),
.A2(n_657),
.B(n_602),
.Y(n_924)
);

NOR2x1p5_ASAP7_75t_SL g925 ( 
.A(n_753),
.B(n_680),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_831),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_712),
.Y(n_927)
);

AOI21x1_ASAP7_75t_L g928 ( 
.A1(n_704),
.A2(n_657),
.B(n_602),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_SL g929 ( 
.A1(n_704),
.A2(n_272),
.B(n_337),
.C(n_20),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_SL g930 ( 
.A(n_718),
.B(n_337),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_758),
.A2(n_657),
.B(n_602),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_841),
.A2(n_602),
.B(n_594),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_782),
.A2(n_594),
.B(n_580),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_773),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_754),
.A2(n_15),
.B(n_16),
.C(n_20),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_702),
.B(n_337),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_748),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_764),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_712),
.Y(n_939)
);

BUFx4f_ASAP7_75t_L g940 ( 
.A(n_703),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_703),
.B(n_89),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_735),
.B(n_594),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_721),
.B(n_594),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_778),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_762),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_819),
.A2(n_594),
.B(n_580),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_816),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_699),
.B(n_16),
.Y(n_948)
);

INVx5_ASAP7_75t_L g949 ( 
.A(n_762),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_820),
.A2(n_580),
.B(n_95),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_721),
.B(n_580),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_691),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_829),
.A2(n_580),
.B(n_84),
.Y(n_953)
);

OR2x6_ASAP7_75t_L g954 ( 
.A(n_796),
.B(n_24),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_703),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_762),
.A2(n_806),
.B(n_798),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_755),
.B(n_25),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_835),
.B(n_26),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_673),
.A2(n_106),
.B1(n_164),
.B2(n_159),
.Y(n_959)
);

AOI21x1_ASAP7_75t_L g960 ( 
.A1(n_800),
.A2(n_74),
.B(n_156),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_762),
.A2(n_167),
.B(n_153),
.Y(n_961)
);

NAND3xp33_ASAP7_75t_L g962 ( 
.A(n_785),
.B(n_28),
.C(n_29),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_706),
.A2(n_138),
.B(n_135),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_832),
.A2(n_133),
.B1(n_131),
.B2(n_119),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_792),
.A2(n_118),
.B(n_111),
.Y(n_965)
);

BUFx12f_ASAP7_75t_L g966 ( 
.A(n_802),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_835),
.B(n_30),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_825),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_698),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_969)
);

BUFx4f_ASAP7_75t_L g970 ( 
.A(n_770),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_793),
.A2(n_811),
.B(n_717),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_797),
.A2(n_110),
.B(n_98),
.Y(n_972)
);

AOI21xp33_ASAP7_75t_L g973 ( 
.A1(n_698),
.A2(n_39),
.B(n_40),
.Y(n_973)
);

AOI21xp33_ASAP7_75t_L g974 ( 
.A1(n_710),
.A2(n_39),
.B(n_40),
.Y(n_974)
);

NOR3xp33_ASAP7_75t_L g975 ( 
.A(n_709),
.B(n_751),
.C(n_823),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_796),
.B(n_45),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_710),
.B(n_46),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_720),
.A2(n_50),
.B(n_46),
.C(n_47),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_723),
.A2(n_731),
.B(n_727),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_770),
.B(n_826),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_726),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_720),
.B(n_730),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_770),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_757),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_839),
.B(n_740),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_725),
.A2(n_812),
.B(n_815),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_759),
.A2(n_750),
.B(n_714),
.C(n_729),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_739),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_733),
.B(n_814),
.Y(n_989)
);

NOR2x1p5_ASAP7_75t_L g990 ( 
.A(n_787),
.B(n_728),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_734),
.B(n_805),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_759),
.A2(n_794),
.B(n_830),
.Y(n_992)
);

AOI21x1_ASAP7_75t_L g993 ( 
.A1(n_794),
.A2(n_828),
.B(n_830),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_818),
.A2(n_837),
.B(n_807),
.Y(n_994)
);

BUFx4f_ASAP7_75t_L g995 ( 
.A(n_769),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_747),
.A2(n_786),
.B1(n_807),
.B2(n_822),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_788),
.A2(n_828),
.B(n_771),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_780),
.A2(n_817),
.B(n_713),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_789),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_799),
.A2(n_834),
.B(n_775),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_777),
.B(n_730),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_760),
.B(n_823),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_724),
.B(n_768),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_724),
.B(n_836),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_824),
.A2(n_718),
.B(n_728),
.C(n_801),
.Y(n_1005)
);

AOI21xp33_ASAP7_75t_L g1006 ( 
.A1(n_822),
.A2(n_722),
.B(n_824),
.Y(n_1006)
);

OAI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_719),
.A2(n_786),
.B(n_765),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_747),
.A2(n_683),
.B(n_684),
.C(n_679),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_765),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_679),
.A2(n_684),
.B(n_541),
.C(n_553),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_682),
.A2(n_546),
.B(n_561),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_682),
.A2(n_546),
.B(n_561),
.Y(n_1012)
);

NAND3xp33_ASAP7_75t_L g1013 ( 
.A(n_679),
.B(n_553),
.C(n_541),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_711),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_684),
.B(n_679),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_682),
.A2(n_546),
.B(n_561),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_827),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_693),
.A2(n_592),
.B(n_561),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_682),
.A2(n_546),
.B(n_561),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_784),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_682),
.A2(n_546),
.B(n_561),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_682),
.A2(n_546),
.B(n_561),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_679),
.A2(n_684),
.B(n_541),
.C(n_553),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_682),
.A2(n_546),
.B(n_561),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_684),
.B(n_716),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_693),
.A2(n_592),
.B(n_561),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_745),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_827),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_827),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_784),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_682),
.A2(n_546),
.B(n_561),
.Y(n_1031)
);

BUFx8_ASAP7_75t_L g1032 ( 
.A(n_739),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_934),
.B(n_938),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_850),
.B(n_1015),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_1010),
.A2(n_1023),
.B(n_1013),
.C(n_923),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1018),
.B(n_1026),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_855),
.Y(n_1037)
);

OAI22x1_ASAP7_75t_L g1038 ( 
.A1(n_990),
.A2(n_982),
.B1(n_919),
.B2(n_980),
.Y(n_1038)
);

AOI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_1008),
.A2(n_1003),
.B(n_1001),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_968),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_876),
.A2(n_889),
.B(n_906),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_934),
.B(n_944),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_855),
.B(n_870),
.Y(n_1043)
);

O2A1O1Ixp5_ASAP7_75t_L g1044 ( 
.A1(n_958),
.A2(n_967),
.B(n_1025),
.C(n_844),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_908),
.A2(n_904),
.B(n_949),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_1014),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_945),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1018),
.B(n_1026),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_860),
.A2(n_996),
.B1(n_1009),
.B2(n_1007),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_913),
.B(n_910),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_949),
.A2(n_994),
.B(n_1011),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_1012),
.A2(n_1019),
.B(n_1016),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_860),
.A2(n_1004),
.B1(n_852),
.B2(n_1002),
.Y(n_1053)
);

AO221x2_ASAP7_75t_L g1054 ( 
.A1(n_962),
.A2(n_897),
.B1(n_965),
.B2(n_972),
.C(n_963),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_863),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_849),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_890),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_949),
.A2(n_1022),
.B(n_1021),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_949),
.A2(n_1031),
.B(n_1024),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_891),
.A2(n_901),
.B(n_914),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_SL g1061 ( 
.A1(n_963),
.A2(n_853),
.B(n_965),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_909),
.B(n_898),
.Y(n_1062)
);

NAND2x1_ASAP7_75t_L g1063 ( 
.A(n_890),
.B(n_1027),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_983),
.B(n_980),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_892),
.B(n_977),
.Y(n_1065)
);

NOR2xp67_ASAP7_75t_L g1066 ( 
.A(n_907),
.B(n_984),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_997),
.A2(n_846),
.B(n_956),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_878),
.A2(n_880),
.B(n_905),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_976),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_865),
.A2(n_857),
.B(n_867),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_975),
.A2(n_1006),
.B1(n_930),
.B2(n_939),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_926),
.B(n_927),
.Y(n_1072)
);

AOI21x1_ASAP7_75t_L g1073 ( 
.A1(n_920),
.A2(n_928),
.B(n_895),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_864),
.A2(n_979),
.B(n_851),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_871),
.A2(n_986),
.B(n_885),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_926),
.B(n_854),
.Y(n_1076)
);

AO31x2_ASAP7_75t_L g1077 ( 
.A1(n_847),
.A2(n_852),
.A3(n_874),
.B(n_887),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_987),
.A2(n_888),
.B(n_1005),
.C(n_1000),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_983),
.B(n_955),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_947),
.B(n_899),
.Y(n_1080)
);

NAND3xp33_ASAP7_75t_L g1081 ( 
.A(n_930),
.B(n_973),
.C(n_974),
.Y(n_1081)
);

INVxp67_ASAP7_75t_SL g1082 ( 
.A(n_945),
.Y(n_1082)
);

AOI211x1_ASAP7_75t_L g1083 ( 
.A1(n_972),
.A2(n_915),
.B(n_992),
.C(n_1030),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_872),
.B(n_1020),
.Y(n_1084)
);

AOI21x1_ASAP7_75t_SL g1085 ( 
.A1(n_957),
.A2(n_948),
.B(n_942),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_903),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_902),
.A2(n_912),
.B(n_993),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_858),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_945),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_903),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_862),
.B(n_866),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_999),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_966),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_873),
.B(n_875),
.Y(n_1094)
);

O2A1O1Ixp5_ASAP7_75t_L g1095 ( 
.A1(n_896),
.A2(n_911),
.B(n_924),
.C(n_933),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_1002),
.B(n_917),
.Y(n_1096)
);

AOI221xp5_ASAP7_75t_L g1097 ( 
.A1(n_935),
.A2(n_922),
.B1(n_918),
.B2(n_969),
.C(n_978),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_903),
.B(n_940),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_886),
.A2(n_900),
.B(n_971),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_864),
.A2(n_881),
.B(n_992),
.Y(n_1100)
);

AO21x1_ASAP7_75t_L g1101 ( 
.A1(n_884),
.A2(n_964),
.B(n_921),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_933),
.A2(n_931),
.B(n_943),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_931),
.A2(n_951),
.B(n_884),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_894),
.A2(n_916),
.B1(n_859),
.B2(n_941),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_879),
.B(n_937),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_932),
.A2(n_946),
.B(n_877),
.Y(n_1106)
);

AOI21x1_ASAP7_75t_L g1107 ( 
.A1(n_936),
.A2(n_985),
.B(n_877),
.Y(n_1107)
);

AO21x1_ASAP7_75t_L g1108 ( 
.A1(n_882),
.A2(n_924),
.B(n_845),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_SL g1109 ( 
.A1(n_959),
.A2(n_941),
.B(n_918),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_SL g1110 ( 
.A(n_954),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_883),
.B(n_894),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_952),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_1027),
.B(n_843),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1017),
.B(n_1029),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_998),
.A2(n_989),
.B(n_991),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_950),
.A2(n_953),
.B(n_869),
.Y(n_1116)
);

INVx4_ASAP7_75t_L g1117 ( 
.A(n_843),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_940),
.B(n_970),
.Y(n_1118)
);

AO31x2_ASAP7_75t_L g1119 ( 
.A1(n_1028),
.A2(n_981),
.A3(n_961),
.B(n_881),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_861),
.A2(n_960),
.B(n_925),
.Y(n_1120)
);

OAI21xp33_ASAP7_75t_L g1121 ( 
.A1(n_954),
.A2(n_843),
.B(n_868),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_868),
.A2(n_893),
.B(n_995),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_L g1123 ( 
.A1(n_995),
.A2(n_868),
.B(n_893),
.Y(n_1123)
);

AOI21x1_ASAP7_75t_SL g1124 ( 
.A1(n_929),
.A2(n_970),
.B(n_893),
.Y(n_1124)
);

O2A1O1Ixp5_ASAP7_75t_L g1125 ( 
.A1(n_954),
.A2(n_988),
.B(n_1032),
.C(n_848),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1032),
.B(n_856),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_891),
.A2(n_901),
.B(n_914),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_1014),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_983),
.B(n_980),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_903),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1013),
.B(n_1010),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_L g1132 ( 
.A(n_1013),
.B(n_1023),
.C(n_1010),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_890),
.Y(n_1133)
);

AO31x2_ASAP7_75t_L g1134 ( 
.A1(n_847),
.A2(n_996),
.A3(n_851),
.B(n_852),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_850),
.B(n_1015),
.Y(n_1135)
);

NOR2x1_ASAP7_75t_SL g1136 ( 
.A(n_949),
.B(n_945),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1013),
.B(n_1010),
.Y(n_1137)
);

AOI21x1_ASAP7_75t_L g1138 ( 
.A1(n_844),
.A2(n_928),
.B(n_920),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_876),
.A2(n_546),
.B(n_561),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_876),
.A2(n_546),
.B(n_561),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_891),
.A2(n_901),
.B(n_914),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_842),
.Y(n_1142)
);

AOI21xp33_ASAP7_75t_L g1143 ( 
.A1(n_1013),
.A2(n_1015),
.B(n_850),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1010),
.A2(n_1023),
.B(n_1013),
.C(n_1015),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_850),
.B(n_1015),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_855),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_876),
.A2(n_546),
.B(n_561),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_SL g1148 ( 
.A1(n_963),
.A2(n_853),
.B(n_965),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_1014),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1010),
.A2(n_1023),
.B1(n_1015),
.B2(n_850),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1010),
.A2(n_1023),
.B(n_1012),
.Y(n_1151)
);

NOR2x1_ASAP7_75t_L g1152 ( 
.A(n_858),
.B(n_1013),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1010),
.A2(n_1023),
.B(n_1012),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_891),
.A2(n_901),
.B(n_914),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_1014),
.B(n_761),
.Y(n_1155)
);

OR2x6_ASAP7_75t_L g1156 ( 
.A(n_1014),
.B(n_761),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_891),
.A2(n_901),
.B(n_914),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_850),
.B(n_1015),
.Y(n_1158)
);

NAND3xp33_ASAP7_75t_SL g1159 ( 
.A(n_1013),
.B(n_1023),
.C(n_1010),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_850),
.B(n_1015),
.Y(n_1160)
);

NAND2xp33_ASAP7_75t_L g1161 ( 
.A(n_850),
.B(n_1015),
.Y(n_1161)
);

AND3x2_ASAP7_75t_L g1162 ( 
.A(n_930),
.B(n_923),
.C(n_658),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_891),
.A2(n_901),
.B(n_914),
.Y(n_1163)
);

AOI21xp33_ASAP7_75t_L g1164 ( 
.A1(n_1013),
.A2(n_1015),
.B(n_850),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_890),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_876),
.A2(n_546),
.B(n_561),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1013),
.B(n_1010),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_934),
.B(n_938),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1010),
.A2(n_1023),
.B(n_1012),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_891),
.A2(n_901),
.B(n_914),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_850),
.B(n_1015),
.Y(n_1171)
);

INVxp67_ASAP7_75t_SL g1172 ( 
.A(n_945),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_947),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1010),
.A2(n_1023),
.B(n_1012),
.Y(n_1174)
);

INVx5_ASAP7_75t_L g1175 ( 
.A(n_945),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1013),
.B(n_1010),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_890),
.Y(n_1177)
);

OA21x2_ASAP7_75t_L g1178 ( 
.A1(n_864),
.A2(n_1026),
.B(n_1018),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_876),
.A2(n_546),
.B(n_561),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_850),
.B(n_1015),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_876),
.A2(n_546),
.B(n_561),
.Y(n_1181)
);

AOI21xp33_ASAP7_75t_L g1182 ( 
.A1(n_1013),
.A2(n_1015),
.B(n_850),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1010),
.A2(n_1023),
.B(n_1012),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_876),
.A2(n_546),
.B(n_561),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_891),
.A2(n_901),
.B(n_914),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_842),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_855),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1034),
.B(n_1135),
.Y(n_1188)
);

CKINVDCx6p67_ASAP7_75t_R g1189 ( 
.A(n_1088),
.Y(n_1189)
);

BUFx12f_ASAP7_75t_L g1190 ( 
.A(n_1093),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1060),
.A2(n_1141),
.B(n_1127),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1033),
.B(n_1168),
.Y(n_1192)
);

BUFx4f_ASAP7_75t_L g1193 ( 
.A(n_1155),
.Y(n_1193)
);

O2A1O1Ixp5_ASAP7_75t_SL g1194 ( 
.A1(n_1131),
.A2(n_1167),
.B(n_1137),
.C(n_1176),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1035),
.A2(n_1081),
.B(n_1132),
.C(n_1144),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1040),
.Y(n_1196)
);

BUFx4_ASAP7_75t_SL g1197 ( 
.A(n_1155),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1037),
.B(n_1034),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1187),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1113),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1069),
.B(n_1043),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1041),
.A2(n_1074),
.B(n_1075),
.Y(n_1202)
);

BUFx12f_ASAP7_75t_L g1203 ( 
.A(n_1155),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1074),
.A2(n_1099),
.B(n_1061),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1143),
.A2(n_1164),
.B(n_1182),
.C(n_1039),
.Y(n_1205)
);

INVx5_ASAP7_75t_L g1206 ( 
.A(n_1047),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1161),
.A2(n_1160),
.B(n_1171),
.C(n_1145),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1148),
.A2(n_1070),
.B(n_1052),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1156),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1084),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1037),
.B(n_1158),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1180),
.B(n_1143),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1164),
.B(n_1182),
.Y(n_1213)
);

INVx3_ASAP7_75t_SL g1214 ( 
.A(n_1156),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1069),
.B(n_1055),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1146),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_SL g1217 ( 
.A(n_1156),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1112),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1045),
.A2(n_1166),
.B(n_1184),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1080),
.B(n_1042),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1052),
.A2(n_1179),
.B(n_1147),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1110),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1046),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1128),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1039),
.A2(n_1109),
.B(n_1096),
.C(n_1159),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1149),
.Y(n_1226)
);

AO22x1_ASAP7_75t_L g1227 ( 
.A1(n_1111),
.A2(n_1152),
.B1(n_1064),
.B2(n_1129),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1047),
.Y(n_1228)
);

INVx3_ASAP7_75t_SL g1229 ( 
.A(n_1079),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1173),
.B(n_1092),
.Y(n_1230)
);

INVx5_ASAP7_75t_L g1231 ( 
.A(n_1047),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1150),
.B(n_1050),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1079),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1064),
.B(n_1129),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1139),
.A2(n_1181),
.B(n_1140),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1038),
.B(n_1104),
.Y(n_1236)
);

OR2x6_ASAP7_75t_L g1237 ( 
.A(n_1118),
.B(n_1098),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1150),
.B(n_1050),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1062),
.B(n_1056),
.Y(n_1239)
);

INVx5_ASAP7_75t_L g1240 ( 
.A(n_1089),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1094),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1114),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1090),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1054),
.A2(n_1110),
.B1(n_1053),
.B2(n_1049),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1151),
.A2(n_1174),
.B(n_1183),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_1089),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1049),
.A2(n_1071),
.B1(n_1036),
.B2(n_1048),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1153),
.A2(n_1174),
.B(n_1169),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1036),
.A2(n_1048),
.B1(n_1109),
.B2(n_1053),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1065),
.B(n_1162),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_1126),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1121),
.B(n_1072),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1090),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1051),
.A2(n_1078),
.B(n_1102),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1066),
.B(n_1186),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1058),
.A2(n_1059),
.B(n_1103),
.Y(n_1256)
);

NOR2x1_ASAP7_75t_L g1257 ( 
.A(n_1117),
.B(n_1130),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1082),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1100),
.A2(n_1067),
.B(n_1068),
.Y(n_1259)
);

INVx3_ASAP7_75t_SL g1260 ( 
.A(n_1086),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1142),
.Y(n_1261)
);

BUFx4_ASAP7_75t_SL g1262 ( 
.A(n_1125),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1086),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1126),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1130),
.B(n_1117),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1175),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1105),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1175),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1076),
.B(n_1091),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1175),
.B(n_1172),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1100),
.A2(n_1178),
.B(n_1054),
.Y(n_1271)
);

O2A1O1Ixp5_ASAP7_75t_L g1272 ( 
.A1(n_1044),
.A2(n_1101),
.B(n_1108),
.C(n_1095),
.Y(n_1272)
);

INVxp67_ASAP7_75t_SL g1273 ( 
.A(n_1136),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1091),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1154),
.A2(n_1185),
.B(n_1170),
.Y(n_1275)
);

AOI21xp33_ASAP7_75t_L g1276 ( 
.A1(n_1097),
.A2(n_1178),
.B(n_1116),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1115),
.A2(n_1107),
.B(n_1106),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1122),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_SL g1279 ( 
.A(n_1057),
.B(n_1177),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1123),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1083),
.A2(n_1165),
.B1(n_1133),
.B2(n_1177),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1165),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1119),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1063),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1134),
.A2(n_1138),
.B1(n_1073),
.B2(n_1124),
.Y(n_1285)
);

INVxp67_ASAP7_75t_SL g1286 ( 
.A(n_1120),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1134),
.B(n_1119),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1119),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1085),
.Y(n_1289)
);

OAI21xp33_ASAP7_75t_L g1290 ( 
.A1(n_1087),
.A2(n_1157),
.B(n_1163),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1134),
.B(n_1077),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1077),
.B(n_1034),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1077),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1187),
.Y(n_1294)
);

NAND2xp33_ASAP7_75t_L g1295 ( 
.A(n_1035),
.B(n_1010),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1041),
.A2(n_1074),
.B(n_1075),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1187),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1034),
.B(n_1135),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1034),
.B(n_1135),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1155),
.B(n_1156),
.Y(n_1300)
);

CKINVDCx16_ASAP7_75t_R g1301 ( 
.A(n_1088),
.Y(n_1301)
);

AOI221xp5_ASAP7_75t_L g1302 ( 
.A1(n_1049),
.A2(n_1013),
.B1(n_1023),
.B2(n_1010),
.C(n_982),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1034),
.B(n_1135),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1187),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1034),
.B(n_1135),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1135),
.B(n_1013),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1151),
.A2(n_1169),
.B(n_1153),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1040),
.Y(n_1308)
);

INVx3_ASAP7_75t_SL g1309 ( 
.A(n_1155),
.Y(n_1309)
);

NAND2x1_ASAP7_75t_L g1310 ( 
.A(n_1057),
.B(n_890),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1035),
.A2(n_1023),
.B(n_1010),
.C(n_1013),
.Y(n_1311)
);

AO21x2_ASAP7_75t_L g1312 ( 
.A1(n_1074),
.A2(n_1148),
.B(n_1061),
.Y(n_1312)
);

OR2x6_ASAP7_75t_L g1313 ( 
.A(n_1155),
.B(n_1156),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1113),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1041),
.A2(n_1074),
.B(n_1075),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1034),
.A2(n_1010),
.B1(n_1023),
.B2(n_1015),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1033),
.B(n_934),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1034),
.B(n_1135),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1187),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1041),
.A2(n_1074),
.B(n_1075),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1033),
.B(n_934),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1034),
.B(n_1135),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1135),
.B(n_1013),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1040),
.Y(n_1324)
);

CKINVDCx11_ASAP7_75t_R g1325 ( 
.A(n_1155),
.Y(n_1325)
);

CKINVDCx11_ASAP7_75t_R g1326 ( 
.A(n_1155),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1064),
.B(n_1129),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1047),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1080),
.A2(n_1013),
.B1(n_982),
.B2(n_919),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1040),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1329),
.A2(n_1188),
.B1(n_1305),
.B2(n_1322),
.Y(n_1331)
);

AO21x2_ASAP7_75t_L g1332 ( 
.A1(n_1259),
.A2(n_1221),
.B(n_1277),
.Y(n_1332)
);

BUFx2_ASAP7_75t_R g1333 ( 
.A(n_1222),
.Y(n_1333)
);

AO21x2_ASAP7_75t_L g1334 ( 
.A1(n_1221),
.A2(n_1277),
.B(n_1256),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1327),
.B(n_1237),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1196),
.Y(n_1336)
);

NAND2x1p5_ASAP7_75t_L g1337 ( 
.A(n_1289),
.B(n_1278),
.Y(n_1337)
);

BUFx2_ASAP7_75t_SL g1338 ( 
.A(n_1206),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1244),
.B(n_1274),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1306),
.A2(n_1323),
.B1(n_1236),
.B2(n_1295),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1302),
.A2(n_1250),
.B1(n_1247),
.B2(n_1316),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1188),
.B(n_1298),
.Y(n_1342)
);

BUFx12f_ASAP7_75t_L g1343 ( 
.A(n_1325),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1302),
.A2(n_1250),
.B1(n_1247),
.B2(n_1316),
.Y(n_1344)
);

AOI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1245),
.A2(n_1248),
.B(n_1204),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1249),
.A2(n_1245),
.B1(n_1252),
.B2(n_1312),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1191),
.A2(n_1235),
.B(n_1219),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1215),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1312),
.A2(n_1212),
.B1(n_1213),
.B2(n_1237),
.Y(n_1349)
);

BUFx4f_ASAP7_75t_SL g1350 ( 
.A(n_1223),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1212),
.A2(n_1213),
.B1(n_1237),
.B2(n_1291),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1291),
.A2(n_1307),
.B1(n_1201),
.B2(n_1220),
.Y(n_1352)
);

BUFx5_ASAP7_75t_L g1353 ( 
.A(n_1287),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1229),
.Y(n_1354)
);

CKINVDCx6p67_ASAP7_75t_R g1355 ( 
.A(n_1217),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1294),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1298),
.A2(n_1305),
.B1(n_1303),
.B2(n_1318),
.Y(n_1357)
);

BUFx8_ASAP7_75t_L g1358 ( 
.A(n_1217),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1193),
.A2(n_1255),
.B1(n_1318),
.B2(n_1299),
.Y(n_1359)
);

INVxp67_ASAP7_75t_SL g1360 ( 
.A(n_1297),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1224),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1319),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1299),
.B(n_1303),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1322),
.A2(n_1210),
.B1(n_1198),
.B2(n_1238),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1317),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1192),
.Y(n_1366)
);

AO21x1_ASAP7_75t_SL g1367 ( 
.A1(n_1232),
.A2(n_1238),
.B(n_1292),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1193),
.A2(n_1300),
.B1(n_1313),
.B2(n_1214),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1324),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1232),
.A2(n_1225),
.B1(n_1211),
.B2(n_1195),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1330),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1269),
.B(n_1241),
.Y(n_1372)
);

INVx4_ASAP7_75t_L g1373 ( 
.A(n_1268),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1218),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1300),
.A2(n_1313),
.B1(n_1292),
.B2(n_1279),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1242),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1307),
.A2(n_1264),
.B1(n_1321),
.B2(n_1304),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1254),
.A2(n_1208),
.B(n_1320),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1199),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1216),
.A2(n_1289),
.B1(n_1203),
.B2(n_1326),
.Y(n_1380)
);

AOI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1204),
.A2(n_1296),
.B(n_1315),
.Y(n_1381)
);

CKINVDCx6p67_ASAP7_75t_R g1382 ( 
.A(n_1309),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1267),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1226),
.Y(n_1384)
);

BUFx2_ASAP7_75t_R g1385 ( 
.A(n_1209),
.Y(n_1385)
);

BUFx12f_ASAP7_75t_L g1386 ( 
.A(n_1190),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1293),
.A2(n_1327),
.B1(n_1271),
.B2(n_1313),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1268),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1206),
.Y(n_1389)
);

INVx4_ASAP7_75t_L g1390 ( 
.A(n_1268),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1230),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1207),
.A2(n_1205),
.B1(n_1233),
.B2(n_1258),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1189),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1239),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1271),
.B(n_1288),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1251),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1300),
.A2(n_1234),
.B1(n_1276),
.B2(n_1261),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1194),
.B(n_1311),
.Y(n_1398)
);

AO21x1_ASAP7_75t_SL g1399 ( 
.A1(n_1276),
.A2(n_1280),
.B(n_1290),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1231),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1200),
.B(n_1314),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1283),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1282),
.Y(n_1403)
);

BUFx2_ASAP7_75t_R g1404 ( 
.A(n_1260),
.Y(n_1404)
);

BUFx8_ASAP7_75t_SL g1405 ( 
.A(n_1243),
.Y(n_1405)
);

CKINVDCx11_ASAP7_75t_R g1406 ( 
.A(n_1301),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1253),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1275),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1202),
.A2(n_1315),
.B(n_1285),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1197),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1314),
.B(n_1227),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1286),
.A2(n_1281),
.B(n_1310),
.Y(n_1412)
);

BUFx4_ASAP7_75t_SL g1413 ( 
.A(n_1266),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1265),
.B(n_1270),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1273),
.A2(n_1265),
.B1(n_1263),
.B2(n_1257),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1246),
.B(n_1279),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1270),
.A2(n_1284),
.B1(n_1328),
.B2(n_1228),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1228),
.A2(n_1328),
.B1(n_1246),
.B2(n_1240),
.Y(n_1418)
);

CKINVDCx11_ASAP7_75t_R g1419 ( 
.A(n_1228),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1231),
.B(n_1240),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1240),
.B(n_1262),
.Y(n_1421)
);

AO21x1_ASAP7_75t_L g1422 ( 
.A1(n_1295),
.A2(n_1311),
.B(n_1150),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1244),
.B(n_1274),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1297),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1297),
.Y(n_1425)
);

INVxp67_ASAP7_75t_L g1426 ( 
.A(n_1201),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1244),
.A2(n_1013),
.B1(n_919),
.B2(n_1054),
.Y(n_1427)
);

INVxp67_ASAP7_75t_SL g1428 ( 
.A(n_1297),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1329),
.A2(n_1013),
.B1(n_982),
.B2(n_919),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1244),
.A2(n_1013),
.B1(n_919),
.B2(n_1054),
.Y(n_1430)
);

INVx8_ASAP7_75t_L g1431 ( 
.A(n_1206),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1244),
.A2(n_1013),
.B1(n_919),
.B2(n_1054),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1308),
.Y(n_1433)
);

NAND2x1p5_ASAP7_75t_L g1434 ( 
.A(n_1289),
.B(n_1278),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1223),
.Y(n_1435)
);

BUFx12f_ASAP7_75t_L g1436 ( 
.A(n_1325),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1197),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1272),
.A2(n_1259),
.B(n_1254),
.Y(n_1438)
);

INVxp33_ASAP7_75t_L g1439 ( 
.A(n_1201),
.Y(n_1439)
);

INVx4_ASAP7_75t_L g1440 ( 
.A(n_1268),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1244),
.A2(n_1013),
.B1(n_919),
.B2(n_1054),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1188),
.B(n_1298),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1201),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1308),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1308),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1353),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1367),
.B(n_1342),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1409),
.A2(n_1378),
.B(n_1347),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1409),
.A2(n_1378),
.B(n_1347),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1424),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1335),
.B(n_1402),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1424),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1367),
.B(n_1342),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1408),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1395),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1395),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1353),
.Y(n_1457)
);

CKINVDCx6p67_ASAP7_75t_R g1458 ( 
.A(n_1406),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1331),
.B(n_1357),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1353),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1406),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1425),
.Y(n_1462)
);

AOI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1381),
.A2(n_1398),
.B(n_1345),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1364),
.B(n_1372),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1339),
.B(n_1423),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1339),
.B(n_1423),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1346),
.B(n_1349),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1425),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1353),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1362),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1353),
.Y(n_1471)
);

AO21x2_ASAP7_75t_L g1472 ( 
.A1(n_1332),
.A2(n_1334),
.B(n_1422),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1439),
.B(n_1366),
.Y(n_1473)
);

OR2x6_ASAP7_75t_L g1474 ( 
.A(n_1337),
.B(n_1434),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1438),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1394),
.Y(n_1476)
);

INVxp67_ASAP7_75t_SL g1477 ( 
.A(n_1422),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1372),
.B(n_1363),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1348),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1341),
.B(n_1344),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1412),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1352),
.B(n_1370),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1351),
.B(n_1365),
.Y(n_1483)
);

INVxp67_ASAP7_75t_SL g1484 ( 
.A(n_1337),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1439),
.B(n_1426),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1434),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1434),
.A2(n_1392),
.B(n_1387),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1360),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1377),
.B(n_1443),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1437),
.Y(n_1490)
);

INVxp67_ASAP7_75t_L g1491 ( 
.A(n_1428),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1411),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1340),
.B(n_1383),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1336),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1427),
.A2(n_1441),
.B(n_1430),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1411),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1416),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1432),
.A2(n_1397),
.B(n_1403),
.Y(n_1498)
);

AO21x2_ASAP7_75t_L g1499 ( 
.A1(n_1429),
.A2(n_1371),
.B(n_1369),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1442),
.B(n_1376),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1391),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1359),
.A2(n_1375),
.B(n_1401),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1399),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1335),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1407),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1445),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1379),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1444),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1433),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1374),
.B(n_1399),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1368),
.A2(n_1435),
.B1(n_1380),
.B2(n_1343),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_SL g1512 ( 
.A(n_1358),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1338),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1389),
.Y(n_1514)
);

BUFx8_ASAP7_75t_SL g1515 ( 
.A(n_1490),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1471),
.B(n_1414),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1471),
.B(n_1414),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1484),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1447),
.B(n_1388),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1447),
.B(n_1355),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1455),
.B(n_1421),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1464),
.B(n_1459),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_SL g1523 ( 
.A1(n_1502),
.A2(n_1415),
.B(n_1400),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1453),
.B(n_1454),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1453),
.B(n_1355),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1472),
.B(n_1420),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1474),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1472),
.B(n_1440),
.Y(n_1528)
);

NOR2x1_ASAP7_75t_L g1529 ( 
.A(n_1499),
.B(n_1440),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1472),
.B(n_1440),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1464),
.B(n_1356),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1472),
.B(n_1373),
.Y(n_1532)
);

AOI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1459),
.A2(n_1393),
.B1(n_1384),
.B2(n_1361),
.C(n_1435),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1455),
.B(n_1382),
.Y(n_1534)
);

NOR2x1_ASAP7_75t_L g1535 ( 
.A(n_1499),
.B(n_1390),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1456),
.B(n_1417),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1457),
.B(n_1460),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1456),
.B(n_1382),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1499),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1495),
.A2(n_1358),
.B1(n_1343),
.B2(n_1436),
.Y(n_1540)
);

INVx5_ASAP7_75t_L g1541 ( 
.A(n_1503),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1481),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1495),
.A2(n_1480),
.B1(n_1482),
.B2(n_1467),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1475),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1477),
.B(n_1418),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1469),
.B(n_1354),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1474),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1499),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1494),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1488),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1469),
.B(n_1354),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1446),
.B(n_1463),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1522),
.B(n_1531),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_SL g1554 ( 
.A1(n_1523),
.A2(n_1495),
.B1(n_1480),
.B2(n_1467),
.Y(n_1554)
);

OAI21xp5_ASAP7_75t_SL g1555 ( 
.A1(n_1540),
.A2(n_1543),
.B(n_1533),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1524),
.B(n_1497),
.Y(n_1556)
);

OAI21xp33_ASAP7_75t_L g1557 ( 
.A1(n_1543),
.A2(n_1482),
.B(n_1465),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1524),
.B(n_1526),
.Y(n_1558)
);

OAI221xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1533),
.A2(n_1511),
.B1(n_1465),
.B2(n_1466),
.C(n_1489),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1540),
.A2(n_1502),
.B(n_1466),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1531),
.A2(n_1495),
.B1(n_1512),
.B2(n_1458),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1521),
.B(n_1479),
.Y(n_1562)
);

NAND3xp33_ASAP7_75t_L g1563 ( 
.A(n_1545),
.B(n_1489),
.C(n_1495),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1521),
.B(n_1501),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1523),
.B(n_1493),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1545),
.A2(n_1512),
.B1(n_1458),
.B2(n_1483),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1549),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1521),
.B(n_1476),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1526),
.B(n_1519),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1550),
.B(n_1462),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_L g1571 ( 
.A(n_1534),
.B(n_1493),
.C(n_1510),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1550),
.B(n_1462),
.Y(n_1572)
);

OA21x2_ASAP7_75t_L g1573 ( 
.A1(n_1539),
.A2(n_1449),
.B(n_1448),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1526),
.B(n_1492),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1529),
.A2(n_1477),
.B(n_1500),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1534),
.B(n_1450),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1538),
.B(n_1468),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1538),
.B(n_1470),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1519),
.B(n_1492),
.Y(n_1579)
);

OAI221xp5_ASAP7_75t_L g1580 ( 
.A1(n_1538),
.A2(n_1485),
.B1(n_1473),
.B2(n_1483),
.C(n_1452),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1546),
.B(n_1491),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1546),
.B(n_1452),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1520),
.B(n_1458),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1551),
.B(n_1478),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1551),
.B(n_1478),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1551),
.B(n_1505),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1529),
.B(n_1451),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1516),
.B(n_1507),
.Y(n_1588)
);

AOI211xp5_ASAP7_75t_SL g1589 ( 
.A1(n_1539),
.A2(n_1486),
.B(n_1510),
.C(n_1504),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1516),
.B(n_1492),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1536),
.A2(n_1396),
.B1(n_1461),
.B2(n_1496),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1516),
.B(n_1496),
.Y(n_1592)
);

NAND2xp33_ASAP7_75t_SL g1593 ( 
.A(n_1520),
.B(n_1503),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1544),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1517),
.B(n_1496),
.Y(n_1595)
);

AOI221xp5_ASAP7_75t_L g1596 ( 
.A1(n_1536),
.A2(n_1500),
.B1(n_1506),
.B2(n_1508),
.C(n_1509),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1518),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1520),
.B(n_1525),
.Y(n_1598)
);

NAND3xp33_ASAP7_75t_L g1599 ( 
.A(n_1535),
.B(n_1498),
.C(n_1514),
.Y(n_1599)
);

NAND3xp33_ASAP7_75t_L g1600 ( 
.A(n_1535),
.B(n_1498),
.C(n_1514),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1541),
.A2(n_1396),
.B1(n_1503),
.B2(n_1504),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1567),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1594),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1567),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1562),
.B(n_1548),
.Y(n_1605)
);

INVx4_ASAP7_75t_L g1606 ( 
.A(n_1573),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1594),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1597),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1558),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1558),
.B(n_1528),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1573),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1570),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1553),
.B(n_1537),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1573),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1572),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1573),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1564),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1569),
.B(n_1528),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1568),
.B(n_1548),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1581),
.B(n_1552),
.Y(n_1620)
);

NOR2xp67_ASAP7_75t_L g1621 ( 
.A(n_1599),
.B(n_1542),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1574),
.B(n_1528),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1556),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1575),
.B(n_1537),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1587),
.B(n_1547),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1579),
.B(n_1530),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1556),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1579),
.B(n_1530),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1583),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1590),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1588),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1592),
.B(n_1530),
.Y(n_1632)
);

AND2x2_ASAP7_75t_SL g1633 ( 
.A(n_1598),
.B(n_1527),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1582),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1578),
.B(n_1525),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1586),
.B(n_1552),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1587),
.B(n_1547),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1595),
.B(n_1532),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1602),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1602),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1608),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1604),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1617),
.B(n_1584),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1603),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1604),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1609),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1609),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1612),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1612),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1624),
.A2(n_1555),
.B(n_1563),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1607),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1633),
.B(n_1589),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1607),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1633),
.B(n_1519),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1603),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1603),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1633),
.B(n_1525),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1617),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1615),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1615),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1625),
.B(n_1571),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1624),
.B(n_1585),
.Y(n_1662)
);

OAI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1629),
.A2(n_1560),
.B1(n_1561),
.B2(n_1580),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1631),
.B(n_1576),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1623),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1618),
.B(n_1610),
.Y(n_1666)
);

NOR2x1p5_ASAP7_75t_L g1667 ( 
.A(n_1629),
.B(n_1436),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1605),
.B(n_1577),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1605),
.B(n_1600),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1623),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1635),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1631),
.B(n_1554),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1625),
.B(n_1547),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1613),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1625),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1627),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1650),
.B(n_1630),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1652),
.B(n_1666),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1639),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1652),
.B(n_1618),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1644),
.Y(n_1681)
);

OR2x6_ASAP7_75t_L g1682 ( 
.A(n_1667),
.B(n_1621),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1675),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1641),
.Y(n_1684)
);

NAND2x1_ASAP7_75t_L g1685 ( 
.A(n_1661),
.B(n_1621),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_SL g1686 ( 
.A(n_1663),
.B(n_1385),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1662),
.B(n_1636),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1671),
.B(n_1630),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1672),
.B(n_1630),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1675),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1664),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1666),
.B(n_1618),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1658),
.B(n_1674),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1640),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1659),
.B(n_1630),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1662),
.B(n_1668),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1663),
.B(n_1629),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1642),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1661),
.B(n_1610),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1645),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1661),
.B(n_1566),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1660),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1648),
.B(n_1632),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1657),
.A2(n_1557),
.B1(n_1565),
.B2(n_1593),
.Y(n_1704)
);

INVxp67_ASAP7_75t_L g1705 ( 
.A(n_1649),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1654),
.B(n_1610),
.Y(n_1706)
);

INVxp67_ASAP7_75t_SL g1707 ( 
.A(n_1675),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1643),
.B(n_1632),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1668),
.B(n_1632),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1651),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1651),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1665),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1654),
.B(n_1622),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1670),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1676),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1653),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1669),
.B(n_1638),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1646),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1669),
.B(n_1636),
.Y(n_1719)
);

AND2x4_ASAP7_75t_SL g1720 ( 
.A(n_1682),
.B(n_1657),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1710),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1684),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1684),
.B(n_1673),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1677),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1711),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1678),
.B(n_1673),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1679),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1678),
.B(n_1673),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1694),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1691),
.B(n_1647),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1699),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1697),
.A2(n_1557),
.B1(n_1559),
.B2(n_1565),
.C(n_1591),
.Y(n_1732)
);

CKINVDCx16_ASAP7_75t_R g1733 ( 
.A(n_1686),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1697),
.B(n_1638),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1704),
.B(n_1625),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1698),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1680),
.B(n_1622),
.Y(n_1737)
);

AOI222xp33_ASAP7_75t_L g1738 ( 
.A1(n_1701),
.A2(n_1596),
.B1(n_1608),
.B2(n_1593),
.C1(n_1634),
.C2(n_1637),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1680),
.B(n_1622),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1699),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1701),
.B(n_1515),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1705),
.B(n_1638),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1700),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1682),
.B(n_1626),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1696),
.B(n_1619),
.Y(n_1745)
);

INVxp67_ASAP7_75t_L g1746 ( 
.A(n_1693),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1716),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1712),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1682),
.A2(n_1637),
.B1(n_1601),
.B2(n_1620),
.Y(n_1749)
);

CKINVDCx16_ASAP7_75t_R g1750 ( 
.A(n_1682),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1713),
.B(n_1626),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1683),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1714),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1689),
.B(n_1634),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1688),
.Y(n_1755)
);

CKINVDCx16_ASAP7_75t_R g1756 ( 
.A(n_1713),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1721),
.Y(n_1757)
);

NAND2x1p5_ASAP7_75t_L g1758 ( 
.A(n_1722),
.B(n_1685),
.Y(n_1758)
);

NOR2xp67_ASAP7_75t_SL g1759 ( 
.A(n_1733),
.B(n_1386),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1756),
.B(n_1706),
.Y(n_1760)
);

AOI21xp33_ASAP7_75t_SL g1761 ( 
.A1(n_1750),
.A2(n_1437),
.B(n_1719),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1722),
.B(n_1706),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1734),
.B(n_1717),
.Y(n_1763)
);

O2A1O1Ixp33_ASAP7_75t_SL g1764 ( 
.A1(n_1741),
.A2(n_1690),
.B(n_1683),
.C(n_1707),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1721),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1726),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1720),
.B(n_1690),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1732),
.A2(n_1702),
.B1(n_1498),
.B2(n_1487),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1731),
.B(n_1709),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1738),
.A2(n_1703),
.B1(n_1687),
.B2(n_1708),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1725),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1724),
.B(n_1746),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1755),
.B(n_1386),
.Y(n_1773)
);

AO21x1_ASAP7_75t_L g1774 ( 
.A1(n_1720),
.A2(n_1718),
.B(n_1715),
.Y(n_1774)
);

NAND2x1p5_ASAP7_75t_L g1775 ( 
.A(n_1723),
.B(n_1541),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1731),
.B(n_1692),
.Y(n_1776)
);

NOR3xp33_ASAP7_75t_L g1777 ( 
.A(n_1735),
.B(n_1410),
.C(n_1695),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1749),
.A2(n_1637),
.B1(n_1692),
.B2(n_1606),
.Y(n_1778)
);

OAI21xp33_ASAP7_75t_L g1779 ( 
.A1(n_1740),
.A2(n_1681),
.B(n_1333),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1725),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1740),
.B(n_1626),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1727),
.B(n_1628),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1766),
.B(n_1760),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1761),
.B(n_1723),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1767),
.B(n_1726),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1762),
.B(n_1772),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1767),
.Y(n_1787)
);

NAND2x1_ASAP7_75t_L g1788 ( 
.A(n_1759),
.B(n_1723),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1777),
.A2(n_1744),
.B1(n_1728),
.B2(n_1745),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1758),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1757),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1765),
.Y(n_1792)
);

NAND2x1_ASAP7_75t_L g1793 ( 
.A(n_1771),
.B(n_1744),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1780),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1775),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1773),
.B(n_1768),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1776),
.B(n_1728),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1774),
.B(n_1752),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1779),
.B(n_1737),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1779),
.B(n_1737),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1768),
.B(n_1770),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1764),
.B(n_1730),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1769),
.Y(n_1803)
);

AOI222xp33_ASAP7_75t_SL g1804 ( 
.A1(n_1787),
.A2(n_1778),
.B1(n_1748),
.B2(n_1727),
.C1(n_1736),
.C2(n_1753),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1801),
.A2(n_1763),
.B1(n_1778),
.B2(n_1742),
.Y(n_1805)
);

NAND4xp25_ASAP7_75t_SL g1806 ( 
.A(n_1798),
.B(n_1782),
.C(n_1781),
.D(n_1739),
.Y(n_1806)
);

NOR3xp33_ASAP7_75t_L g1807 ( 
.A(n_1788),
.B(n_1736),
.C(n_1729),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1798),
.A2(n_1788),
.B(n_1802),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1796),
.A2(n_1743),
.B(n_1729),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1793),
.A2(n_1747),
.B(n_1743),
.Y(n_1810)
);

OAI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1784),
.A2(n_1747),
.B1(n_1748),
.B2(n_1753),
.C(n_1745),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1790),
.A2(n_1793),
.B1(n_1783),
.B2(n_1786),
.Y(n_1812)
);

NOR3xp33_ASAP7_75t_L g1813 ( 
.A(n_1803),
.B(n_1754),
.C(n_1419),
.Y(n_1813)
);

OAI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1789),
.A2(n_1739),
.B1(n_1751),
.B2(n_1681),
.C(n_1619),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1803),
.B(n_1350),
.Y(n_1815)
);

NAND4xp25_ASAP7_75t_L g1816 ( 
.A(n_1808),
.B(n_1785),
.C(n_1799),
.D(n_1800),
.Y(n_1816)
);

NAND4xp75_ASAP7_75t_SL g1817 ( 
.A(n_1815),
.B(n_1800),
.C(n_1799),
.D(n_1785),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1812),
.B(n_1797),
.Y(n_1818)
);

NOR2xp67_ASAP7_75t_SL g1819 ( 
.A(n_1811),
.B(n_1361),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1805),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1807),
.B(n_1797),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_SL g1822 ( 
.A(n_1806),
.B(n_1404),
.Y(n_1822)
);

NOR3x1_ASAP7_75t_L g1823 ( 
.A(n_1814),
.B(n_1792),
.C(n_1791),
.Y(n_1823)
);

NOR2xp67_ASAP7_75t_L g1824 ( 
.A(n_1810),
.B(n_1795),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1816),
.B(n_1813),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1820),
.A2(n_1809),
.B1(n_1795),
.B2(n_1794),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1822),
.B(n_1751),
.Y(n_1827)
);

AOI211x1_ASAP7_75t_L g1828 ( 
.A1(n_1819),
.A2(n_1804),
.B(n_1656),
.C(n_1655),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1821),
.B(n_1384),
.Y(n_1829)
);

NAND3x1_ASAP7_75t_L g1830 ( 
.A(n_1825),
.B(n_1818),
.C(n_1817),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1826),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1828),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1829),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1827),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1829),
.B(n_1823),
.Y(n_1835)
);

XNOR2xp5_ASAP7_75t_L g1836 ( 
.A(n_1830),
.B(n_1824),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_R g1837 ( 
.A(n_1831),
.B(n_1419),
.Y(n_1837)
);

NAND4xp25_ASAP7_75t_L g1838 ( 
.A(n_1834),
.B(n_1413),
.C(n_1405),
.D(n_1637),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1831),
.Y(n_1839)
);

BUFx6f_ASAP7_75t_L g1840 ( 
.A(n_1833),
.Y(n_1840)
);

XNOR2xp5_ASAP7_75t_L g1841 ( 
.A(n_1836),
.B(n_1835),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1839),
.Y(n_1842)
);

XOR2x2_ASAP7_75t_L g1843 ( 
.A(n_1837),
.B(n_1832),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1843),
.Y(n_1844)
);

NAND2x1_ASAP7_75t_L g1845 ( 
.A(n_1844),
.B(n_1842),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1845),
.A2(n_1840),
.B1(n_1841),
.B2(n_1838),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1845),
.Y(n_1847)
);

OA21x2_ASAP7_75t_L g1848 ( 
.A1(n_1846),
.A2(n_1644),
.B(n_1614),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1847),
.B(n_1620),
.Y(n_1849)
);

XNOR2xp5_ASAP7_75t_L g1850 ( 
.A(n_1849),
.B(n_1848),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1849),
.A2(n_1606),
.B1(n_1616),
.B2(n_1614),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1850),
.A2(n_1431),
.B(n_1405),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1852),
.Y(n_1853)
);

OAI221xp5_ASAP7_75t_R g1854 ( 
.A1(n_1853),
.A2(n_1851),
.B1(n_1431),
.B2(n_1606),
.C(n_1614),
.Y(n_1854)
);

AOI211xp5_ASAP7_75t_L g1855 ( 
.A1(n_1854),
.A2(n_1513),
.B(n_1611),
.C(n_1616),
.Y(n_1855)
);


endmodule