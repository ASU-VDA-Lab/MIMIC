module fake_jpeg_15397_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_1),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_51),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_49),
.B1(n_47),
.B2(n_50),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_49),
.B1(n_53),
.B2(n_43),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_74),
.B1(n_64),
.B2(n_62),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_3),
.Y(n_90)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_54),
.B1(n_52),
.B2(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_42),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_6),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_8),
.B(n_9),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_86),
.B1(n_67),
.B2(n_65),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_85),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_56),
.B1(n_20),
.B2(n_22),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_67),
.B1(n_6),
.B2(n_7),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_4),
.B(n_5),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_4),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_8),
.C(n_9),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_96),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_97),
.A2(n_83),
.B1(n_87),
.B2(n_85),
.Y(n_106)
);

XNOR2x1_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_5),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_104),
.B1(n_10),
.B2(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_103),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_26),
.B(n_38),
.C(n_37),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_106),
.B(n_104),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_92),
.B1(n_89),
.B2(n_15),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_109),
.A2(n_97),
.B1(n_101),
.B2(n_98),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_99),
.B(n_107),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_102),
.B(n_14),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_11),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_118),
.A2(n_108),
.B(n_17),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_121),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_106),
.C(n_23),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_117),
.B1(n_116),
.B2(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_16),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_39),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_27),
.B(n_28),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_29),
.C(n_30),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_33),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_34),
.Y(n_130)
);


endmodule