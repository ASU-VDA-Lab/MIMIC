module fake_ariane_307_n_288 (n_8, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_288);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_288;

wire n_83;
wire n_233;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_195;
wire n_213;
wire n_110;
wire n_197;
wire n_221;
wire n_153;
wire n_86;
wire n_269;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_237;
wire n_172;
wire n_69;
wire n_259;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_242;
wire n_260;
wire n_274;
wire n_115;
wire n_272;
wire n_133;
wire n_66;
wire n_205;
wire n_236;
wire n_265;
wire n_71;
wire n_267;
wire n_208;
wire n_109;
wire n_245;
wire n_96;
wire n_156;
wire n_281;
wire n_209;
wire n_262;
wire n_286;
wire n_174;
wire n_275;
wire n_100;
wire n_283;
wire n_187;
wire n_132;
wire n_62;
wire n_210;
wire n_147;
wire n_204;
wire n_225;
wire n_235;
wire n_200;
wire n_166;
wire n_253;
wire n_76;
wire n_218;
wire n_103;
wire n_79;
wire n_246;
wire n_226;
wire n_244;
wire n_271;
wire n_220;
wire n_84;
wire n_247;
wire n_261;
wire n_199;
wire n_159;
wire n_189;
wire n_107;
wire n_91;
wire n_72;
wire n_128;
wire n_105;
wire n_217;
wire n_240;
wire n_82;
wire n_178;
wire n_224;
wire n_57;
wire n_131;
wire n_263;
wire n_201;
wire n_229;
wire n_70;
wire n_250;
wire n_222;
wire n_117;
wire n_139;
wire n_165;
wire n_287;
wire n_85;
wire n_144;
wire n_130;
wire n_256;
wire n_214;
wire n_227;
wire n_101;
wire n_94;
wire n_243;
wire n_284;
wire n_134;
wire n_188;
wire n_185;
wire n_249;
wire n_58;
wire n_65;
wire n_123;
wire n_212;
wire n_138;
wire n_112;
wire n_162;
wire n_264;
wire n_129;
wire n_126;
wire n_137;
wire n_255;
wire n_278;
wire n_122;
wire n_268;
wire n_257;
wire n_266;
wire n_198;
wire n_282;
wire n_148;
wire n_232;
wire n_164;
wire n_52;
wire n_277;
wire n_157;
wire n_248;
wire n_184;
wire n_177;
wire n_135;
wire n_258;
wire n_73;
wire n_77;
wire n_171;
wire n_228;
wire n_121;
wire n_118;
wire n_93;
wire n_276;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_81;
wire n_87;
wire n_206;
wire n_279;
wire n_207;
wire n_241;
wire n_254;
wire n_238;
wire n_219;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_231;
wire n_192;
wire n_80;
wire n_146;
wire n_234;
wire n_230;
wire n_211;
wire n_270;
wire n_194;
wire n_97;
wire n_154;
wire n_280;
wire n_215;
wire n_252;
wire n_142;
wire n_251;
wire n_161;
wire n_285;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_78;
wire n_193;
wire n_63;
wire n_59;
wire n_99;
wire n_216;
wire n_155;
wire n_127;
wire n_239;
wire n_223;
wire n_273;
wire n_54;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

INVxp67_ASAP7_75t_SL g60 ( 
.A(n_10),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_27),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_1),
.Y(n_90)
);

OA21x2_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_1),
.B(n_2),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_3),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_4),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_4),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_55),
.A2(n_5),
.B1(n_6),
.B2(n_50),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_5),
.Y(n_106)
);

NAND2x1p5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_8),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_9),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_59),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_65),
.A2(n_68),
.B1(n_60),
.B2(n_81),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_83),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_82),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_76),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_68),
.B1(n_65),
.B2(n_60),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_77),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_52),
.B1(n_18),
.B2(n_20),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_16),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_26),
.Y(n_129)
);

AND2x6_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_28),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_86),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

NAND3x1_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_29),
.C(n_31),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_88),
.B(n_32),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_113),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_100),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_115),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_84),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_107),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_107),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_121),
.B(n_105),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_94),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_129),
.B(n_124),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_84),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

AND2x4_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_140),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_141),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_116),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_123),
.B(n_94),
.C(n_93),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

AND2x4_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_125),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_104),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_149),
.Y(n_171)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_99),
.Y(n_172)
);

AND2x4_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_108),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

CKINVDCx6p67_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_149),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_152),
.B(n_150),
.C(n_137),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_167),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

AO21x2_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_155),
.B(n_142),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_173),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_149),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_149),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_176),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_180),
.A2(n_161),
.B(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_178),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_173),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

OAI31xp33_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_169),
.A3(n_171),
.B(n_180),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_189),
.B(n_186),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_169),
.Y(n_220)
);

OAI322xp33_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_166),
.A3(n_170),
.B1(n_143),
.B2(n_145),
.C1(n_136),
.C2(n_163),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

OAI31xp33_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_170),
.A3(n_172),
.B(n_173),
.Y(n_224)
);

OAI211xp5_ASAP7_75t_SL g225 ( 
.A1(n_205),
.A2(n_162),
.B(n_158),
.C(n_174),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_160),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_163),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_200),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_91),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_178),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

AOI211xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_109),
.B(n_161),
.C(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_209),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_227),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_216),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_219),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_240),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_215),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_215),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_211),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_216),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_135),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_229),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_130),
.Y(n_259)
);

OAI33xp33_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_225),
.A3(n_142),
.B1(n_151),
.B2(n_194),
.B3(n_203),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

AOI211xp5_ASAP7_75t_L g263 ( 
.A1(n_259),
.A2(n_249),
.B(n_253),
.C(n_247),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_256),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_247),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_245),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_254),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_265),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_260),
.B(n_257),
.Y(n_269)
);

AND3x4_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_255),
.C(n_161),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_266),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_245),
.B1(n_251),
.B2(n_262),
.Y(n_274)
);

XOR2x2_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_235),
.Y(n_275)
);

NOR4xp25_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_193),
.C(n_158),
.D(n_174),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_275),
.B(n_224),
.Y(n_277)
);

NOR3xp33_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_188),
.C(n_174),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_277),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_35),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_277),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_281),
.Y(n_283)
);

AOI221xp5_ASAP7_75t_L g284 ( 
.A1(n_279),
.A2(n_190),
.B1(n_223),
.B2(n_153),
.C(n_151),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_190),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_209),
.B(n_186),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_283),
.Y(n_287)
);

AOI221xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.C(n_189),
.Y(n_288)
);


endmodule