module fake_jpeg_985_n_348 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_49),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_50),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_76),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_59),
.Y(n_114)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_62),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_6),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_21),
.B(n_6),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_80),
.Y(n_126)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_19),
.B(n_7),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_74),
.B(n_92),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_34),
.Y(n_75)
);

NAND2x1_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_24),
.B(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_85),
.Y(n_111)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_23),
.B(n_8),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_23),
.B(n_8),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_87),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_26),
.B(n_32),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_94),
.Y(n_121)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_46),
.Y(n_117)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_45),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_75),
.A2(n_48),
.B1(n_47),
.B2(n_32),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_99),
.A2(n_113),
.B1(n_122),
.B2(n_124),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_47),
.B1(n_26),
.B2(n_35),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_55),
.A2(n_38),
.B1(n_37),
.B2(n_35),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_62),
.A2(n_38),
.B1(n_37),
.B2(n_40),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_51),
.A2(n_46),
.B1(n_45),
.B2(n_40),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_141),
.B1(n_142),
.B2(n_151),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_126),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_137),
.B1(n_147),
.B2(n_141),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_10),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_132),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_72),
.B(n_10),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_13),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_143),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_74),
.A2(n_22),
.B1(n_28),
.B2(n_30),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_52),
.A2(n_28),
.B1(n_30),
.B2(n_16),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_93),
.A2(n_28),
.B1(n_30),
.B2(n_16),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_14),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_54),
.B(n_14),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_146),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_15),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_56),
.A2(n_28),
.B1(n_30),
.B2(n_15),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_63),
.A2(n_28),
.B1(n_30),
.B2(n_68),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_161),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_102),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_181),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_111),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_159),
.B(n_165),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_104),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_182),
.Y(n_201)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_124),
.A2(n_70),
.B1(n_79),
.B2(n_59),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_164),
.A2(n_190),
.B1(n_157),
.B2(n_163),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_104),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_100),
.A2(n_142),
.B(n_119),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_166),
.A2(n_171),
.B(n_155),
.Y(n_214)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_169),
.B(n_186),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_116),
.A2(n_133),
.B1(n_119),
.B2(n_136),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_183),
.B1(n_194),
.B2(n_189),
.Y(n_210)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_105),
.A2(n_118),
.B1(n_110),
.B2(n_139),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_180),
.A2(n_193),
.B1(n_196),
.B2(n_175),
.Y(n_209)
);

NAND2x1_ASAP7_75t_L g181 ( 
.A(n_98),
.B(n_110),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_97),
.B(n_127),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g183 ( 
.A1(n_99),
.A2(n_113),
.B1(n_122),
.B2(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_149),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_181),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_115),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_140),
.B(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_189),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_149),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_120),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_106),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_197),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_134),
.A2(n_130),
.B1(n_138),
.B2(n_120),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_107),
.A2(n_108),
.B1(n_138),
.B2(n_130),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_137),
.A2(n_50),
.B1(n_75),
.B2(n_88),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

AO21x2_ASAP7_75t_L g199 ( 
.A1(n_160),
.A2(n_181),
.B(n_185),
.Y(n_199)
);

OA22x2_ASAP7_75t_L g249 ( 
.A1(n_199),
.A2(n_203),
.B1(n_209),
.B2(n_216),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g200 ( 
.A(n_182),
.B(n_152),
.C(n_155),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_206),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_156),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_204),
.B(n_214),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_171),
.B1(n_169),
.B2(n_188),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_207),
.A2(n_210),
.B1(n_212),
.B2(n_216),
.Y(n_250)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_169),
.A2(n_166),
.B1(n_153),
.B2(n_183),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_153),
.A2(n_168),
.B1(n_172),
.B2(n_191),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_153),
.B(n_170),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_174),
.C(n_179),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_158),
.B(n_176),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_227),
.Y(n_229)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_211),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_242),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_217),
.B(n_153),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_233),
.B(n_240),
.Y(n_258)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_195),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_235),
.B(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_211),
.Y(n_237)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_214),
.B(n_173),
.CI(n_184),
.CON(n_239),
.SN(n_239)
);

AOI221xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.C(n_256),
.Y(n_261)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_167),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_199),
.A2(n_178),
.B1(n_210),
.B2(n_207),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_199),
.B1(n_205),
.B2(n_203),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_247),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_212),
.C(n_206),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_249),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_208),
.B(n_228),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_201),
.A2(n_198),
.B(n_202),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_228),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_253),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_225),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_254),
.Y(n_262)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_202),
.B(n_201),
.C(n_205),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_199),
.B1(n_247),
.B2(n_238),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_248),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_270),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_254),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_231),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_246),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_244),
.A2(n_205),
.B1(n_204),
.B2(n_223),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_277),
.A2(n_205),
.B1(n_249),
.B2(n_239),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_232),
.B1(n_245),
.B2(n_250),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_279),
.A2(n_281),
.B1(n_290),
.B2(n_199),
.Y(n_303)
);

XOR2x2_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_230),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_295),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_233),
.C(n_240),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_286),
.C(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_264),
.B(n_255),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_292),
.Y(n_298)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_256),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_230),
.C(n_252),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_266),
.A2(n_244),
.B(n_249),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_289),
.A2(n_270),
.B(n_199),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_249),
.C(n_236),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_257),
.C(n_262),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_215),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

XOR2x2_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_239),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_267),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_274),
.C(n_265),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_304),
.C(n_295),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_294),
.B1(n_293),
.B2(n_276),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_288),
.C(n_280),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_307),
.Y(n_311)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_289),
.B(n_281),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_319),
.C(n_296),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_291),
.B(n_278),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_312),
.A2(n_314),
.B(n_306),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_313),
.A2(n_260),
.B(n_259),
.C(n_272),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_297),
.B(n_275),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_316),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_263),
.Y(n_318)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_318),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_272),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_268),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_287),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_322),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_304),
.C(n_302),
.Y(n_322)
);

AOI21x1_ASAP7_75t_L g333 ( 
.A1(n_323),
.A2(n_313),
.B(n_315),
.Y(n_333)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_324),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_300),
.C(n_268),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_328),
.B1(n_311),
.B2(n_317),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_309),
.C(n_267),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_329),
.A2(n_260),
.B(n_259),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_330),
.B(n_335),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_332),
.A2(n_333),
.B(n_329),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_314),
.B1(n_299),
.B2(n_200),
.Y(n_335)
);

AO21x1_ASAP7_75t_L g343 ( 
.A1(n_336),
.A2(n_337),
.B(n_338),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_334),
.B(n_322),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_332),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_327),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_340),
.A2(n_243),
.B(n_224),
.Y(n_342)
);

O2A1O1Ixp33_ASAP7_75t_SL g341 ( 
.A1(n_336),
.A2(n_200),
.B(n_334),
.C(n_299),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_341),
.B(n_342),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_339),
.C(n_221),
.Y(n_344)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_344),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_345),
.C(n_234),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_241),
.Y(n_348)
);


endmodule