module fake_jpeg_8999_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx6p67_ASAP7_75t_R g80 ( 
.A(n_36),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_25),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_22),
.B1(n_30),
.B2(n_29),
.Y(n_66)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_45),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_49),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_51),
.B(n_53),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_63),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_78),
.B1(n_16),
.B2(n_27),
.Y(n_98)
);

NAND2x1_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_23),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_66),
.B(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_26),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_13),
.C(n_15),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_18),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_23),
.B1(n_21),
.B2(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_21),
.B1(n_34),
.B2(n_30),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_87),
.B(n_115),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_85),
.A2(n_10),
.B(n_14),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_34),
.B1(n_30),
.B2(n_29),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_94),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_15),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_54),
.A2(n_29),
.B1(n_31),
.B2(n_26),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_93),
.A2(n_95),
.B1(n_32),
.B2(n_61),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_52),
.A2(n_31),
.B1(n_16),
.B2(n_27),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_55),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_105),
.B(n_107),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_70),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_108),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_114),
.Y(n_121)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_74),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_61),
.A2(n_16),
.B1(n_28),
.B2(n_19),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_61),
.A2(n_28),
.B1(n_19),
.B2(n_32),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_58),
.B(n_56),
.Y(n_143)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_74),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_53),
.Y(n_123)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_120),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_123),
.B(n_130),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_142),
.Y(n_154)
);

AOI32xp33_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_65),
.A3(n_73),
.B1(n_72),
.B2(n_63),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_86),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_134),
.B(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_86),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_141),
.B(n_148),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_66),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_143),
.A2(n_109),
.B(n_67),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_77),
.B1(n_71),
.B2(n_65),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_149),
.B1(n_99),
.B2(n_103),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_88),
.B(n_60),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_89),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_151),
.B(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_77),
.B1(n_71),
.B2(n_72),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_110),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_0),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_152),
.B(n_150),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_159),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_SL g197 ( 
.A(n_155),
.B(n_156),
.C(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_160),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_166),
.B(n_143),
.Y(n_189)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_104),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_101),
.B1(n_100),
.B2(n_105),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_86),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_169),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_102),
.B(n_94),
.C(n_120),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_163),
.A2(n_138),
.B(n_122),
.Y(n_205)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_177),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_90),
.B1(n_71),
.B2(n_69),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_168),
.B1(n_182),
.B2(n_144),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_118),
.B1(n_81),
.B2(n_102),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_106),
.B1(n_73),
.B2(n_117),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_81),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_170),
.B(n_171),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_118),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_172),
.B(n_175),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_10),
.B(n_12),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_124),
.A2(n_106),
.B1(n_113),
.B2(n_108),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_127),
.B1(n_123),
.B2(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_82),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_122),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_179),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_171),
.B(n_151),
.Y(n_208)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_183),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_135),
.A2(n_111),
.B1(n_96),
.B2(n_109),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_96),
.C(n_1),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_184),
.B(n_149),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_186),
.B(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_189),
.A2(n_199),
.B(n_203),
.Y(n_234)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_200),
.B1(n_201),
.B2(n_214),
.Y(n_225)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_175),
.Y(n_221)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_209),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_124),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_156),
.A2(n_121),
.B1(n_147),
.B2(n_145),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_8),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_151),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_205),
.B(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_153),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_151),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_137),
.B(n_130),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_172),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_216),
.Y(n_245)
);

OA22x2_ASAP7_75t_SL g213 ( 
.A1(n_162),
.A2(n_154),
.B1(n_155),
.B2(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_154),
.A2(n_138),
.B1(n_134),
.B2(n_137),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_169),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_167),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_130),
.C(n_10),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_203),
.A2(n_178),
.B1(n_165),
.B2(n_160),
.Y(n_219)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_221),
.A2(n_222),
.B(n_226),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_187),
.A2(n_157),
.B1(n_158),
.B2(n_184),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_164),
.Y(n_224)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_144),
.C(n_159),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_233),
.C(n_202),
.Y(n_252)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_229),
.B(n_238),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_186),
.Y(n_250)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_242),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_144),
.C(n_183),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_129),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_237),
.B1(n_243),
.B2(n_218),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_0),
.Y(n_236)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_240),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_217),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_201),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_228),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_246),
.B(n_248),
.Y(n_279)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_261),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_267),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_253),
.C(n_254),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_244),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_197),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_209),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_197),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_260),
.C(n_234),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_208),
.C(n_189),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_196),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_263),
.A2(n_243),
.B1(n_237),
.B2(n_240),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_216),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_221),
.Y(n_272)
);

NAND2x1_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_241),
.Y(n_267)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_257),
.A2(n_191),
.B1(n_214),
.B2(n_219),
.Y(n_269)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_191),
.B1(n_222),
.B2(n_223),
.Y(n_271)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_277),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_233),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_223),
.C(n_226),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_282),
.C(n_285),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_255),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_194),
.B1(n_220),
.B2(n_212),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_281),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_200),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_199),
.B1(n_212),
.B2(n_232),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_266),
.B1(n_262),
.B2(n_248),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_199),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_265),
.B(n_205),
.Y(n_286)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_292),
.B(n_300),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_260),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_270),
.C(n_273),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_291),
.A2(n_293),
.B1(n_282),
.B2(n_272),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_265),
.B(n_255),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_276),
.A2(n_253),
.B1(n_264),
.B2(n_249),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_204),
.B(n_210),
.Y(n_297)
);

AOI221xp5_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_274),
.B1(n_204),
.B2(n_210),
.C(n_285),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_279),
.A2(n_207),
.B(n_247),
.Y(n_300)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_305),
.C(n_306),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_270),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_292),
.C(n_290),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_312),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_273),
.C(n_275),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_309),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_289),
.A2(n_236),
.B1(n_207),
.B2(n_192),
.Y(n_309)
);

AO221x1_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_3),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_4),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_4),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_298),
.B(n_294),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_314),
.A2(n_320),
.B(n_5),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_7),
.Y(n_325)
);

AOI211xp5_ASAP7_75t_L g318 ( 
.A1(n_302),
.A2(n_299),
.B(n_287),
.C(n_286),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_293),
.A3(n_306),
.B1(n_308),
.B2(n_304),
.C1(n_305),
.C2(n_7),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_307),
.A2(n_297),
.B(n_287),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_312),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_322),
.B(n_326),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_313),
.A2(n_316),
.B(n_320),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_319),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_326),
.B(n_327),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_331),
.A2(n_332),
.B(n_330),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_319),
.B(n_315),
.Y(n_332)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_6),
.B(n_332),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_6),
.Y(n_336)
);


endmodule