module real_jpeg_18870_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_2),
.B(n_133),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_2),
.B(n_289),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_2),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_2),
.B(n_438),
.Y(n_437)
);

NAND2xp33_ASAP7_75t_SL g475 ( 
.A(n_2),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_2),
.B(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_2),
.B(n_508),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_3),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_3),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_3),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_3),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_3),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_3),
.B(n_136),
.Y(n_135)
);

NAND2x1p5_ASAP7_75t_L g223 ( 
.A(n_3),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_4),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g479 ( 
.A(n_4),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_5),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_5),
.Y(n_350)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_5),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_6),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_6),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_6),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_6),
.B(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_6),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_6),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_6),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_6),
.B(n_217),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_7),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g296 ( 
.A(n_7),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_7),
.Y(n_462)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_8),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_8),
.Y(n_353)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_8),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_9),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_9),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_9),
.B(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_9),
.B(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g299 ( 
.A(n_9),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_9),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_9),
.B(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_9),
.B(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_10),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_10),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_10),
.B(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_10),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_10),
.B(n_433),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_10),
.B(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_10),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_10),
.B(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_11),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_11),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g215 ( 
.A(n_11),
.Y(n_215)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_12),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_12),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_12),
.B(n_56),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_12),
.A2(n_17),
.B1(n_310),
.B2(n_314),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_12),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_12),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_12),
.B(n_494),
.Y(n_493)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_13),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_13),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_13),
.Y(n_291)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_14),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_14),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_14),
.B(n_274),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_14),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_14),
.B(n_296),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_15),
.Y(n_111)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g213 ( 
.A(n_16),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_16),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_16),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_17),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_17),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_17),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_17),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_17),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_17),
.B(n_132),
.Y(n_237)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_17),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

A2O1A1O1Ixp25_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_257),
.B(n_530),
.C(n_537),
.D(n_539),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_227),
.C(n_245),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_180),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21x1_ASAP7_75t_SL g532 ( 
.A1(n_26),
.A2(n_533),
.B(n_534),
.Y(n_532)
);

NOR2xp67_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_148),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_27),
.B(n_148),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_112),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_28),
.B(n_113),
.C(n_125),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_78),
.C(n_94),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_29),
.B(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_48),
.C(n_63),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_30),
.B(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_41),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_32),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_32),
.A2(n_39),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_32),
.B(n_40),
.C(n_41),
.Y(n_124)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_32),
.B(n_298),
.C(n_299),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_32),
.A2(n_39),
.B1(n_298),
.B2(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_34),
.Y(n_445)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_35),
.B(n_97),
.C(n_100),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_35),
.A2(n_40),
.B1(n_97),
.B2(n_98),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_35),
.B(n_216),
.Y(n_328)
);

XNOR2x1_ASAP7_75t_SL g409 ( 
.A(n_35),
.B(n_307),
.Y(n_409)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_37),
.Y(n_164)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_37),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_38),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_39),
.B(n_116),
.C(n_119),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_42),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_42),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_47),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_47),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_48),
.B(n_63),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.C(n_58),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_49),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_166)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_58),
.A2(n_59),
.B1(n_116),
.B2(n_118),
.Y(n_319)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_59),
.B(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_59),
.B(n_116),
.C(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_62),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_64),
.B(n_72),
.C(n_76),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_64),
.B(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_64),
.B(n_139),
.C(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_72),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_72),
.A2(n_77),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_77),
.B(n_139),
.C(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_78),
.B(n_94),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_88),
.B2(n_93),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_83),
.C(n_88),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_82),
.B(n_169),
.C(n_172),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_82),
.B(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_87),
.Y(n_316)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_88),
.A2(n_93),
.B1(n_251),
.B2(n_254),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_L g538 ( 
.A(n_88),
.B(n_252),
.C(n_253),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_92),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.C(n_108),
.Y(n_94)
);

AO22x1_ASAP7_75t_SL g177 ( 
.A1(n_95),
.A2(n_96),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_159),
.C(n_162),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_97),
.A2(n_98),
.B1(n_162),
.B2(n_163),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_97),
.B(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_98),
.B(n_417),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_99),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_100),
.B(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_100),
.A2(n_249),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_100),
.Y(n_252)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_104),
.A2(n_248),
.B(n_538),
.Y(n_539)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_105),
.B(n_108),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_108),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_108),
.A2(n_144),
.B1(n_174),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_111),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_125),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_123),
.C(n_124),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_118),
.B1(n_135),
.B2(n_139),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_118),
.B(n_135),
.C(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_124),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_140),
.B2(n_141),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_128),
.B(n_129),
.C(n_140),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_130),
.Y(n_239)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_135),
.A2(n_139),
.B1(n_222),
.B2(n_223),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_135),
.A2(n_139),
.B1(n_196),
.B2(n_267),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_136),
.Y(n_282)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_142),
.B(n_144),
.C(n_146),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_168),
.C(n_174),
.Y(n_167)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_151),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_167),
.C(n_177),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_155),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_165),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_156),
.B(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_158),
.B(n_165),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_160),
.B(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_160),
.B(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_162),
.A2(n_163),
.B1(n_294),
.B2(n_295),
.Y(n_345)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_163),
.B(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_167),
.B(n_177),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_194),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_171),
.Y(n_300)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

OR2x2_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_181),
.B(n_183),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_190),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_184),
.B(n_188),
.Y(n_394)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_190),
.B(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_203),
.C(n_207),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_191),
.A2(n_192),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.C(n_200),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g379 ( 
.A(n_193),
.B(n_380),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_195),
.B(n_201),
.Y(n_380)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_196),
.Y(n_267)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_219),
.C(n_222),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_209),
.A2(n_210),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.C(n_216),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_211),
.A2(n_216),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_211),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_214),
.B(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_216),
.Y(n_307)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_218),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_221),
.Y(n_275)
);

BUFx2_ASAP7_75t_R g249 ( 
.A(n_222),
.Y(n_249)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

A2O1A1O1Ixp25_ASAP7_75t_L g531 ( 
.A1(n_228),
.A2(n_246),
.B(n_532),
.C(n_535),
.D(n_536),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_244),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_229),
.B(n_244),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_232),
.C(n_243),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_242),
.B2(n_243),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_238),
.C(n_240),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_256),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_247),
.B(n_256),
.Y(n_536)
);

BUFx24_ASAP7_75t_SL g540 ( 
.A(n_247),
.Y(n_540)
);

FAx1_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_250),
.CI(n_255),
.CON(n_247),
.SN(n_247)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_251),
.Y(n_254)
);

NAND2x1_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_524),
.Y(n_257)
);

NAND4xp25_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_381),
.C(n_395),
.D(n_400),
.Y(n_258)
);

NOR2x1_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_358),
.Y(n_259)
);

NOR2xp67_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_334),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_261),
.B(n_334),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_301),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_262),
.B(n_302),
.C(n_317),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_279),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_264),
.Y(n_362)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_268),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_277),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_272),
.B1(n_273),
.B2(n_276),
.Y(n_269)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g374 ( 
.A1(n_270),
.A2(n_273),
.B(n_277),
.C(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_272),
.B(n_276),
.Y(n_375)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_275),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_279),
.B(n_362),
.C(n_363),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_292),
.C(n_297),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_280),
.B(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_284),
.C(n_288),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_288),
.Y(n_283)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_292),
.A2(n_293),
.B1(n_297),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx12f_ASAP7_75t_L g517 ( 
.A(n_296),
.Y(n_517)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_298),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_299),
.B(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_317),
.Y(n_301)
);

XOR2x2_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_309),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_304),
.B(n_368),
.C(n_369),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_308),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_321),
.B(n_323),
.Y(n_320)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_309),
.Y(n_368)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_SL g495 ( 
.A(n_312),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_314),
.Y(n_322)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_316),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.C(n_327),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_320),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_327),
.B(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.C(n_332),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_328),
.B(n_407),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_329),
.A2(n_330),
.B1(n_332),
.B2(n_333),
.Y(n_407)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_337),
.C(n_341),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_335),
.B(n_423),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_337),
.A2(n_338),
.B1(n_341),
.B2(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_341),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_345),
.C(n_346),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_342),
.B(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_345),
.B(n_346),
.Y(n_405)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_351),
.C(n_354),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_347),
.B(n_354),
.Y(n_447)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_351),
.B(n_447),
.Y(n_446)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

OAI21x1_ASAP7_75t_SL g525 ( 
.A1(n_358),
.A2(n_526),
.B(n_527),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_359),
.B(n_360),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_361),
.B(n_365),
.C(n_379),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_365),
.A2(n_366),
.B1(n_378),
.B2(n_379),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_374),
.B1(n_376),
.B2(n_377),
.Y(n_370)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_371),
.Y(n_376)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_374),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_374),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_389),
.C(n_390),
.Y(n_388)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

A2O1A1O1Ixp25_ASAP7_75t_L g524 ( 
.A1(n_381),
.A2(n_395),
.B(n_525),
.C(n_528),
.D(n_529),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_393),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_382),
.B(n_393),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_387),
.C(n_391),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_383),
.A2(n_384),
.B1(n_391),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_385),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_388),
.B(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_391),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_396),
.B(n_397),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_425),
.B(n_523),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_422),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_402),
.B(n_422),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_406),
.C(n_408),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_403),
.A2(n_404),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_406),
.B(n_408),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.C(n_416),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_409),
.A2(n_410),
.B1(n_411),
.B2(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_409),
.Y(n_430)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_416),
.B(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_421),
.Y(n_492)
);

AOI21x1_ASAP7_75t_SL g425 ( 
.A1(n_426),
.A2(n_451),
.B(n_522),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_448),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_427),
.B(n_448),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_431),
.C(n_446),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_428),
.B(n_469),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_446),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_437),
.C(n_443),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_456),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_436),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_443),
.Y(n_456)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_470),
.B(n_521),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_468),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_453),
.B(n_468),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_457),
.C(n_466),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_454),
.A2(n_455),
.B1(n_481),
.B2(n_483),
.Y(n_480)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_457),
.A2(n_466),
.B1(n_467),
.B2(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_457),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_463),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_458),
.A2(n_459),
.B1(n_463),
.B2(n_464),
.Y(n_473)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_484),
.B(n_520),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_480),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_472),
.B(n_480),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.C(n_478),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_473),
.B(n_497),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_474),
.A2(n_475),
.B1(n_478),
.B2(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_478),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_481),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_485),
.A2(n_499),
.B(n_519),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_496),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_486),
.B(n_496),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_493),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_487),
.B(n_493),
.Y(n_505)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_506),
.B(n_518),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_505),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_501),
.B(n_505),
.Y(n_518)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_514),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx6_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_538),
.Y(n_537)
);


endmodule