module fake_jpeg_23168_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_41),
.B(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_48),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_55),
.Y(n_100)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_39),
.Y(n_56)
);

OR2x4_ASAP7_75t_L g129 ( 
.A(n_56),
.B(n_29),
.Y(n_129)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_63),
.Y(n_104)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_17),
.B1(n_32),
.B2(n_30),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_60),
.A2(n_73),
.B(n_85),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_30),
.B1(n_17),
.B2(n_32),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_61),
.A2(n_70),
.B1(n_92),
.B2(n_29),
.Y(n_121)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_66),
.Y(n_113)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_72),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_17),
.B1(n_32),
.B2(n_20),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_71),
.Y(n_102)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_38),
.B1(n_39),
.B2(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_76),
.Y(n_124)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_86),
.Y(n_125)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_19),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_26),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_38),
.B1(n_39),
.B2(n_37),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_40),
.B(n_25),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_90),
.B(n_35),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_37),
.B1(n_34),
.B2(n_23),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_95),
.B(n_97),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_35),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_98),
.B(n_99),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_23),
.A3(n_31),
.B1(n_27),
.B2(n_24),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_23),
.C(n_33),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_107),
.B(n_109),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_81),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_56),
.A2(n_18),
.B(n_26),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_33),
.B(n_31),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_29),
.B(n_18),
.C(n_23),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_117),
.B(n_119),
.Y(n_163)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_85),
.B(n_13),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_121),
.B1(n_27),
.B2(n_24),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_65),
.B(n_13),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

AND2x4_ASAP7_75t_SL g128 ( 
.A(n_68),
.B(n_22),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_54),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_68),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_103),
.B1(n_121),
.B2(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_134),
.B1(n_139),
.B2(n_148),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_60),
.B(n_78),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_132),
.A2(n_137),
.B(n_145),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_91),
.B1(n_57),
.B2(n_62),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_133),
.A2(n_138),
.B1(n_146),
.B2(n_112),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_136),
.A2(n_113),
.B(n_115),
.C(n_102),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_91),
.B1(n_93),
.B2(n_77),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_22),
.B1(n_33),
.B2(n_31),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_71),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_160),
.Y(n_177)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_144),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_108),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_0),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_105),
.B1(n_118),
.B2(n_101),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_147),
.B(n_100),
.Y(n_166)
);

AOI22x1_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_22),
.B1(n_27),
.B2(n_24),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_108),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_107),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_151),
.B1(n_106),
.B2(n_127),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_110),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_161),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_0),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_114),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_167),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_166),
.A2(n_186),
.B(n_197),
.Y(n_225)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_157),
.B(n_98),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_168),
.B(n_172),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_147),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_188),
.B1(n_195),
.B2(n_139),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_112),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_173),
.B(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_178),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_127),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_180),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_126),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_183),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_126),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_146),
.A2(n_123),
.B1(n_94),
.B2(n_106),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_184),
.A2(n_199),
.B1(n_6),
.B2(n_8),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_162),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_132),
.A2(n_123),
.B1(n_96),
.B2(n_115),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_189),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_190),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_114),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_151),
.B(n_140),
.C(n_143),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_96),
.Y(n_193)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_131),
.A2(n_102),
.B1(n_1),
.B2(n_2),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_160),
.B(n_8),
.Y(n_196)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_8),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_134),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_199)
);

NOR2x1p5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_148),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g249 ( 
.A1(n_201),
.A2(n_226),
.B1(n_11),
.B2(n_12),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_223),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_219),
.C(n_179),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_163),
.B1(n_153),
.B2(n_137),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_211),
.B1(n_217),
.B2(n_218),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_137),
.B1(n_149),
.B2(n_133),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_177),
.B(n_138),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_227),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_184),
.A2(n_183),
.B1(n_166),
.B2(n_175),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_173),
.C(n_177),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_1),
.B(n_3),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_199),
.Y(n_238)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_175),
.A2(n_135),
.B1(n_144),
.B2(n_130),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_9),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_180),
.Y(n_229)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_200),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_231),
.B(n_238),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_236),
.Y(n_269)
);

AOI211xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_191),
.B(n_195),
.C(n_186),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_234),
.B(n_248),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_169),
.Y(n_235)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_206),
.C(n_205),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_182),
.C(n_178),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_244),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_197),
.C(n_171),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_242),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_208),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_241),
.Y(n_255)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_246),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_208),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_192),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_249),
.A2(n_220),
.B1(n_222),
.B2(n_204),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_215),
.C(n_209),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_251),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_181),
.C(n_174),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_218),
.B1(n_201),
.B2(n_203),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_252),
.A2(n_258),
.B1(n_249),
.B2(n_202),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_243),
.A2(n_201),
.B(n_221),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_254),
.A2(n_267),
.B1(n_249),
.B2(n_238),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_213),
.B1(n_207),
.B2(n_227),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_245),
.B(n_228),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_245),
.Y(n_271)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_240),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_236),
.Y(n_272)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_239),
.B1(n_234),
.B2(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_230),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_279),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_233),
.C(n_248),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_269),
.C(n_265),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_256),
.B(n_220),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_283),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_229),
.B1(n_242),
.B2(n_235),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_281),
.Y(n_297)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_280),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_300)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_263),
.B(n_222),
.Y(n_282)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_255),
.B(n_213),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_252),
.A2(n_249),
.B1(n_204),
.B2(n_202),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_167),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_254),
.B(n_265),
.Y(n_288)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_290),
.C(n_295),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_270),
.C(n_257),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_264),
.B(n_259),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_268),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_264),
.C(n_260),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_279),
.B(n_274),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_297),
.B1(n_300),
.B2(n_299),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_306),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_300),
.A2(n_278),
.B1(n_284),
.B2(n_281),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_307),
.B1(n_260),
.B2(n_189),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_290),
.Y(n_316)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_298),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_286),
.B1(n_273),
.B2(n_275),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_266),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_294),
.C(n_287),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_310),
.A2(n_305),
.B1(n_223),
.B2(n_15),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_SL g311 ( 
.A(n_303),
.B(n_289),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_314),
.B(n_302),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_295),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_316),
.Y(n_321)
);

AOI31xp33_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_267),
.A3(n_292),
.B(n_273),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_317),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_309),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_318),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_322),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_313),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_324),
.B(n_322),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_320),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.C(n_325),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_316),
.B1(n_214),
.B2(n_15),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_11),
.C(n_14),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_16),
.B(n_14),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_15),
.Y(n_332)
);


endmodule