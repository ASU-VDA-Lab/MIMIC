module fake_jpeg_28886_n_535 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_535);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_535;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_55),
.Y(n_143)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_6),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_58),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_10),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_66),
.Y(n_166)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_67),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_17),
.B(n_10),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_83),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g125 ( 
.A(n_74),
.Y(n_125)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

HAxp5_ASAP7_75t_SL g76 ( 
.A(n_24),
.B(n_15),
.CON(n_76),
.SN(n_76)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_34),
.Y(n_110)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_17),
.B(n_5),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_33),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_84),
.B(n_89),
.Y(n_169)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_92),
.B(n_94),
.Y(n_171)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_25),
.B(n_5),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_100),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_25),
.B(n_4),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_101),
.B(n_32),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_102),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_104),
.Y(n_163)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_110),
.B(n_29),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_31),
.B1(n_46),
.B2(n_38),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_118),
.A2(n_124),
.B1(n_136),
.B2(n_146),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_31),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_119),
.B(n_39),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_32),
.B1(n_46),
.B2(n_38),
.Y(n_124)
);

BUFx10_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_126),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_135),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_76),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_86),
.A2(n_20),
.B1(n_43),
.B2(n_34),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_107),
.A2(n_34),
.B1(n_40),
.B2(n_20),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_141),
.A2(n_44),
.B1(n_54),
.B2(n_63),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_90),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_59),
.A2(n_20),
.B1(n_43),
.B2(n_29),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_106),
.B1(n_103),
.B2(n_100),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_60),
.B(n_28),
.C(n_47),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_162),
.B(n_44),
.C(n_39),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_109),
.A2(n_43),
.B1(n_48),
.B2(n_52),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_164),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_55),
.B(n_23),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_165),
.B(n_125),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_SL g173 ( 
.A(n_85),
.Y(n_173)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_74),
.Y(n_186)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_176),
.Y(n_230)
);

AOI32xp33_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_111),
.A3(n_110),
.B1(n_122),
.B2(n_169),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_177),
.B(n_186),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_181),
.B(n_194),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_182),
.A2(n_185),
.B1(n_196),
.B2(n_198),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_134),
.B(n_65),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_183),
.B(n_211),
.C(n_214),
.Y(n_260)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_123),
.A2(n_98),
.B1(n_87),
.B2(n_96),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_113),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_190),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_74),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_191),
.B(n_197),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_192),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_126),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_151),
.A2(n_108),
.B1(n_91),
.B2(n_88),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_126),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_149),
.A2(n_89),
.B1(n_102),
.B2(n_104),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_202),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_263)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_150),
.A2(n_138),
.B1(n_144),
.B2(n_53),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_204),
.A2(n_120),
.B(n_167),
.Y(n_256)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_205),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_122),
.A2(n_35),
.B1(n_28),
.B2(n_23),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_116),
.A2(n_71),
.B1(n_61),
.B2(n_35),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_140),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_215),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_111),
.B(n_72),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_139),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_130),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_213),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_67),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_164),
.A2(n_47),
.B(n_45),
.C(n_16),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_216),
.A2(n_120),
.B(n_44),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_223),
.Y(n_245)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_141),
.A2(n_89),
.B1(n_45),
.B2(n_16),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_219),
.A2(n_221),
.B1(n_127),
.B2(n_158),
.Y(n_265)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_220),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_116),
.A2(n_44),
.B1(n_70),
.B2(n_39),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_114),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_225),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_70),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_229),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_125),
.B(n_39),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_227),
.Y(n_250)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_143),
.Y(n_228)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

AO21x2_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_173),
.B(n_44),
.Y(n_243)
);

AO22x2_ASAP7_75t_L g300 ( 
.A1(n_243),
.A2(n_212),
.B1(n_133),
.B2(n_142),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_248),
.B(n_256),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_223),
.A2(n_143),
.B1(n_127),
.B2(n_121),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_251),
.Y(n_291)
);

OR2x2_ASAP7_75t_SL g254 ( 
.A(n_177),
.B(n_115),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_SL g289 ( 
.A(n_254),
.B(n_224),
.C(n_183),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_267),
.B1(n_268),
.B2(n_183),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g264 ( 
.A(n_222),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_197),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_204),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_180),
.A2(n_158),
.B1(n_112),
.B2(n_166),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_180),
.A2(n_112),
.B1(n_166),
.B2(n_157),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_254),
.C(n_252),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_272),
.B(n_263),
.C(n_265),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_226),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_273),
.B(n_281),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_274),
.A2(n_283),
.B(n_286),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_275),
.Y(n_318)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_277),
.A2(n_290),
.B1(n_280),
.B2(n_291),
.Y(n_316)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_280),
.A2(n_299),
.B1(n_301),
.B2(n_231),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_241),
.B(n_229),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_211),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_285),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_248),
.A2(n_214),
.B(n_181),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_181),
.C(n_211),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_284),
.B(n_290),
.Y(n_331)
);

O2A1O1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_243),
.A2(n_194),
.B(n_178),
.C(n_216),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_242),
.A2(n_179),
.B(n_214),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_178),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_292),
.Y(n_314)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_289),
.B(n_293),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_259),
.A2(n_215),
.B(n_208),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

AOI32xp33_ASAP7_75t_L g293 ( 
.A1(n_260),
.A2(n_218),
.A3(n_128),
.B1(n_170),
.B2(n_205),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_294),
.B(n_295),
.Y(n_302)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_257),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_259),
.B(n_188),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_297),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_298),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_263),
.A2(n_182),
.B1(n_157),
.B2(n_139),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_243),
.B1(n_238),
.B2(n_266),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_234),
.B(n_210),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_307),
.A2(n_310),
.B1(n_311),
.B2(n_315),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_309),
.B(n_264),
.C(n_239),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_299),
.A2(n_243),
.B1(n_209),
.B2(n_236),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_280),
.A2(n_243),
.B1(n_236),
.B2(n_207),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_317),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_277),
.A2(n_279),
.B1(n_273),
.B2(n_289),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_283),
.A2(n_201),
.B1(n_235),
.B2(n_176),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_323),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_272),
.B(n_284),
.C(n_282),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_331),
.C(n_328),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_300),
.A2(n_235),
.B1(n_187),
.B2(n_184),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_300),
.A2(n_200),
.B1(n_189),
.B2(n_246),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_325),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_300),
.A2(n_285),
.B1(n_281),
.B2(n_291),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_300),
.A2(n_213),
.B1(n_190),
.B2(n_220),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_296),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_305),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_332),
.B(n_351),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_330),
.A2(n_270),
.B(n_271),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_334),
.A2(n_337),
.B(n_341),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_312),
.B(n_288),
.Y(n_336)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_330),
.A2(n_276),
.B(n_278),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_345),
.C(n_360),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_311),
.A2(n_295),
.B(n_294),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_349),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_298),
.Y(n_344)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_293),
.C(n_286),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_325),
.A2(n_247),
.B(n_190),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_346),
.A2(n_353),
.B(n_316),
.Y(n_372)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_315),
.A2(n_244),
.B(n_239),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_358),
.Y(n_364)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_237),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_350),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_319),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_233),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_352),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_328),
.A2(n_247),
.B(n_213),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_306),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_354),
.Y(n_382)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_306),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_306),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_356),
.B(n_303),
.Y(n_366)
);

XOR2x2_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_233),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_357),
.A2(n_309),
.B(n_303),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_232),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_308),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_359),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_232),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_366),
.B(n_368),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_360),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_317),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_380),
.C(n_357),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_371),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_372),
.A2(n_381),
.B(n_343),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_339),
.A2(n_329),
.B1(n_327),
.B2(n_307),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_373),
.A2(n_385),
.B1(n_387),
.B2(n_390),
.Y(n_413)
);

INVxp33_ASAP7_75t_L g401 ( 
.A(n_375),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_338),
.A2(n_310),
.B1(n_324),
.B2(n_323),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_376),
.A2(n_347),
.B1(n_335),
.B2(n_341),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_327),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_384),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_345),
.B(n_314),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_333),
.A2(n_320),
.B(n_314),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_336),
.B(n_320),
.Y(n_383)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_383),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_345),
.B(n_302),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_339),
.A2(n_318),
.B1(n_302),
.B2(n_313),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_338),
.A2(n_326),
.B1(n_313),
.B2(n_308),
.Y(n_386)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_386),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_347),
.A2(n_326),
.B1(n_246),
.B2(n_262),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_347),
.A2(n_262),
.B1(n_244),
.B2(n_255),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_367),
.B(n_352),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_391),
.B(n_397),
.Y(n_429)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_392),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_395),
.B(n_410),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_356),
.C(n_357),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_404),
.C(n_406),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_344),
.Y(n_397)
);

INVx4_ASAP7_75t_SL g399 ( 
.A(n_382),
.Y(n_399)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_399),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_362),
.B(n_358),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g423 ( 
.A(n_400),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_402),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_334),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_403),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_356),
.C(n_333),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_365),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_405),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_353),
.C(n_349),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_388),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_407),
.B(n_409),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_370),
.B(n_346),
.C(n_334),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_366),
.C(n_384),
.Y(n_426)
);

INVx8_ASAP7_75t_L g409 ( 
.A(n_361),
.Y(n_409)
);

AOI221xp5_ASAP7_75t_L g410 ( 
.A1(n_371),
.A2(n_337),
.B1(n_341),
.B2(n_335),
.C(n_332),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_411),
.A2(n_419),
.B1(n_387),
.B2(n_390),
.Y(n_438)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_388),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_412),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_354),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_414),
.A2(n_393),
.B1(n_399),
.B2(n_418),
.Y(n_425)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_379),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_416),
.B(n_417),
.Y(n_437)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_379),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_364),
.A2(n_347),
.B1(n_337),
.B2(n_350),
.Y(n_419)
);

XOR2x2_ASAP7_75t_L g420 ( 
.A(n_418),
.B(n_380),
.Y(n_420)
);

XOR2x2_ASAP7_75t_L g463 ( 
.A(n_420),
.B(n_199),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_413),
.A2(n_364),
.B1(n_398),
.B2(n_372),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_422),
.A2(n_433),
.B1(n_439),
.B2(n_441),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_425),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_394),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_378),
.C(n_377),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_430),
.C(n_415),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_395),
.C(n_415),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_413),
.A2(n_364),
.B1(n_376),
.B2(n_373),
.Y(n_433)
);

FAx1_ASAP7_75t_SL g434 ( 
.A(n_396),
.B(n_377),
.CI(n_381),
.CON(n_434),
.SN(n_434)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_434),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_438),
.A2(n_392),
.B1(n_412),
.B2(n_405),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_411),
.A2(n_363),
.B1(n_369),
.B2(n_359),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_419),
.A2(n_369),
.B1(n_348),
.B2(n_342),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_402),
.A2(n_355),
.B1(n_228),
.B2(n_255),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_443),
.A2(n_355),
.B1(n_409),
.B2(n_401),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_446),
.A2(n_457),
.B1(n_230),
.B2(n_203),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_435),
.A2(n_403),
.B(n_429),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_447),
.B(n_450),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_452),
.Y(n_468)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_436),
.Y(n_451)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_451),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_394),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_453),
.A2(n_431),
.B1(n_428),
.B2(n_440),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_432),
.B(n_408),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_454),
.B(n_426),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_422),
.A2(n_401),
.B(n_264),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_456),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_437),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_438),
.A2(n_133),
.B1(n_142),
.B2(n_192),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_436),
.Y(n_458)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_458),
.Y(n_476)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_421),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_459),
.Y(n_479)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_428),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_460),
.B(n_442),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_423),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_461),
.B(n_443),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_433),
.A2(n_195),
.B1(n_230),
.B2(n_237),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_462),
.A2(n_174),
.B1(n_193),
.B2(n_12),
.Y(n_481)
);

XNOR2x1_ASAP7_75t_L g464 ( 
.A(n_463),
.B(n_427),
.Y(n_464)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_475),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_424),
.C(n_430),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_466),
.B(n_474),
.C(n_457),
.Y(n_495)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_467),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_477),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_448),
.C(n_449),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_424),
.C(n_420),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_445),
.B(n_434),
.Y(n_475)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_447),
.B(n_434),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_444),
.A2(n_439),
.B1(n_437),
.B2(n_441),
.Y(n_478)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_478),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_480),
.A2(n_462),
.B1(n_479),
.B2(n_476),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_481),
.B(n_453),
.Y(n_484)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_484),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_466),
.B(n_449),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_486),
.B(n_487),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_469),
.B(n_444),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_474),
.A2(n_455),
.B(n_452),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_488),
.A2(n_471),
.B1(n_479),
.B2(n_468),
.Y(n_502)
);

FAx1_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_463),
.CI(n_446),
.CON(n_489),
.SN(n_489)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_489),
.B(n_494),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_470),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_491),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_492),
.B(n_468),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g494 ( 
.A(n_473),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_495),
.B(n_496),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_464),
.B(n_39),
.C(n_193),
.Y(n_496)
);

XNOR2x1_ASAP7_75t_L g515 ( 
.A(n_498),
.B(n_501),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_495),
.B(n_465),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_505),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_481),
.Y(n_504)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_504),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_485),
.A2(n_4),
.B1(n_13),
.B2(n_12),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_496),
.B(n_4),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_507),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_485),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_507)
);

INVx11_ASAP7_75t_L g510 ( 
.A(n_489),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_510),
.B(n_14),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_508),
.A2(n_482),
.B(n_493),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_511),
.A2(n_514),
.B(n_509),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_500),
.A2(n_497),
.B(n_489),
.Y(n_514)
);

NOR2xp67_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_11),
.Y(n_516)
);

A2O1A1Ixp33_ASAP7_75t_L g524 ( 
.A1(n_516),
.A2(n_518),
.B(n_503),
.C(n_513),
.Y(n_524)
);

OAI21xp33_ASAP7_75t_L g518 ( 
.A1(n_499),
.A2(n_11),
.B(n_13),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_507),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_515),
.B(n_498),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_521),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_517),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g528 ( 
.A1(n_522),
.A2(n_524),
.B(n_525),
.Y(n_528)
);

O2A1O1Ixp5_ASAP7_75t_L g527 ( 
.A1(n_523),
.A2(n_506),
.B(n_14),
.C(n_2),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_512),
.A2(n_504),
.B(n_501),
.Y(n_525)
);

O2A1O1Ixp33_ASAP7_75t_SL g529 ( 
.A1(n_527),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_529)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_529),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_528),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_531),
.B(n_526),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_530),
.C(n_1),
.Y(n_533)
);

A2O1A1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_534)
);

OA21x2_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_3),
.B(n_531),
.Y(n_535)
);


endmodule