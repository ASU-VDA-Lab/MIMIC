module fake_jpeg_12496_n_173 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_34),
.A2(n_18),
.B(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_44),
.Y(n_65)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_46),
.Y(n_82)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_14),
.Y(n_77)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_12),
.Y(n_84)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

CKINVDCx6p67_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g60 ( 
.A1(n_34),
.A2(n_20),
.B(n_16),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_42),
.B(n_54),
.C(n_21),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_18),
.B1(n_30),
.B2(n_20),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_39),
.B1(n_2),
.B2(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_40),
.B(n_25),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_8),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_33),
.A2(n_35),
.B1(n_47),
.B2(n_50),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_73),
.B1(n_37),
.B2(n_41),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_81),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_12),
.B1(n_16),
.B2(n_28),
.Y(n_73)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_46),
.B(n_25),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_26),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_85),
.B(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_48),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_95),
.Y(n_118)
);

AO22x1_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_42),
.B1(n_49),
.B2(n_54),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_105),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_55),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_102),
.Y(n_108)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_21),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_103),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_107),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_8),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_11),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_104),
.A2(n_71),
.B1(n_63),
.B2(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_1),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_76),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_4),
.C(n_6),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_97),
.C(n_99),
.Y(n_128)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_69),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_122),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_64),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_70),
.B1(n_58),
.B2(n_57),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_57),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_98),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_127),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_133),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_105),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_125),
.C(n_111),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_95),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_116),
.B(n_108),
.C(n_112),
.D(n_94),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_121),
.Y(n_144)
);

AO22x1_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_92),
.B1(n_112),
.B2(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_109),
.B(n_63),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_144),
.B(n_117),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_128),
.B(n_135),
.C(n_137),
.D(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_145),
.B(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

OAI321xp33_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_138),
.A3(n_137),
.B1(n_134),
.B2(n_131),
.C(n_108),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_151),
.B1(n_152),
.B2(n_155),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_134),
.B(n_78),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_113),
.C(n_93),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_142),
.B1(n_143),
.B2(n_146),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_86),
.B(n_58),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_140),
.B1(n_156),
.B2(n_145),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_124),
.B(n_113),
.C(n_89),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_163),
.B(n_164),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_61),
.B(n_68),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_157),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_166),
.B(n_167),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_157),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_161),
.C(n_68),
.Y(n_170)
);

AOI21x1_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_161),
.B(n_68),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_169),
.Y(n_173)
);


endmodule