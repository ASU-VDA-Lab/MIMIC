module fake_netlist_5_991_n_1711 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1711);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1711;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1556;
wire n_1384;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1534;
wire n_560;
wire n_1354;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_109),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_39),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_64),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_61),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_96),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_91),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_77),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_124),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_75),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_117),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_100),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_86),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_13),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_139),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_7),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_45),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_110),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_113),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_76),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_20),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_47),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_47),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_25),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_69),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_56),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_120),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_38),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_154),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_44),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_34),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_51),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_92),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_37),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_123),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_84),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_14),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_41),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_11),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_30),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_43),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_79),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_150),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_144),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_34),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_23),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_155),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_98),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_146),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_127),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_49),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_38),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_24),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_17),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_133),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_82),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_105),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_28),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_142),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_153),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_102),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_115),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_23),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_42),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_99),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_71),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_20),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_1),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_28),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_36),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_95),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_112),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_93),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_52),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_43),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_108),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_21),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_128),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_134),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_42),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_19),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_74),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_141),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_114),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_27),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_15),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_19),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_33),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_130),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_106),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_83),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_81),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_94),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_41),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_48),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_37),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_104),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_55),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_103),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_4),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_12),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_131),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_58),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_1),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_18),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_25),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_107),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_63),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_27),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_89),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_73),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_60),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_36),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_57),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_48),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_80),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_17),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_30),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_31),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_136),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_15),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_5),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_156),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_140),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_21),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_101),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_119),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_31),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_52),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_55),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_152),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_68),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_151),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_125),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_10),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_4),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_26),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_14),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_78),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_85),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_5),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_8),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_8),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_9),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_59),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_32),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_65),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_90),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_277),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_170),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_157),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_277),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_240),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_160),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_277),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_277),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_170),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_277),
.B(n_0),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_161),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_277),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_181),
.B(n_0),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_181),
.B(n_2),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_182),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_163),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_162),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_165),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_166),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_310),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_158),
.B(n_2),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_219),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_182),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_164),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_182),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_187),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_167),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_187),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_182),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_182),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_194),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_169),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_172),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_248),
.B(n_3),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_194),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_200),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_200),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_159),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_174),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_177),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_229),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_295),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_168),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_178),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_173),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_226),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_226),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_179),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_180),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_278),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_278),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_302),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_291),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_183),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_175),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_199),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_291),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_180),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_191),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_199),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_185),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_185),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_193),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_302),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_193),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_L g382 ( 
.A(n_248),
.B(n_3),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_202),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_210),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_222),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_202),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_204),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_331),
.Y(n_389)
);

CKINVDCx6p67_ASAP7_75t_R g390 ( 
.A(n_336),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_313),
.B(n_323),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_372),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_196),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_331),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_344),
.B(n_368),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_312),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_339),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_198),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_339),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_372),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_372),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_341),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_341),
.B(n_345),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_345),
.B(n_158),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_315),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_346),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_346),
.B(n_205),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_350),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_376),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_315),
.B(n_184),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_318),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_318),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_320),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_320),
.B(n_242),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_322),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_314),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_337),
.B(n_239),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_326),
.B(n_184),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_371),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_326),
.B(n_206),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_316),
.B(n_192),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_374),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_327),
.B(n_192),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_350),
.Y(n_429)
);

OAI21x1_ASAP7_75t_L g430 ( 
.A1(n_327),
.A2(n_283),
.B(n_242),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_329),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_378),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_378),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_379),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_329),
.Y(n_435)
);

OA21x2_ASAP7_75t_L g436 ( 
.A1(n_324),
.A2(n_209),
.B(n_204),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_347),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_347),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_351),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_351),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_352),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_352),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_353),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_353),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_362),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_362),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_354),
.Y(n_447)
);

CKINVDCx8_ASAP7_75t_R g448 ( 
.A(n_317),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_366),
.Y(n_451)
);

CKINVDCx11_ASAP7_75t_R g452 ( 
.A(n_333),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_328),
.A2(n_171),
.B1(n_186),
.B2(n_280),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_367),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_367),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_421),
.A2(n_330),
.B1(n_321),
.B2(n_382),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_L g458 ( 
.A(n_409),
.B(n_429),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_421),
.B(n_319),
.Y(n_459)
);

OR2x6_ASAP7_75t_L g460 ( 
.A(n_391),
.B(n_225),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_418),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_391),
.B(n_325),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_409),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_332),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_436),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_418),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_452),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_418),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_388),
.Y(n_470)
);

AND3x2_ASAP7_75t_L g471 ( 
.A(n_393),
.B(n_283),
.C(n_235),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_423),
.B(n_336),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_423),
.B(n_357),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_436),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_419),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_453),
.B(n_340),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_453),
.A2(n_190),
.B1(n_217),
.B2(n_201),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_420),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_417),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_419),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_425),
.B(n_334),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_397),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_419),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_392),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_420),
.B(n_357),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_436),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_431),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_425),
.B(n_335),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_394),
.B(n_343),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_392),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_394),
.B(n_348),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_431),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_431),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

BUFx4f_ASAP7_75t_L g499 ( 
.A(n_436),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_435),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_392),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_396),
.B(n_411),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_392),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_436),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_399),
.B(n_349),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_399),
.B(n_355),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_435),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_393),
.B(n_358),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_392),
.Y(n_509)
);

AND2x2_ASAP7_75t_SL g510 ( 
.A(n_436),
.B(n_199),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_392),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_408),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_397),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_397),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_426),
.A2(n_382),
.B1(n_354),
.B2(n_268),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_452),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_401),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_397),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_411),
.B(n_199),
.Y(n_519)
);

NAND3xp33_ASAP7_75t_L g520 ( 
.A(n_426),
.B(n_422),
.C(n_411),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_447),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_406),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_401),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_406),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_393),
.B(n_358),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_406),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_406),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_447),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_413),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_408),
.B(n_356),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_401),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_422),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_401),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_447),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_413),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_390),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_422),
.B(n_360),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_448),
.A2(n_370),
.B1(n_375),
.B2(n_317),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_413),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_413),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_401),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_414),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_414),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_414),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_414),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_415),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_448),
.B(n_289),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_415),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_401),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_448),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_R g551 ( 
.A(n_428),
.B(n_176),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_415),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_428),
.B(n_369),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_428),
.B(n_207),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_390),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_415),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_389),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_417),
.B(n_225),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_389),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_389),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_417),
.B(n_377),
.C(n_365),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_430),
.B(n_235),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_401),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_389),
.B(n_417),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_390),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_417),
.A2(n_290),
.B1(n_241),
.B2(n_311),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_417),
.A2(n_273),
.B1(n_269),
.B2(n_259),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_424),
.B(n_427),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_424),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_395),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_430),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_395),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_410),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_404),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_427),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_395),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_398),
.B(n_211),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_398),
.B(n_212),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_401),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_439),
.B(n_373),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_432),
.B(n_289),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_432),
.B(n_289),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_433),
.B(n_189),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_404),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_398),
.Y(n_585)
);

INVx6_ASAP7_75t_L g586 ( 
.A(n_405),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_433),
.B(n_189),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_400),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_400),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_434),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_402),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_430),
.B(n_405),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_400),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_439),
.B(n_373),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_434),
.B(n_262),
.C(n_245),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_439),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_403),
.B(n_213),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_402),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_405),
.B(n_189),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_402),
.Y(n_600)
);

CKINVDCx16_ASAP7_75t_R g601 ( 
.A(n_405),
.Y(n_601)
);

AO22x2_ASAP7_75t_L g602 ( 
.A1(n_405),
.A2(n_243),
.B1(n_209),
.B2(n_215),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_405),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_SL g604 ( 
.A(n_444),
.B(n_188),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_403),
.B(n_218),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_462),
.B(n_359),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_SL g607 ( 
.A(n_459),
.B(n_245),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_512),
.A2(n_384),
.B1(n_361),
.B2(n_364),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_502),
.B(n_442),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_502),
.B(n_442),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_532),
.A2(n_296),
.B1(n_262),
.B2(n_270),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_532),
.B(n_270),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_506),
.B(n_574),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_463),
.B(n_385),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_574),
.B(n_442),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_463),
.B(n_220),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_532),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_557),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_584),
.B(n_442),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_569),
.B(n_223),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_584),
.B(n_485),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_492),
.B(n_442),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_575),
.B(n_224),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_493),
.B(n_195),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_570),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_590),
.B(n_228),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_553),
.B(n_456),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_537),
.B(n_234),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_495),
.B(n_456),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_557),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_505),
.B(n_197),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_530),
.B(n_456),
.Y(n_632)
);

XOR2x2_ASAP7_75t_L g633 ( 
.A(n_481),
.B(n_6),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_566),
.B(n_203),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_458),
.B(n_208),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_471),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_520),
.B(n_403),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_570),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_601),
.B(n_236),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_568),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_601),
.B(n_457),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_572),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_520),
.B(n_407),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_553),
.B(n_407),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_568),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_551),
.A2(n_460),
.B1(n_586),
.B2(n_465),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_460),
.A2(n_252),
.B1(n_308),
.B2(n_303),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_528),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_554),
.B(n_407),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_461),
.B(n_467),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_461),
.B(n_437),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_559),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_564),
.A2(n_410),
.B(n_441),
.Y(n_653)
);

NAND3xp33_ASAP7_75t_L g654 ( 
.A(n_515),
.B(n_261),
.C(n_263),
.Y(n_654)
);

AOI221xp5_ASAP7_75t_L g655 ( 
.A1(n_481),
.A2(n_244),
.B1(n_243),
.B2(n_230),
.C(n_221),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_460),
.B(n_444),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_538),
.B(n_246),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_460),
.A2(n_247),
.B1(n_253),
.B2(n_254),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_467),
.B(n_437),
.Y(n_659)
);

NOR2xp67_ASAP7_75t_L g660 ( 
.A(n_561),
.B(n_444),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_460),
.A2(n_296),
.B1(n_275),
.B2(n_199),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_567),
.B(n_255),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_559),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_472),
.B(n_214),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_469),
.B(n_437),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_572),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_567),
.B(n_534),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_473),
.B(n_216),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_534),
.B(n_256),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_547),
.B(n_227),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_469),
.B(n_437),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_SL g672 ( 
.A(n_596),
.B(n_275),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_SL g673 ( 
.A(n_565),
.B(n_189),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_576),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_560),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_560),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_576),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_478),
.A2(n_504),
.B1(n_490),
.B2(n_562),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_561),
.B(n_276),
.C(n_231),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_479),
.B(n_437),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_479),
.B(n_437),
.Y(n_681)
);

AOI221xp5_ASAP7_75t_L g682 ( 
.A1(n_480),
.A2(n_250),
.B1(n_221),
.B2(n_230),
.C(n_244),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_484),
.B(n_437),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_484),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_585),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_483),
.B(n_260),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_585),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_521),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_483),
.B(n_265),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_489),
.B(n_232),
.Y(n_690)
);

INVx5_ASAP7_75t_L g691 ( 
.A(n_592),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_508),
.B(n_233),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_588),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_487),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_487),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_588),
.Y(n_696)
);

OR2x2_ASAP7_75t_SL g697 ( 
.A(n_550),
.B(n_480),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_491),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_562),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_483),
.B(n_482),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_478),
.A2(n_437),
.B1(n_438),
.B2(n_443),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_499),
.A2(n_271),
.B1(n_274),
.B2(n_279),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_491),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_496),
.B(n_438),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_466),
.B(n_287),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_478),
.A2(n_438),
.B1(n_443),
.B2(n_215),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_496),
.Y(n_707)
);

INVxp33_ASAP7_75t_L g708 ( 
.A(n_525),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_562),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_497),
.Y(n_710)
);

NAND2x1p5_ASAP7_75t_L g711 ( 
.A(n_592),
.B(n_402),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_490),
.A2(n_438),
.B1(n_443),
.B2(n_250),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_562),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_589),
.Y(n_714)
);

O2A1O1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_466),
.A2(n_257),
.B(n_258),
.C(n_264),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_497),
.B(n_438),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_589),
.Y(n_717)
);

NOR3xp33_ASAP7_75t_L g718 ( 
.A(n_550),
.B(n_249),
.C(n_238),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_498),
.B(n_438),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_592),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_593),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_593),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_490),
.A2(n_257),
.B(n_258),
.C(n_264),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_500),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_507),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_483),
.B(n_294),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_507),
.B(n_438),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_604),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_510),
.B(n_438),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_510),
.B(n_443),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_592),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_510),
.B(n_443),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_580),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_580),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_577),
.B(n_443),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_581),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_578),
.B(n_443),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_605),
.B(n_443),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_573),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_482),
.B(n_297),
.Y(n_740)
);

NOR3xp33_ASAP7_75t_L g741 ( 
.A(n_582),
.B(n_304),
.C(n_251),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_597),
.B(n_440),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_468),
.B(n_379),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_586),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_504),
.A2(n_268),
.B1(n_300),
.B2(n_299),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_573),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_573),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_571),
.B(n_440),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_482),
.B(n_286),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_L g750 ( 
.A(n_519),
.B(n_402),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_602),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_594),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_482),
.B(n_603),
.Y(n_753)
);

BUFx6f_ASAP7_75t_SL g754 ( 
.A(n_558),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_518),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_594),
.Y(n_756)
);

NOR2xp67_ASAP7_75t_L g757 ( 
.A(n_595),
.B(n_449),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_518),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_571),
.B(n_440),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_518),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_602),
.B(n_455),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_586),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_603),
.B(n_286),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_526),
.Y(n_764)
);

NOR3xp33_ASAP7_75t_L g765 ( 
.A(n_583),
.B(n_237),
.C(n_266),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_571),
.B(n_440),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_586),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_602),
.B(n_449),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_513),
.B(n_441),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_513),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_526),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_514),
.B(n_441),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_514),
.B(n_522),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_522),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_524),
.B(n_441),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_729),
.A2(n_499),
.B(n_504),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_730),
.A2(n_499),
.B(n_558),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_691),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_732),
.A2(n_759),
.B(n_748),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_613),
.B(n_524),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_699),
.A2(n_558),
.B(n_464),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_699),
.A2(n_713),
.B(n_709),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_709),
.A2(n_558),
.B(n_464),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_621),
.A2(n_599),
.B1(n_558),
.B2(n_603),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_678),
.A2(n_646),
.B1(n_731),
.B2(n_720),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_624),
.A2(n_603),
.B1(n_587),
.B2(n_602),
.Y(n_786)
);

NAND2xp33_ASAP7_75t_SL g787 ( 
.A(n_708),
.B(n_536),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_713),
.A2(n_476),
.B(n_486),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_766),
.A2(n_545),
.B(n_527),
.Y(n_789)
);

O2A1O1Ixp5_ASAP7_75t_L g790 ( 
.A1(n_637),
.A2(n_595),
.B(n_598),
.C(n_600),
.Y(n_790)
);

AOI33xp33_ASAP7_75t_L g791 ( 
.A1(n_682),
.A2(n_305),
.A3(n_272),
.B1(n_284),
.B2(n_293),
.B3(n_298),
.Y(n_791)
);

A2O1A1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_631),
.A2(n_544),
.B(n_527),
.C(n_535),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_691),
.B(n_536),
.Y(n_793)
);

INVx8_ASAP7_75t_L g794 ( 
.A(n_754),
.Y(n_794)
);

INVx5_ASAP7_75t_L g795 ( 
.A(n_720),
.Y(n_795)
);

AOI21xp33_ASAP7_75t_L g796 ( 
.A1(n_634),
.A2(n_555),
.B(n_267),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_609),
.A2(n_470),
.B(n_475),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_691),
.A2(n_488),
.B(n_511),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_617),
.B(n_535),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_720),
.A2(n_555),
.B1(n_544),
.B2(n_545),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_640),
.B(n_516),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_691),
.B(n_286),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_691),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_688),
.B(n_281),
.Y(n_804)
);

BUFx5_ASAP7_75t_L g805 ( 
.A(n_762),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_617),
.Y(n_806)
);

BUFx4f_ASAP7_75t_SL g807 ( 
.A(n_614),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_640),
.A2(n_540),
.B(n_526),
.C(n_552),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_648),
.B(n_282),
.Y(n_809)
);

AO21x2_ASAP7_75t_L g810 ( 
.A1(n_705),
.A2(n_529),
.B(n_556),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_743),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_635),
.B(n_286),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_641),
.A2(n_519),
.B1(n_486),
.B2(n_470),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_670),
.A2(n_529),
.B(n_475),
.C(n_476),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_739),
.Y(n_815)
);

OAI21xp33_ASAP7_75t_L g816 ( 
.A1(n_655),
.A2(n_285),
.B(n_288),
.Y(n_816)
);

OAI21xp33_ASAP7_75t_L g817 ( 
.A1(n_664),
.A2(n_292),
.B(n_301),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_606),
.B(n_306),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_752),
.A2(n_539),
.B1(n_548),
.B2(n_542),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_684),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_743),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_742),
.A2(n_488),
.B(n_511),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_667),
.B(n_307),
.Y(n_823)
);

BUFx6f_ASAP7_75t_SL g824 ( 
.A(n_636),
.Y(n_824)
);

OAI21xp33_ASAP7_75t_L g825 ( 
.A1(n_668),
.A2(n_293),
.B(n_284),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_711),
.Y(n_826)
);

AO21x1_ASAP7_75t_L g827 ( 
.A1(n_607),
.A2(n_298),
.B(n_299),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_739),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_735),
.A2(n_488),
.B(n_511),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_708),
.B(n_474),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_737),
.A2(n_488),
.B(n_511),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_752),
.B(n_539),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_645),
.B(n_523),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_684),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_738),
.A2(n_610),
.B(n_629),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_728),
.A2(n_542),
.B1(n_543),
.B2(n_546),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_636),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_733),
.B(n_381),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_627),
.B(n_649),
.Y(n_839)
);

NOR2xp67_ASAP7_75t_L g840 ( 
.A(n_736),
.B(n_381),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_627),
.B(n_734),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_622),
.A2(n_523),
.B(n_541),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_756),
.B(n_383),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_632),
.A2(n_523),
.B(n_541),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_746),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_656),
.A2(n_543),
.B(n_546),
.C(n_548),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_711),
.A2(n_523),
.B(n_541),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_711),
.A2(n_705),
.B(n_744),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_744),
.A2(n_767),
.B(n_619),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_656),
.B(n_615),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_643),
.A2(n_552),
.B1(n_556),
.B2(n_540),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_694),
.B(n_540),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_L g853 ( 
.A(n_767),
.B(n_519),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_706),
.A2(n_600),
.B(n_598),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_695),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_762),
.A2(n_519),
.B1(n_598),
.B2(n_600),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_761),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_695),
.B(n_474),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_698),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_723),
.A2(n_272),
.B(n_300),
.C(n_305),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_692),
.B(n_383),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_698),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_703),
.B(n_474),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_761),
.B(n_386),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_703),
.B(n_474),
.Y(n_865)
);

AOI21xp33_ASAP7_75t_L g866 ( 
.A1(n_690),
.A2(n_449),
.B(n_451),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_712),
.A2(n_600),
.B(n_598),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_673),
.B(n_523),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_746),
.Y(n_869)
);

NOR3xp33_ASAP7_75t_L g870 ( 
.A(n_608),
.B(n_386),
.C(n_387),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_707),
.Y(n_871)
);

BUFx12f_ASAP7_75t_L g872 ( 
.A(n_636),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_747),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_707),
.B(n_477),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_662),
.B(n_477),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_745),
.A2(n_725),
.B1(n_710),
.B2(n_724),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_620),
.B(n_477),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_710),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_724),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_616),
.B(n_387),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_725),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_747),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_650),
.A2(n_501),
.B(n_579),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_660),
.B(n_477),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_672),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_612),
.B(n_494),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_644),
.A2(n_501),
.B(n_579),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_618),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_661),
.A2(n_501),
.B1(n_579),
.B2(n_563),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_669),
.B(n_451),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_612),
.B(n_494),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_751),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_612),
.B(n_494),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_651),
.A2(n_494),
.B(n_563),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_607),
.A2(n_503),
.B(n_563),
.C(n_509),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_618),
.B(n_503),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_630),
.B(n_503),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_647),
.B(n_523),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_659),
.A2(n_671),
.B(n_665),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_751),
.A2(n_533),
.B1(n_563),
.B2(n_517),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_625),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_658),
.B(n_541),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_680),
.A2(n_531),
.B(n_517),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_697),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_768),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_630),
.B(n_503),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_623),
.B(n_533),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_626),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_768),
.B(n_451),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_625),
.Y(n_910)
);

CKINVDCx20_ASAP7_75t_R g911 ( 
.A(n_697),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_681),
.A2(n_531),
.B(n_509),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_652),
.B(n_509),
.Y(n_913)
);

CKINVDCx10_ASAP7_75t_R g914 ( 
.A(n_754),
.Y(n_914)
);

AOI21x1_ASAP7_75t_L g915 ( 
.A1(n_683),
.A2(n_410),
.B(n_450),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_652),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_740),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_654),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_628),
.B(n_591),
.Y(n_919)
);

OAI321xp33_ASAP7_75t_L g920 ( 
.A1(n_657),
.A2(n_454),
.A3(n_455),
.B1(n_450),
.B2(n_445),
.C(n_446),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_749),
.B(n_533),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_704),
.A2(n_533),
.B(n_531),
.Y(n_922)
);

NOR3xp33_ASAP7_75t_L g923 ( 
.A(n_718),
.B(n_454),
.C(n_455),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_639),
.B(n_531),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_633),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_663),
.B(n_517),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_638),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_675),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_675),
.B(n_519),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_676),
.Y(n_930)
);

NAND2x1_ASAP7_75t_L g931 ( 
.A(n_755),
.B(n_591),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_611),
.A2(n_676),
.B1(n_679),
.B2(n_687),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_770),
.B(n_519),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_770),
.B(n_519),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_638),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_773),
.A2(n_412),
.B(n_450),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_716),
.A2(n_591),
.B(n_549),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_702),
.B(n_591),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_719),
.A2(n_591),
.B(n_549),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_715),
.A2(n_454),
.B(n_445),
.C(n_446),
.Y(n_940)
);

INVx11_ASAP7_75t_L g941 ( 
.A(n_741),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_727),
.A2(n_591),
.B(n_549),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_765),
.B(n_450),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_774),
.B(n_549),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_774),
.B(n_549),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_701),
.A2(n_549),
.B(n_541),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_753),
.B(n_541),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_642),
.A2(n_412),
.B(n_445),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_666),
.A2(n_412),
.B(n_445),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_653),
.A2(n_412),
.B(n_402),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_769),
.A2(n_412),
.B(n_402),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_666),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_763),
.A2(n_446),
.B(n_7),
.C(n_9),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_754),
.Y(n_954)
);

NAND2x1_ASAP7_75t_L g955 ( 
.A(n_755),
.B(n_402),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_700),
.B(n_446),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_633),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_686),
.B(n_6),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_861),
.B(n_757),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_820),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_839),
.B(n_721),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_784),
.A2(n_689),
.B1(n_726),
.B2(n_722),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_841),
.B(n_909),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_909),
.B(n_721),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_811),
.B(n_717),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_821),
.B(n_717),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_864),
.B(n_714),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_780),
.A2(n_722),
.B(n_677),
.C(n_685),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_848),
.A2(n_750),
.B(n_775),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_834),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_935),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_864),
.B(n_696),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_835),
.A2(n_938),
.B(n_779),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_946),
.A2(n_750),
.B(n_772),
.Y(n_974)
);

OAI22xp33_ASAP7_75t_L g975 ( 
.A1(n_807),
.A2(n_696),
.B1(n_677),
.B2(n_685),
.Y(n_975)
);

NAND3xp33_ASAP7_75t_L g976 ( 
.A(n_818),
.B(n_714),
.C(n_674),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_857),
.B(n_693),
.Y(n_977)
);

AOI221xp5_ASAP7_75t_L g978 ( 
.A1(n_957),
.A2(n_693),
.B1(n_687),
.B2(n_674),
.C(n_758),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_850),
.B(n_764),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_R g980 ( 
.A(n_787),
.B(n_771),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_876),
.A2(n_771),
.B(n_764),
.C(n_760),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_946),
.A2(n_760),
.B(n_758),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_776),
.A2(n_416),
.B(n_148),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_801),
.Y(n_984)
);

BUFx4f_ASAP7_75t_L g985 ( 
.A(n_872),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_958),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_892),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_954),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_855),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_823),
.A2(n_416),
.B(n_16),
.C(n_18),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_918),
.A2(n_13),
.B(n_16),
.C(n_22),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_R g992 ( 
.A(n_904),
.B(n_911),
.Y(n_992)
);

AOI21x1_ASAP7_75t_L g993 ( 
.A1(n_777),
.A2(n_416),
.B(n_147),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_857),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_885),
.B(n_22),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_857),
.B(n_905),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_859),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_871),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_785),
.A2(n_416),
.B1(n_145),
.B2(n_138),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_908),
.A2(n_416),
.B1(n_137),
.B2(n_135),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_905),
.B(n_416),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_777),
.A2(n_786),
.B(n_817),
.C(n_796),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_905),
.B(n_24),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_776),
.A2(n_416),
.B(n_126),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_804),
.B(n_26),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_790),
.A2(n_416),
.B(n_116),
.Y(n_1006)
);

NAND2x1p5_ASAP7_75t_L g1007 ( 
.A(n_803),
.B(n_416),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_862),
.B(n_29),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_930),
.B(n_97),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_837),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_866),
.A2(n_29),
.B(n_32),
.C(n_33),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_847),
.A2(n_88),
.B(n_87),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_880),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_794),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_794),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_875),
.A2(n_924),
.B(n_907),
.C(n_877),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_829),
.A2(n_72),
.B(n_70),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_935),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_825),
.A2(n_35),
.B(n_39),
.C(n_40),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_879),
.A2(n_35),
.B(n_40),
.C(n_44),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_838),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_778),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_830),
.B(n_45),
.Y(n_1023)
);

AO21x1_ASAP7_75t_L g1024 ( 
.A1(n_812),
.A2(n_46),
.B(n_49),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_778),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_781),
.A2(n_46),
.B(n_50),
.C(n_51),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_890),
.B(n_50),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_854),
.A2(n_67),
.B(n_66),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_928),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_831),
.A2(n_62),
.B(n_54),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_878),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_878),
.B(n_53),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_881),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_943),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_925),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_881),
.B(n_53),
.Y(n_1036)
);

NOR2xp67_ASAP7_75t_SL g1037 ( 
.A(n_795),
.B(n_54),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_781),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_809),
.B(n_917),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_943),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_888),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_941),
.B(n_930),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_842),
.A2(n_844),
.B(n_822),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_843),
.B(n_888),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_940),
.A2(n_860),
.B(n_792),
.C(n_832),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_826),
.A2(n_930),
.B1(n_916),
.B2(n_795),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_806),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_SL g1048 ( 
.A1(n_921),
.A2(n_923),
.B(n_870),
.C(n_920),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_783),
.A2(n_953),
.B(n_782),
.C(n_932),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_789),
.A2(n_893),
.B(n_891),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_886),
.A2(n_898),
.B(n_902),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_778),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_846),
.A2(n_900),
.B(n_895),
.C(n_800),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_795),
.B(n_840),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_833),
.A2(n_868),
.B(n_814),
.C(n_852),
.Y(n_1055)
);

NOR3xp33_ASAP7_75t_SL g1056 ( 
.A(n_816),
.B(n_793),
.C(n_802),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_819),
.A2(n_916),
.B(n_836),
.C(n_808),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_826),
.B(n_824),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_901),
.B(n_910),
.Y(n_1059)
);

OAI21xp33_ASAP7_75t_L g1060 ( 
.A1(n_791),
.A2(n_813),
.B(n_874),
.Y(n_1060)
);

NAND2xp33_ASAP7_75t_SL g1061 ( 
.A(n_824),
.B(n_803),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_795),
.A2(n_945),
.B1(n_944),
.B2(n_929),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_927),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_827),
.A2(n_952),
.B1(n_805),
.B2(n_919),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_815),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_851),
.A2(n_799),
.B(n_865),
.C(n_863),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_914),
.Y(n_1067)
);

NAND3xp33_ASAP7_75t_L g1068 ( 
.A(n_783),
.B(n_782),
.C(n_884),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_899),
.B(n_882),
.Y(n_1069)
);

AOI221xp5_ASAP7_75t_L g1070 ( 
.A1(n_794),
.A2(n_899),
.B1(n_887),
.B2(n_889),
.C(n_947),
.Y(n_1070)
);

OAI21xp33_ASAP7_75t_L g1071 ( 
.A1(n_858),
.A2(n_906),
.B(n_926),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_828),
.B(n_873),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_845),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_896),
.A2(n_913),
.B(n_897),
.C(n_869),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_798),
.A2(n_849),
.B(n_853),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_933),
.A2(n_934),
.B1(n_856),
.B2(n_854),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_887),
.B(n_805),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_915),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_805),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_805),
.B(n_797),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_788),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_805),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_788),
.Y(n_1083)
);

INVx6_ASAP7_75t_L g1084 ( 
.A(n_931),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_955),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_867),
.A2(n_883),
.B1(n_937),
.B2(n_939),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_956),
.A2(n_810),
.B1(n_883),
.B2(n_894),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_894),
.B(n_903),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_936),
.B(n_903),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_912),
.A2(n_922),
.B(n_939),
.C(n_942),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_912),
.A2(n_922),
.B1(n_810),
.B2(n_948),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_949),
.A2(n_613),
.B1(n_678),
.B2(n_621),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_951),
.B(n_950),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_951),
.B(n_950),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_861),
.B(n_613),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_823),
.A2(n_613),
.B(n_621),
.C(n_958),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_811),
.B(n_613),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_848),
.A2(n_691),
.B(n_699),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_SL g1099 ( 
.A(n_811),
.B(n_482),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_811),
.B(n_613),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_935),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_821),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_861),
.B(n_613),
.Y(n_1103)
);

NAND2x1p5_ASAP7_75t_L g1104 ( 
.A(n_803),
.B(n_691),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_984),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1051),
.A2(n_1098),
.B(n_1094),
.Y(n_1106)
);

INVx3_ASAP7_75t_SL g1107 ( 
.A(n_1067),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_992),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1097),
.B(n_1100),
.Y(n_1109)
);

OR2x6_ASAP7_75t_L g1110 ( 
.A(n_1014),
.B(n_1015),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1005),
.A2(n_1034),
.B1(n_1040),
.B2(n_1021),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1069),
.A2(n_1093),
.B(n_1075),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_960),
.Y(n_1113)
);

INVx8_ASAP7_75t_L g1114 ( 
.A(n_1014),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_L g1115 ( 
.A(n_1096),
.B(n_1002),
.C(n_1095),
.Y(n_1115)
);

AO32x2_ASAP7_75t_L g1116 ( 
.A1(n_1086),
.A2(n_1062),
.A3(n_1092),
.B1(n_1076),
.B2(n_962),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1103),
.B(n_963),
.Y(n_1117)
);

CKINVDCx16_ASAP7_75t_R g1118 ( 
.A(n_988),
.Y(n_1118)
);

OAI22x1_ASAP7_75t_L g1119 ( 
.A1(n_995),
.A2(n_1039),
.B1(n_1042),
.B2(n_1013),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_SL g1120 ( 
.A1(n_1024),
.A2(n_1053),
.B(n_1028),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_970),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1043),
.A2(n_969),
.B(n_1050),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1044),
.A2(n_1013),
.B1(n_996),
.B2(n_959),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_965),
.B(n_972),
.Y(n_1124)
);

NOR2x1_ASAP7_75t_L g1125 ( 
.A(n_1052),
.B(n_1010),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1049),
.A2(n_976),
.B(n_1055),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_1035),
.B(n_1102),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_982),
.A2(n_974),
.B(n_981),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_987),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1080),
.A2(n_1068),
.B(n_1090),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1055),
.A2(n_1070),
.B(n_1045),
.Y(n_1131)
);

AOI221x1_ASAP7_75t_L g1132 ( 
.A1(n_983),
.A2(n_990),
.B1(n_1006),
.B2(n_1023),
.C(n_1038),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_1052),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_994),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1045),
.A2(n_1060),
.B(n_961),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1053),
.A2(n_1074),
.B(n_979),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1102),
.B(n_1027),
.Y(n_1137)
);

BUFx10_ASAP7_75t_L g1138 ( 
.A(n_1058),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_986),
.B(n_1011),
.C(n_1056),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1066),
.A2(n_1074),
.B(n_1088),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1066),
.A2(n_1091),
.B(n_1071),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_SL g1142 ( 
.A1(n_1048),
.A2(n_1026),
.B(n_1009),
.C(n_1032),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_964),
.A2(n_1064),
.B(n_1057),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_1087),
.A2(n_1078),
.B(n_1089),
.Y(n_1144)
);

NAND3xp33_ASAP7_75t_L g1145 ( 
.A(n_986),
.B(n_1011),
.C(n_1056),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_1004),
.A2(n_1083),
.A3(n_1081),
.B(n_999),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1057),
.A2(n_1019),
.B(n_1030),
.C(n_1008),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1019),
.A2(n_991),
.B(n_1020),
.C(n_1003),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_967),
.B(n_1029),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1077),
.A2(n_968),
.B(n_981),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_SL g1151 ( 
.A1(n_1036),
.A2(n_1089),
.B(n_1059),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_980),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_989),
.A2(n_998),
.B1(n_997),
.B2(n_1047),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1015),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1063),
.B(n_966),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_SL g1156 ( 
.A(n_985),
.B(n_1099),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_1046),
.A2(n_1017),
.A3(n_1079),
.B(n_1082),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_968),
.A2(n_1054),
.B(n_975),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_1061),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1063),
.B(n_1031),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1012),
.A2(n_1072),
.B(n_977),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_971),
.Y(n_1162)
);

NOR2xp67_ASAP7_75t_L g1163 ( 
.A(n_1022),
.B(n_1025),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_1033),
.B(n_1041),
.Y(n_1164)
);

AOI21x1_ASAP7_75t_L g1165 ( 
.A1(n_993),
.A2(n_1085),
.B(n_1001),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_991),
.A2(n_1020),
.B(n_1073),
.C(n_1065),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_1018),
.A2(n_1101),
.A3(n_1037),
.B(n_978),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_985),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1104),
.A2(n_1000),
.B(n_1022),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1025),
.B(n_1104),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1084),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1084),
.A2(n_1096),
.B(n_1005),
.C(n_613),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1084),
.A2(n_1086),
.A3(n_1090),
.B(n_1093),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1007),
.A2(n_1095),
.B1(n_613),
.B2(n_1096),
.Y(n_1174)
);

OAI22x1_ASAP7_75t_L g1175 ( 
.A1(n_1007),
.A2(n_1005),
.B1(n_481),
.B2(n_480),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1097),
.B(n_333),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_SL g1177 ( 
.A1(n_1024),
.A2(n_1053),
.B(n_1028),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_982),
.A2(n_936),
.B(n_1075),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_982),
.A2(n_936),
.B(n_1075),
.Y(n_1179)
);

INVx5_ASAP7_75t_L g1180 ( 
.A(n_994),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1095),
.B(n_613),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_973),
.A2(n_1016),
.B(n_835),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_973),
.A2(n_1016),
.B(n_835),
.Y(n_1183)
);

NAND3xp33_ASAP7_75t_SL g1184 ( 
.A(n_1005),
.B(n_457),
.C(n_448),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_1005),
.B(n_1096),
.C(n_818),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1095),
.B(n_613),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_973),
.A2(n_1016),
.B(n_835),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_960),
.Y(n_1188)
);

NOR2xp67_ASAP7_75t_SL g1189 ( 
.A(n_988),
.B(n_448),
.Y(n_1189)
);

OR2x6_ASAP7_75t_L g1190 ( 
.A(n_1014),
.B(n_794),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_973),
.A2(n_1016),
.B(n_835),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1096),
.A2(n_1005),
.B(n_613),
.C(n_1002),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_973),
.A2(n_1016),
.B(n_835),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1097),
.B(n_333),
.Y(n_1194)
);

OAI22x1_ASAP7_75t_L g1195 ( 
.A1(n_1005),
.A2(n_481),
.B1(n_480),
.B2(n_1034),
.Y(n_1195)
);

OAI21xp33_ASAP7_75t_L g1196 ( 
.A1(n_1005),
.A2(n_481),
.B(n_634),
.Y(n_1196)
);

AOI221x1_ASAP7_75t_L g1197 ( 
.A1(n_1002),
.A2(n_973),
.B1(n_1096),
.B2(n_1005),
.C(n_1028),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1097),
.B(n_333),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_982),
.A2(n_936),
.B(n_1075),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1005),
.A2(n_1096),
.B(n_613),
.C(n_606),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1096),
.A2(n_613),
.B(n_1095),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_982),
.A2(n_936),
.B(n_1075),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_982),
.A2(n_936),
.B(n_1075),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1095),
.B(n_613),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_960),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_973),
.A2(n_1016),
.B(n_835),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1095),
.B(n_613),
.Y(n_1207)
);

AO32x2_ASAP7_75t_L g1208 ( 
.A1(n_1086),
.A2(n_1062),
.A3(n_1092),
.B1(n_876),
.B2(n_1076),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_SL g1209 ( 
.A1(n_1096),
.A2(n_1002),
.B(n_1048),
.C(n_990),
.Y(n_1209)
);

CKINVDCx11_ASAP7_75t_R g1210 ( 
.A(n_988),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_994),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_973),
.A2(n_1016),
.B(n_835),
.Y(n_1212)
);

AO32x2_ASAP7_75t_L g1213 ( 
.A1(n_1086),
.A2(n_1062),
.A3(n_1092),
.B1(n_876),
.B2(n_1076),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1039),
.A2(n_608),
.B1(n_340),
.B2(n_359),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1096),
.A2(n_613),
.B(n_1095),
.Y(n_1215)
);

AO32x2_ASAP7_75t_L g1216 ( 
.A1(n_1086),
.A2(n_1062),
.A3(n_1092),
.B1(n_876),
.B2(n_1076),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_960),
.Y(n_1217)
);

OAI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1095),
.A2(n_481),
.B1(n_811),
.B2(n_807),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_973),
.A2(n_1016),
.B(n_835),
.Y(n_1219)
);

INVxp67_ASAP7_75t_SL g1220 ( 
.A(n_1044),
.Y(n_1220)
);

NOR2xp67_ASAP7_75t_SL g1221 ( 
.A(n_988),
.B(n_448),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1096),
.A2(n_613),
.B(n_1095),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1096),
.A2(n_613),
.B(n_1095),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_973),
.A2(n_1016),
.B(n_835),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1095),
.B(n_613),
.Y(n_1225)
);

NAND3xp33_ASAP7_75t_L g1226 ( 
.A(n_1005),
.B(n_1096),
.C(n_818),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1095),
.B(n_613),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_973),
.A2(n_1016),
.B(n_835),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1096),
.A2(n_613),
.B(n_1095),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1086),
.A2(n_1090),
.A3(n_1093),
.B(n_1002),
.Y(n_1230)
);

OAI22x1_ASAP7_75t_L g1231 ( 
.A1(n_1005),
.A2(n_481),
.B1(n_480),
.B2(n_1034),
.Y(n_1231)
);

OA21x2_ASAP7_75t_L g1232 ( 
.A1(n_1006),
.A2(n_1090),
.B(n_983),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1097),
.B(n_1100),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_982),
.A2(n_936),
.B(n_1075),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_982),
.A2(n_936),
.B(n_1075),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_982),
.A2(n_936),
.B(n_1075),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_973),
.A2(n_1016),
.B(n_835),
.Y(n_1237)
);

OA21x2_ASAP7_75t_L g1238 ( 
.A1(n_1006),
.A2(n_1090),
.B(n_983),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1097),
.B(n_1100),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_973),
.A2(n_1016),
.B(n_835),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1107),
.Y(n_1241)
);

INVx6_ASAP7_75t_L g1242 ( 
.A(n_1180),
.Y(n_1242)
);

BUFx4f_ASAP7_75t_SL g1243 ( 
.A(n_1108),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1196),
.A2(n_1204),
.B1(n_1186),
.B2(n_1181),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1185),
.A2(n_1226),
.B1(n_1184),
.B2(n_1195),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1180),
.B(n_1133),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1231),
.A2(n_1156),
.B1(n_1214),
.B2(n_1225),
.Y(n_1247)
);

INVx6_ASAP7_75t_L g1248 ( 
.A(n_1114),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1207),
.B(n_1227),
.Y(n_1249)
);

INVx6_ASAP7_75t_L g1250 ( 
.A(n_1114),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1154),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1154),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1176),
.A2(n_1198),
.B1(n_1194),
.B2(n_1175),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1139),
.A2(n_1145),
.B1(n_1192),
.B2(n_1131),
.Y(n_1254)
);

BUFx8_ASAP7_75t_L g1255 ( 
.A(n_1154),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1124),
.A2(n_1233),
.B1(n_1239),
.B2(n_1119),
.Y(n_1256)
);

INVx6_ASAP7_75t_L g1257 ( 
.A(n_1110),
.Y(n_1257)
);

CKINVDCx11_ASAP7_75t_R g1258 ( 
.A(n_1210),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1121),
.Y(n_1259)
);

BUFx8_ASAP7_75t_L g1260 ( 
.A(n_1129),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1218),
.A2(n_1109),
.B1(n_1111),
.B2(n_1152),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1110),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1188),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1115),
.A2(n_1177),
.B1(n_1120),
.B2(n_1222),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1201),
.B(n_1215),
.Y(n_1265)
);

AOI22x1_ASAP7_75t_SL g1266 ( 
.A1(n_1168),
.A2(n_1105),
.B1(n_1220),
.B2(n_1217),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_1118),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1232),
.A2(n_1238),
.B1(n_1126),
.B2(n_1229),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1223),
.A2(n_1123),
.B1(n_1137),
.B2(n_1232),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1188),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1205),
.Y(n_1271)
);

BUFx12f_ASAP7_75t_L g1272 ( 
.A(n_1138),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1238),
.A2(n_1135),
.B1(n_1136),
.B2(n_1141),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1205),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1118),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1117),
.A2(n_1174),
.B1(n_1143),
.B2(n_1127),
.Y(n_1276)
);

BUFx2_ASAP7_75t_SL g1277 ( 
.A(n_1134),
.Y(n_1277)
);

INVx4_ASAP7_75t_L g1278 ( 
.A(n_1134),
.Y(n_1278)
);

CKINVDCx11_ASAP7_75t_R g1279 ( 
.A(n_1138),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1182),
.A2(n_1240),
.B1(n_1187),
.B2(n_1183),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1153),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1191),
.A2(n_1237),
.B1(n_1228),
.B2(n_1224),
.Y(n_1282)
);

OAI21xp33_ASAP7_75t_L g1283 ( 
.A1(n_1200),
.A2(n_1172),
.B(n_1147),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1155),
.B(n_1149),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1189),
.A2(n_1221),
.B1(n_1193),
.B2(n_1212),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1190),
.Y(n_1286)
);

INVx6_ASAP7_75t_L g1287 ( 
.A(n_1171),
.Y(n_1287)
);

CKINVDCx6p67_ASAP7_75t_R g1288 ( 
.A(n_1211),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1206),
.A2(n_1219),
.B1(n_1160),
.B2(n_1162),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1159),
.A2(n_1130),
.B1(n_1164),
.B2(n_1140),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1158),
.A2(n_1169),
.B1(n_1161),
.B2(n_1144),
.Y(n_1291)
);

INVx6_ASAP7_75t_L g1292 ( 
.A(n_1211),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1167),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_1125),
.Y(n_1294)
);

BUFx4f_ASAP7_75t_SL g1295 ( 
.A(n_1133),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1197),
.B(n_1150),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1148),
.A2(n_1112),
.B1(n_1166),
.B2(n_1144),
.Y(n_1297)
);

BUFx8_ASAP7_75t_SL g1298 ( 
.A(n_1165),
.Y(n_1298)
);

BUFx4_ASAP7_75t_R g1299 ( 
.A(n_1163),
.Y(n_1299)
);

INVx4_ASAP7_75t_L g1300 ( 
.A(n_1170),
.Y(n_1300)
);

INVx3_ASAP7_75t_L g1301 ( 
.A(n_1173),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1173),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1132),
.A2(n_1106),
.B(n_1122),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1151),
.Y(n_1304)
);

CKINVDCx11_ASAP7_75t_R g1305 ( 
.A(n_1142),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1209),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1230),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1128),
.A2(n_1236),
.B1(n_1235),
.B2(n_1234),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1230),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1157),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1178),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1116),
.A2(n_1216),
.B1(n_1213),
.B2(n_1208),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1116),
.A2(n_1216),
.B1(n_1213),
.B2(n_1208),
.Y(n_1313)
);

OAI22x1_ASAP7_75t_L g1314 ( 
.A1(n_1116),
.A2(n_1216),
.B1(n_1213),
.B2(n_1208),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1146),
.A2(n_1179),
.B1(n_1199),
.B2(n_1202),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1203),
.A2(n_925),
.B1(n_1145),
.B2(n_1139),
.Y(n_1316)
);

INVx4_ASAP7_75t_L g1317 ( 
.A(n_1180),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1196),
.A2(n_1095),
.B1(n_1186),
.B2(n_1181),
.Y(n_1318)
);

CKINVDCx11_ASAP7_75t_R g1319 ( 
.A(n_1107),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1129),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1181),
.B(n_1186),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1196),
.A2(n_1095),
.B1(n_1186),
.B2(n_1181),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_SL g1323 ( 
.A1(n_1195),
.A2(n_1231),
.B1(n_1175),
.B2(n_1005),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1185),
.A2(n_1005),
.B1(n_1226),
.B2(n_673),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1181),
.B(n_1186),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1196),
.A2(n_1095),
.B1(n_1186),
.B2(n_1181),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1196),
.A2(n_1176),
.B1(n_1198),
.B2(n_1194),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1196),
.A2(n_1226),
.B1(n_1185),
.B2(n_1184),
.Y(n_1328)
);

INVx4_ASAP7_75t_SL g1329 ( 
.A(n_1171),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1196),
.A2(n_1226),
.B1(n_1185),
.B2(n_1184),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1196),
.A2(n_1226),
.B1(n_1185),
.B2(n_1184),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1105),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1113),
.Y(n_1333)
);

CKINVDCx11_ASAP7_75t_R g1334 ( 
.A(n_1107),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1113),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_SL g1336 ( 
.A(n_1190),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1180),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1196),
.A2(n_1226),
.B1(n_1185),
.B2(n_1184),
.Y(n_1338)
);

CKINVDCx11_ASAP7_75t_R g1339 ( 
.A(n_1107),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1196),
.A2(n_1095),
.B1(n_1186),
.B2(n_1181),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1196),
.A2(n_1095),
.B1(n_1186),
.B2(n_1181),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1129),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1196),
.A2(n_1176),
.B1(n_1198),
.B2(n_1194),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1310),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1293),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1254),
.A2(n_1324),
.B(n_1283),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1281),
.B(n_1302),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1315),
.A2(n_1308),
.B(n_1291),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1315),
.A2(n_1303),
.B(n_1297),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1309),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1298),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1301),
.A2(n_1296),
.B(n_1307),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1296),
.B(n_1254),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1319),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1259),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1328),
.A2(n_1330),
.B(n_1331),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1263),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1270),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1305),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1271),
.Y(n_1360)
);

NAND3xp33_ASAP7_75t_L g1361 ( 
.A(n_1338),
.B(n_1245),
.C(n_1276),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1274),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1332),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1333),
.B(n_1335),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1260),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1332),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1265),
.A2(n_1264),
.B(n_1285),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1284),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1327),
.A2(n_1343),
.B1(n_1253),
.B2(n_1247),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1273),
.B(n_1268),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1320),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1244),
.B(n_1318),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1269),
.B(n_1313),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1244),
.B(n_1249),
.Y(n_1374)
);

NAND2x1_ASAP7_75t_L g1375 ( 
.A(n_1289),
.B(n_1290),
.Y(n_1375)
);

AO21x2_ASAP7_75t_L g1376 ( 
.A1(n_1312),
.A2(n_1256),
.B(n_1322),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1314),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1311),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1342),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1249),
.B(n_1321),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1261),
.A2(n_1306),
.B1(n_1325),
.B2(n_1321),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1280),
.Y(n_1382)
);

NOR2x1_ASAP7_75t_R g1383 ( 
.A(n_1258),
.B(n_1275),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1242),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1282),
.Y(n_1385)
);

AO21x2_ASAP7_75t_L g1386 ( 
.A1(n_1318),
.A2(n_1341),
.B(n_1322),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1300),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1326),
.A2(n_1341),
.B(n_1340),
.Y(n_1388)
);

AO21x2_ASAP7_75t_L g1389 ( 
.A1(n_1326),
.A2(n_1340),
.B(n_1325),
.Y(n_1389)
);

AO21x2_ASAP7_75t_L g1390 ( 
.A1(n_1316),
.A2(n_1304),
.B(n_1323),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1246),
.A2(n_1337),
.B(n_1317),
.Y(n_1391)
);

AOI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1294),
.A2(n_1299),
.B(n_1266),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1257),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1337),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1336),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1334),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1286),
.Y(n_1397)
);

BUFx2_ASAP7_75t_SL g1398 ( 
.A(n_1336),
.Y(n_1398)
);

BUFx12f_ASAP7_75t_L g1399 ( 
.A(n_1339),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1329),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1329),
.Y(n_1401)
);

INVx4_ASAP7_75t_SL g1402 ( 
.A(n_1295),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1272),
.A2(n_1279),
.B1(n_1260),
.B2(n_1267),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1262),
.B(n_1277),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1288),
.A2(n_1292),
.B(n_1241),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1344),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1344),
.Y(n_1407)
);

AND2x2_ASAP7_75t_SL g1408 ( 
.A(n_1370),
.B(n_1278),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1345),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1369),
.A2(n_1361),
.B(n_1356),
.Y(n_1410)
);

INVx4_ASAP7_75t_L g1411 ( 
.A(n_1405),
.Y(n_1411)
);

NOR2x1_ASAP7_75t_SL g1412 ( 
.A(n_1386),
.B(n_1252),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1369),
.A2(n_1252),
.B(n_1251),
.C(n_1255),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1361),
.A2(n_1243),
.B(n_1287),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1377),
.B(n_1370),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1344),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1396),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1356),
.A2(n_1248),
.B1(n_1250),
.B2(n_1292),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1363),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1368),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1381),
.A2(n_1248),
.B1(n_1250),
.B2(n_1346),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1347),
.B(n_1373),
.Y(n_1422)
);

A2O1A1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1346),
.A2(n_1388),
.B(n_1375),
.C(n_1372),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1347),
.B(n_1373),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1396),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1347),
.B(n_1364),
.Y(n_1426)
);

AOI221xp5_ASAP7_75t_L g1427 ( 
.A1(n_1388),
.A2(n_1374),
.B1(n_1386),
.B2(n_1385),
.C(n_1382),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1371),
.B(n_1379),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1375),
.A2(n_1367),
.B(n_1374),
.C(n_1385),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1364),
.B(n_1355),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1353),
.B(n_1378),
.Y(n_1431)
);

INVx5_ASAP7_75t_SL g1432 ( 
.A(n_1386),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1353),
.B(n_1378),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1364),
.B(n_1355),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1357),
.B(n_1360),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1357),
.B(n_1360),
.Y(n_1436)
);

NOR2x1_ASAP7_75t_SL g1437 ( 
.A(n_1386),
.B(n_1389),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1366),
.Y(n_1438)
);

NOR2x1_ASAP7_75t_R g1439 ( 
.A(n_1396),
.B(n_1399),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1382),
.A2(n_1389),
.B(n_1380),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1390),
.A2(n_1380),
.B(n_1387),
.C(n_1351),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1405),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1390),
.A2(n_1351),
.B1(n_1376),
.B2(n_1389),
.Y(n_1443)
);

NAND2xp33_ASAP7_75t_L g1444 ( 
.A(n_1359),
.B(n_1397),
.Y(n_1444)
);

OR2x2_ASAP7_75t_SL g1445 ( 
.A(n_1405),
.B(n_1397),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1351),
.A2(n_1359),
.B1(n_1397),
.B2(n_1399),
.Y(n_1446)
);

OAI21xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1367),
.A2(n_1349),
.B(n_1358),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1399),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1431),
.B(n_1349),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1406),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1430),
.B(n_1434),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1440),
.B(n_1389),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1407),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1434),
.B(n_1348),
.Y(n_1454)
);

NAND2x1_ASAP7_75t_L g1455 ( 
.A(n_1411),
.B(n_1405),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1442),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1415),
.B(n_1352),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1415),
.B(n_1352),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1432),
.B(n_1416),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1427),
.B(n_1376),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1442),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1433),
.B(n_1376),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1445),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1423),
.A2(n_1359),
.B1(n_1392),
.B2(n_1398),
.Y(n_1464)
);

INVxp67_ASAP7_75t_SL g1465 ( 
.A(n_1433),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1426),
.B(n_1350),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1410),
.A2(n_1376),
.B1(n_1390),
.B2(n_1359),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1420),
.B(n_1362),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1409),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1409),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1435),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1464),
.B(n_1419),
.Y(n_1472)
);

OR2x6_ASAP7_75t_L g1473 ( 
.A(n_1455),
.B(n_1441),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1469),
.Y(n_1474)
);

NAND4xp25_ASAP7_75t_L g1475 ( 
.A(n_1467),
.B(n_1460),
.C(n_1443),
.D(n_1464),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1454),
.B(n_1432),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1456),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1469),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1465),
.B(n_1438),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1469),
.Y(n_1480)
);

AO21x2_ASAP7_75t_L g1481 ( 
.A1(n_1452),
.A2(n_1437),
.B(n_1412),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1462),
.B(n_1432),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1470),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1450),
.Y(n_1484)
);

NOR3xp33_ASAP7_75t_L g1485 ( 
.A(n_1460),
.B(n_1414),
.C(n_1429),
.Y(n_1485)
);

OAI31xp33_ASAP7_75t_L g1486 ( 
.A1(n_1467),
.A2(n_1446),
.A3(n_1413),
.B(n_1395),
.Y(n_1486)
);

AO21x2_ASAP7_75t_L g1487 ( 
.A1(n_1452),
.A2(n_1437),
.B(n_1412),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_L g1488 ( 
.A(n_1462),
.B(n_1421),
.C(n_1444),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1468),
.B(n_1371),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1459),
.B(n_1411),
.Y(n_1490)
);

INVx4_ASAP7_75t_L g1491 ( 
.A(n_1463),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1454),
.B(n_1432),
.Y(n_1492)
);

OAI222xp33_ASAP7_75t_L g1493 ( 
.A1(n_1463),
.A2(n_1421),
.B1(n_1392),
.B2(n_1418),
.C1(n_1424),
.C2(n_1422),
.Y(n_1493)
);

NAND2x1p5_ASAP7_75t_L g1494 ( 
.A(n_1455),
.B(n_1442),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1456),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1449),
.B(n_1432),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1454),
.B(n_1422),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1453),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1465),
.B(n_1435),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1468),
.B(n_1436),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1456),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1489),
.B(n_1466),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1484),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1497),
.B(n_1463),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1489),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1474),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1482),
.B(n_1449),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1497),
.B(n_1463),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1485),
.B(n_1466),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1474),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1497),
.B(n_1451),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1491),
.B(n_1451),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1478),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_1472),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1491),
.B(n_1451),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1482),
.B(n_1449),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1478),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1480),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1479),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1480),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1485),
.B(n_1466),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1491),
.B(n_1461),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1484),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1482),
.B(n_1471),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1499),
.B(n_1471),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1472),
.B(n_1457),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1484),
.Y(n_1527)
);

OR2x6_ASAP7_75t_L g1528 ( 
.A(n_1491),
.B(n_1455),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1499),
.B(n_1471),
.Y(n_1529)
);

AND2x2_ASAP7_75t_SL g1530 ( 
.A(n_1491),
.B(n_1408),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1479),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1495),
.B(n_1461),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1476),
.B(n_1457),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1500),
.B(n_1496),
.Y(n_1534)
);

AND2x6_ASAP7_75t_SL g1535 ( 
.A(n_1473),
.B(n_1439),
.Y(n_1535)
);

NOR2x1_ASAP7_75t_L g1536 ( 
.A(n_1475),
.B(n_1461),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1476),
.B(n_1457),
.Y(n_1537)
);

INVxp67_ASAP7_75t_SL g1538 ( 
.A(n_1495),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1514),
.B(n_1424),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1506),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1506),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1509),
.B(n_1458),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1510),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1510),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1513),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1523),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1513),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1534),
.B(n_1496),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1504),
.B(n_1476),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1521),
.B(n_1458),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1519),
.B(n_1458),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1523),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1517),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1534),
.B(n_1496),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1517),
.Y(n_1555)
);

INVx3_ASAP7_75t_SL g1556 ( 
.A(n_1530),
.Y(n_1556)
);

OAI32xp33_ASAP7_75t_L g1557 ( 
.A1(n_1536),
.A2(n_1475),
.A3(n_1488),
.B1(n_1477),
.B2(n_1447),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1518),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1504),
.B(n_1492),
.Y(n_1559)
);

NOR2xp67_ASAP7_75t_SL g1560 ( 
.A(n_1505),
.B(n_1397),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1523),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1518),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1508),
.B(n_1492),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1520),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1520),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1531),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1527),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1538),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1522),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1536),
.B(n_1488),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1527),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1527),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1503),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1526),
.B(n_1502),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1503),
.Y(n_1575)
);

INVxp33_ASAP7_75t_L g1576 ( 
.A(n_1512),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1525),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1530),
.A2(n_1486),
.B1(n_1390),
.B2(n_1408),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1524),
.B(n_1483),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1508),
.B(n_1492),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1556),
.B(n_1522),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1568),
.B(n_1507),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1570),
.B(n_1512),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1556),
.B(n_1522),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1556),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1546),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1566),
.B(n_1507),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1546),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1580),
.B(n_1522),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1543),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1539),
.B(n_1439),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1543),
.Y(n_1592)
);

AOI221xp5_ASAP7_75t_L g1593 ( 
.A1(n_1557),
.A2(n_1493),
.B1(n_1486),
.B2(n_1516),
.C(n_1446),
.Y(n_1593)
);

NOR2x1_ASAP7_75t_L g1594 ( 
.A(n_1540),
.B(n_1354),
.Y(n_1594)
);

AOI211x1_ASAP7_75t_SL g1595 ( 
.A1(n_1557),
.A2(n_1535),
.B(n_1359),
.C(n_1397),
.Y(n_1595)
);

INVxp67_ASAP7_75t_L g1596 ( 
.A(n_1560),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1549),
.B(n_1515),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1544),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1580),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1544),
.Y(n_1600)
);

AOI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1578),
.A2(n_1493),
.B1(n_1516),
.B2(n_1428),
.C(n_1515),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1574),
.B(n_1511),
.Y(n_1602)
);

NOR3xp33_ASAP7_75t_L g1603 ( 
.A(n_1569),
.B(n_1383),
.C(n_1395),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1548),
.B(n_1524),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1552),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1577),
.B(n_1511),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1545),
.Y(n_1607)
);

AOI31xp33_ASAP7_75t_L g1608 ( 
.A1(n_1576),
.A2(n_1383),
.A3(n_1425),
.B(n_1417),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1580),
.B(n_1530),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1545),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1569),
.B(n_1528),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1549),
.B(n_1533),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1547),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1547),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1577),
.B(n_1533),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_SL g1616 ( 
.A1(n_1595),
.A2(n_1403),
.B(n_1359),
.Y(n_1616)
);

NAND2xp33_ASAP7_75t_SL g1617 ( 
.A(n_1581),
.B(n_1560),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1590),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1585),
.B(n_1559),
.Y(n_1619)
);

AOI332xp33_ASAP7_75t_L g1620 ( 
.A1(n_1590),
.A2(n_1555),
.A3(n_1558),
.B1(n_1553),
.B2(n_1541),
.B3(n_1564),
.C1(n_1565),
.C2(n_1562),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1599),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1594),
.A2(n_1473),
.B(n_1448),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1583),
.B(n_1548),
.Y(n_1623)
);

OAI32xp33_ASAP7_75t_L g1624 ( 
.A1(n_1609),
.A2(n_1554),
.A3(n_1477),
.B1(n_1494),
.B2(n_1550),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1601),
.B(n_1593),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1592),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1592),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_R g1628 ( 
.A(n_1599),
.B(n_1397),
.Y(n_1628)
);

OAI32xp33_ASAP7_75t_L g1629 ( 
.A1(n_1599),
.A2(n_1554),
.A3(n_1494),
.B1(n_1542),
.B2(n_1501),
.Y(n_1629)
);

OAI21xp33_ASAP7_75t_SL g1630 ( 
.A1(n_1581),
.A2(n_1563),
.B(n_1559),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1598),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1612),
.B(n_1563),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1612),
.B(n_1537),
.Y(n_1633)
);

AOI221x1_ASAP7_75t_L g1634 ( 
.A1(n_1603),
.A2(n_1553),
.B1(n_1558),
.B2(n_1555),
.C(n_1573),
.Y(n_1634)
);

OAI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1596),
.A2(n_1608),
.B1(n_1473),
.B2(n_1582),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1602),
.B(n_1551),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1598),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1591),
.A2(n_1473),
.B1(n_1408),
.B2(n_1490),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1584),
.A2(n_1473),
.B(n_1494),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1597),
.B(n_1584),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1625),
.A2(n_1589),
.B1(n_1615),
.B2(n_1597),
.Y(n_1641)
);

NAND2xp33_ASAP7_75t_SL g1642 ( 
.A(n_1628),
.B(n_1582),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1618),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1619),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1617),
.A2(n_1589),
.B1(n_1606),
.B2(n_1473),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1640),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1622),
.A2(n_1589),
.B1(n_1587),
.B2(n_1445),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1621),
.B(n_1587),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1632),
.B(n_1604),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1626),
.Y(n_1650)
);

A2O1A1Ixp33_ASAP7_75t_L g1651 ( 
.A1(n_1622),
.A2(n_1611),
.B(n_1604),
.C(n_1535),
.Y(n_1651)
);

AOI32xp33_ASAP7_75t_L g1652 ( 
.A1(n_1635),
.A2(n_1611),
.A3(n_1610),
.B1(n_1607),
.B2(n_1600),
.Y(n_1652)
);

OA21x2_ASAP7_75t_L g1653 ( 
.A1(n_1634),
.A2(n_1614),
.B(n_1613),
.Y(n_1653)
);

OAI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1638),
.A2(n_1616),
.B1(n_1630),
.B2(n_1639),
.C(n_1623),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1627),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1631),
.B(n_1614),
.Y(n_1656)
);

INVxp33_ASAP7_75t_L g1657 ( 
.A(n_1636),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1637),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1635),
.A2(n_1613),
.B(n_1611),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1641),
.B(n_1637),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1658),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1653),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1651),
.A2(n_1633),
.B1(n_1528),
.B2(n_1532),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1646),
.B(n_1586),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1659),
.A2(n_1653),
.B(n_1642),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1648),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1657),
.B(n_1624),
.Y(n_1667)
);

AOI21xp33_ASAP7_75t_L g1668 ( 
.A1(n_1659),
.A2(n_1629),
.B(n_1588),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1644),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1647),
.A2(n_1528),
.B1(n_1481),
.B2(n_1487),
.Y(n_1670)
);

NOR3xp33_ASAP7_75t_L g1671 ( 
.A(n_1669),
.B(n_1654),
.C(n_1652),
.Y(n_1671)
);

NOR3xp33_ASAP7_75t_L g1672 ( 
.A(n_1665),
.B(n_1650),
.C(n_1643),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1662),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_SL g1674 ( 
.A(n_1661),
.B(n_1649),
.Y(n_1674)
);

NOR4xp25_ASAP7_75t_L g1675 ( 
.A(n_1660),
.B(n_1655),
.C(n_1656),
.D(n_1645),
.Y(n_1675)
);

NAND3xp33_ASAP7_75t_L g1676 ( 
.A(n_1665),
.B(n_1620),
.C(n_1588),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_SL g1677 ( 
.A(n_1667),
.B(n_1379),
.C(n_1586),
.Y(n_1677)
);

NAND4xp75_ASAP7_75t_L g1678 ( 
.A(n_1668),
.B(n_1605),
.C(n_1572),
.D(n_1567),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1663),
.B(n_1605),
.Y(n_1679)
);

OAI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1676),
.A2(n_1666),
.B(n_1664),
.C(n_1670),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1674),
.B(n_1365),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1678),
.A2(n_1671),
.B1(n_1673),
.B2(n_1672),
.Y(n_1682)
);

AOI211xp5_ASAP7_75t_SL g1683 ( 
.A1(n_1677),
.A2(n_1395),
.B(n_1572),
.C(n_1567),
.Y(n_1683)
);

AOI211xp5_ASAP7_75t_SL g1684 ( 
.A1(n_1675),
.A2(n_1395),
.B(n_1573),
.C(n_1404),
.Y(n_1684)
);

AOI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1682),
.A2(n_1679),
.B1(n_1552),
.B2(n_1561),
.C(n_1571),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1681),
.A2(n_1528),
.B1(n_1398),
.B2(n_1365),
.Y(n_1686)
);

AOI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1680),
.A2(n_1365),
.B(n_1404),
.C(n_1571),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1683),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1684),
.A2(n_1561),
.B1(n_1575),
.B2(n_1532),
.C(n_1501),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1682),
.A2(n_1575),
.B1(n_1532),
.B2(n_1495),
.C(n_1501),
.Y(n_1690)
);

NAND4xp75_ASAP7_75t_L g1691 ( 
.A(n_1690),
.B(n_1391),
.C(n_1384),
.D(n_1418),
.Y(n_1691)
);

NAND4xp75_ASAP7_75t_L g1692 ( 
.A(n_1685),
.B(n_1391),
.C(n_1384),
.D(n_1400),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1688),
.Y(n_1693)
);

NAND2x1p5_ASAP7_75t_SL g1694 ( 
.A(n_1687),
.B(n_1402),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1686),
.Y(n_1695)
);

AOI222xp33_ASAP7_75t_L g1696 ( 
.A1(n_1693),
.A2(n_1689),
.B1(n_1532),
.B2(n_1402),
.C1(n_1537),
.C2(n_1447),
.Y(n_1696)
);

INVx4_ASAP7_75t_L g1697 ( 
.A(n_1695),
.Y(n_1697)
);

O2A1O1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1694),
.A2(n_1528),
.B(n_1579),
.C(n_1494),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_1697),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1699),
.Y(n_1700)
);

XNOR2xp5_ASAP7_75t_L g1701 ( 
.A(n_1700),
.B(n_1691),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1700),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1702),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1701),
.B(n_1691),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_SL g1705 ( 
.A1(n_1703),
.A2(n_1704),
.B(n_1698),
.Y(n_1705)
);

AO21x2_ASAP7_75t_L g1706 ( 
.A1(n_1703),
.A2(n_1692),
.B(n_1696),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1706),
.B(n_1579),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1707),
.A2(n_1705),
.B1(n_1529),
.B2(n_1525),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1708),
.Y(n_1709)
);

AOI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1709),
.A2(n_1394),
.B1(n_1490),
.B2(n_1393),
.C(n_1498),
.Y(n_1710)
);

AOI211xp5_ASAP7_75t_L g1711 ( 
.A1(n_1710),
.A2(n_1394),
.B(n_1401),
.C(n_1400),
.Y(n_1711)
);


endmodule