module real_aes_3689_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_1067;
wire n_518;
wire n_673;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_1034;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_666;
wire n_537;
wire n_320;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_1021;
wire n_700;
wire n_1046;
wire n_677;
wire n_948;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_892;
wire n_370;
wire n_994;
wire n_744;
wire n_384;
wire n_938;
wire n_352;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_455;
wire n_725;
wire n_973;
wire n_671;
wire n_960;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_1100;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1103;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_999;
wire n_913;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_713;
wire n_598;
wire n_756;
wire n_1073;
wire n_404;
wire n_728;
wire n_334;
wire n_735;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_1056;
wire n_358;
wire n_385;
wire n_397;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_1043;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_314;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_359;
wire n_1090;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_1101;
wire n_601;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_1104;
wire n_842;
wire n_1061;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_0), .A2(n_3), .B1(n_788), .B2(n_789), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_1), .A2(n_165), .B1(n_459), .B2(n_460), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_2), .A2(n_126), .B1(n_473), .B2(n_474), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_4), .A2(n_139), .B1(n_522), .B2(n_523), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_5), .A2(n_268), .B1(n_553), .B2(n_556), .Y(n_632) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_6), .A2(n_213), .B1(n_408), .B2(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_7), .A2(n_142), .B1(n_416), .B2(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g1094 ( .A(n_8), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_9), .A2(n_181), .B1(n_564), .B2(n_1056), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_10), .A2(n_280), .B1(n_522), .B2(n_564), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_11), .A2(n_255), .B1(n_436), .B2(n_490), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_12), .A2(n_24), .B1(n_430), .B2(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_13), .B(n_343), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_14), .A2(n_218), .B1(n_792), .B2(n_793), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_15), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_16), .A2(n_204), .B1(n_473), .B2(n_474), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_17), .A2(n_144), .B1(n_408), .B2(n_412), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_18), .A2(n_174), .B1(n_464), .B2(n_465), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_19), .B(n_664), .Y(n_663) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_20), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_21), .A2(n_224), .B1(n_843), .B2(n_845), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_22), .A2(n_64), .B1(n_364), .B2(n_373), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_23), .A2(n_125), .B1(n_405), .B2(n_570), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_25), .A2(n_169), .B1(n_843), .B2(n_845), .Y(n_842) );
AOI21xp33_ASAP7_75t_L g1066 ( .A1(n_26), .A2(n_580), .B(n_1067), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_27), .A2(n_187), .B1(n_492), .B2(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g647 ( .A(n_28), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_28), .A2(n_293), .B1(n_847), .B2(n_864), .Y(n_875) );
INVx1_ASAP7_75t_L g703 ( .A(n_29), .Y(n_703) );
INVxp33_ASAP7_75t_SL g865 ( .A(n_30), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_31), .A2(n_177), .B1(n_836), .B2(n_838), .Y(n_913) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_32), .A2(n_438), .B(n_748), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_33), .A2(n_46), .B1(n_828), .B2(n_833), .Y(n_914) );
INVx1_ASAP7_75t_L g749 ( .A(n_34), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_35), .A2(n_83), .B1(n_457), .B2(n_465), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_36), .A2(n_173), .B1(n_427), .B2(n_430), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_37), .A2(n_309), .B1(n_464), .B2(n_465), .Y(n_729) );
XOR2x2_ASAP7_75t_L g445 ( .A(n_38), .B(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_39), .A2(n_45), .B1(n_427), .B2(n_430), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g1057 ( .A1(n_40), .A2(n_44), .B1(n_502), .B2(n_1058), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_41), .A2(n_91), .B1(n_489), .B2(n_490), .Y(n_529) );
INVx1_ASAP7_75t_L g774 ( .A(n_42), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_43), .A2(n_113), .B1(n_489), .B2(n_490), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_47), .A2(n_151), .B1(n_507), .B2(n_744), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_48), .A2(n_88), .B1(n_473), .B2(n_474), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_49), .A2(n_160), .B1(n_408), .B2(n_612), .Y(n_694) );
OA22x2_ASAP7_75t_L g348 ( .A1(n_50), .A2(n_137), .B1(n_343), .B2(n_347), .Y(n_348) );
INVx1_ASAP7_75t_L g370 ( .A(n_50), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_51), .A2(n_262), .B1(n_570), .B2(n_767), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_52), .A2(n_239), .B1(n_847), .B2(n_848), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_53), .A2(n_56), .B1(n_473), .B2(n_474), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_54), .A2(n_102), .B1(n_440), .B2(n_490), .Y(n_1064) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_55), .A2(n_250), .B1(n_459), .B2(n_460), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_57), .A2(n_296), .B1(n_574), .B2(n_575), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_58), .A2(n_209), .B1(n_470), .B2(n_471), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_59), .A2(n_254), .B1(n_473), .B2(n_474), .Y(n_681) );
INVx1_ASAP7_75t_L g953 ( .A(n_60), .Y(n_953) );
AOI22xp5_ASAP7_75t_L g1060 ( .A1(n_61), .A2(n_188), .B1(n_428), .B2(n_1061), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_62), .A2(n_87), .B1(n_459), .B2(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_63), .A2(n_216), .B1(n_464), .B2(n_465), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_65), .A2(n_157), .B1(n_448), .B2(n_450), .C(n_452), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_66), .B(n_153), .Y(n_322) );
INVx1_ASAP7_75t_L g346 ( .A(n_66), .Y(n_346) );
OAI21xp33_ASAP7_75t_L g371 ( .A1(n_66), .A2(n_137), .B(n_372), .Y(n_371) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_67), .A2(n_492), .B(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_68), .A2(n_251), .B1(n_468), .B2(n_470), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_69), .A2(n_121), .B1(n_398), .B2(n_405), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_70), .A2(n_231), .B1(n_408), .B2(n_612), .Y(n_654) );
INVx1_ASAP7_75t_L g677 ( .A(n_71), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_72), .A2(n_155), .B1(n_398), .B2(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_73), .A2(n_127), .B1(n_379), .B2(n_389), .Y(n_378) );
AOI22xp33_ASAP7_75t_SL g655 ( .A1(n_74), .A2(n_179), .B1(n_398), .B2(n_405), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_75), .A2(n_279), .B1(n_364), .B2(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_76), .B(n_777), .Y(n_776) );
INVxp33_ASAP7_75t_L g857 ( .A(n_77), .Y(n_857) );
INVx1_ASAP7_75t_L g832 ( .A(n_78), .Y(n_832) );
AND2x4_ASAP7_75t_L g837 ( .A(n_78), .B(n_227), .Y(n_837) );
HB1xp67_ASAP7_75t_L g1103 ( .A(n_78), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_79), .A2(n_171), .B1(n_389), .B2(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g584 ( .A(n_80), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_81), .A2(n_82), .B1(n_618), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_84), .A2(n_163), .B1(n_440), .B2(n_471), .Y(n_725) );
INVx1_ASAP7_75t_L g810 ( .A(n_85), .Y(n_810) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_86), .A2(n_89), .B1(n_577), .B2(n_578), .C(n_581), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_90), .A2(n_467), .B(n_773), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_92), .A2(n_578), .B(n_722), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_93), .A2(n_269), .B1(n_467), .B2(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_94), .B(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_95), .A2(n_128), .B1(n_507), .B2(n_786), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_96), .A2(n_701), .B(n_702), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_97), .A2(n_129), .B1(n_504), .B2(n_525), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_98), .A2(n_123), .B1(n_615), .B2(n_616), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_99), .A2(n_152), .B1(n_468), .B2(n_471), .Y(n_674) );
INVx1_ASAP7_75t_L g582 ( .A(n_100), .Y(n_582) );
INVx1_ASAP7_75t_L g830 ( .A(n_101), .Y(n_830) );
AND2x4_ASAP7_75t_L g834 ( .A(n_101), .B(n_318), .Y(n_834) );
INVx1_ASAP7_75t_SL g844 ( .A(n_101), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_103), .A2(n_214), .B1(n_440), .B2(n_490), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_104), .A2(n_245), .B1(n_613), .B2(n_616), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g851 ( .A1(n_105), .A2(n_195), .B1(n_847), .B2(n_848), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_106), .A2(n_236), .B1(n_612), .B2(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g635 ( .A(n_107), .Y(n_635) );
INVx1_ASAP7_75t_L g538 ( .A(n_108), .Y(n_538) );
XOR2xp5_ASAP7_75t_L g1077 ( .A(n_109), .B(n_1078), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_110), .A2(n_220), .B1(n_504), .B2(n_505), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_111), .A2(n_285), .B1(n_416), .B2(n_744), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_112), .A2(n_295), .B1(n_467), .B2(n_470), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g1097 ( .A1(n_114), .A2(n_300), .B1(n_450), .B2(n_1098), .C(n_1099), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_115), .A2(n_230), .B1(n_836), .B2(n_838), .Y(n_835) );
XNOR2x1_ASAP7_75t_L g712 ( .A(n_116), .B(n_713), .Y(n_712) );
OAI22x1_ASAP7_75t_L g330 ( .A1(n_117), .A2(n_331), .B1(n_442), .B2(n_443), .Y(n_330) );
NAND3xp33_ASAP7_75t_SL g442 ( .A(n_117), .B(n_396), .C(n_433), .Y(n_442) );
INVx1_ASAP7_75t_L g719 ( .A(n_118), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_119), .A2(n_150), .B1(n_456), .B2(n_457), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_120), .A2(n_298), .B1(n_473), .B2(n_474), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_122), .A2(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g1088 ( .A(n_124), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_130), .B(n_701), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_131), .A2(n_308), .B1(n_828), .B2(n_833), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g1059 ( .A1(n_132), .A2(n_261), .B1(n_507), .B2(n_508), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_133), .A2(n_253), .B1(n_508), .B2(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g710 ( .A(n_134), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_135), .A2(n_288), .B1(n_464), .B2(n_465), .Y(n_630) );
INVx1_ASAP7_75t_L g360 ( .A(n_136), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_136), .B(n_182), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_136), .B(n_368), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_137), .B(n_238), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_138), .A2(n_146), .B1(n_843), .B2(n_845), .Y(n_850) );
INVx1_ASAP7_75t_L g1052 ( .A(n_138), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_138), .A2(n_1075), .B1(n_1077), .B2(n_1101), .Y(n_1074) );
INVx1_ASAP7_75t_L g661 ( .A(n_140), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_141), .A2(n_233), .B1(n_436), .B2(n_779), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_143), .A2(n_149), .B1(n_436), .B2(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_145), .A2(n_199), .B1(n_507), .B2(n_508), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_147), .A2(n_265), .B1(n_795), .B2(n_796), .Y(n_794) );
INVx1_ASAP7_75t_L g494 ( .A(n_148), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_153), .B(n_353), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_154), .A2(n_178), .B1(n_428), .B2(n_505), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_156), .A2(n_310), .B1(n_507), .B2(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g723 ( .A(n_158), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_159), .A2(n_205), .B1(n_362), .B2(n_373), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_161), .A2(n_252), .B1(n_504), .B2(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_162), .B(n_1091), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_164), .A2(n_290), .B1(n_436), .B2(n_485), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_166), .A2(n_513), .B1(n_514), .B2(n_540), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_166), .Y(n_513) );
INVx1_ASAP7_75t_L g1068 ( .A(n_167), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_168), .B(n_577), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_170), .A2(n_311), .B1(n_575), .B2(n_627), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_172), .A2(n_217), .B1(n_862), .B2(n_864), .Y(n_955) );
XNOR2x1_ASAP7_75t_L g763 ( .A(n_175), .B(n_764), .Y(n_763) );
AOI22xp33_ASAP7_75t_SL g846 ( .A1(n_175), .A2(n_229), .B1(n_847), .B2(n_848), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_176), .A2(n_301), .B1(n_802), .B2(n_803), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_180), .A2(n_287), .B1(n_428), .B2(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g344 ( .A(n_182), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g876 ( .A1(n_183), .A2(n_186), .B1(n_843), .B2(n_845), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_184), .A2(n_208), .B1(n_653), .B2(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_185), .B(n_335), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_189), .A2(n_207), .B1(n_651), .B2(n_696), .Y(n_695) );
XNOR2x1_ASAP7_75t_L g541 ( .A(n_190), .B(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_191), .A2(n_283), .B1(n_379), .B2(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_192), .A2(n_235), .B1(n_609), .B2(n_753), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_193), .A2(n_198), .B1(n_609), .B2(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_194), .B(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_196), .A2(n_272), .B1(n_502), .B2(n_564), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_197), .A2(n_248), .B1(n_408), .B2(n_566), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_200), .A2(n_215), .B1(n_456), .B2(n_457), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_201), .A2(n_264), .B1(n_398), .B2(n_519), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_202), .A2(n_247), .B1(n_553), .B2(n_556), .Y(n_1084) );
INVx1_ASAP7_75t_L g954 ( .A(n_203), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_206), .A2(n_266), .B1(n_492), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_210), .A2(n_242), .B1(n_470), .B2(n_471), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_211), .A2(n_243), .B1(n_428), .B2(n_505), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_212), .A2(n_294), .B1(n_519), .B2(n_1061), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_219), .B(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_221), .A2(n_304), .B1(n_598), .B2(n_600), .Y(n_597) );
AOI221xp5_ASAP7_75t_L g805 ( .A1(n_222), .A2(n_223), .B1(n_609), .B2(n_806), .C(n_809), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_225), .A2(n_256), .B1(n_456), .B2(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g1096 ( .A(n_226), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_227), .Y(n_323) );
AND2x4_ASAP7_75t_L g831 ( .A(n_227), .B(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_228), .B(n_532), .Y(n_531) );
XNOR2x2_ASAP7_75t_L g782 ( .A(n_230), .B(n_783), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_232), .A2(n_260), .B1(n_456), .B2(n_457), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_234), .A2(n_305), .B1(n_373), .B2(n_756), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_237), .A2(n_275), .B1(n_467), .B2(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g358 ( .A(n_238), .Y(n_358) );
INVxp67_ASAP7_75t_L g388 ( .A(n_238), .Y(n_388) );
INVx1_ASAP7_75t_L g453 ( .A(n_240), .Y(n_453) );
INVx1_ASAP7_75t_L g640 ( .A(n_241), .Y(n_640) );
AOI22xp5_ASAP7_75t_SL g433 ( .A1(n_244), .A2(n_282), .B1(n_434), .B2(n_438), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_246), .A2(n_263), .B1(n_553), .B2(n_556), .Y(n_680) );
INVx2_ASAP7_75t_L g318 ( .A(n_249), .Y(n_318) );
INVx1_ASAP7_75t_L g859 ( .A(n_257), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_258), .A2(n_259), .B1(n_464), .B2(n_468), .Y(n_546) );
INVx1_ASAP7_75t_L g1100 ( .A(n_267), .Y(n_1100) );
AOI21xp33_ASAP7_75t_L g548 ( .A1(n_270), .A2(n_451), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_271), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_273), .B(n_606), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_274), .A2(n_299), .B1(n_416), .B2(n_421), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_276), .A2(n_286), .B1(n_490), .B2(n_599), .Y(n_775) );
INVx1_ASAP7_75t_L g481 ( .A(n_277), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_278), .A2(n_738), .B(n_757), .Y(n_737) );
INVx1_ASAP7_75t_L g759 ( .A(n_278), .Y(n_759) );
INVx1_ASAP7_75t_L g669 ( .A(n_281), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_284), .A2(n_303), .B1(n_799), .B2(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g641 ( .A(n_289), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_291), .B(n_337), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_292), .A2(n_306), .B1(n_405), .B2(n_693), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_297), .A2(n_580), .B(n_639), .Y(n_638) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_302), .A2(n_451), .B(n_676), .Y(n_675) );
AOI21xp33_ASAP7_75t_SL g534 ( .A1(n_307), .A2(n_535), .B(n_537), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_324), .B(n_820), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx4_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .C(n_323), .Y(n_315) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_316), .B(n_1072), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_316), .B(n_1073), .Y(n_1076) );
AOI21xp5_ASAP7_75t_L g1104 ( .A1(n_316), .A2(n_323), .B(n_844), .Y(n_1104) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AO21x1_ASAP7_75t_L g1102 ( .A1(n_317), .A2(n_1103), .B(n_1104), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g829 ( .A(n_318), .B(n_830), .Y(n_829) );
AND3x4_ASAP7_75t_L g843 ( .A(n_318), .B(n_831), .C(n_844), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g1072 ( .A(n_319), .B(n_1073), .Y(n_1072) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AO21x2_ASAP7_75t_L g392 ( .A1(n_320), .A2(n_393), .B(n_394), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g1073 ( .A(n_323), .Y(n_1073) );
OAI22xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_589), .B2(n_590), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
XNOR2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_476), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AO22x2_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B1(n_444), .B2(n_475), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND3xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_396), .C(n_433), .Y(n_332) );
INVx1_ASAP7_75t_L g443 ( .A(n_333), .Y(n_443) );
AND3x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_361), .C(n_378), .Y(n_333) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_338), .Y(n_533) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx3_ASAP7_75t_L g449 ( .A(n_339), .Y(n_449) );
BUFx3_ASAP7_75t_L g545 ( .A(n_339), .Y(n_545) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_349), .Y(n_339) );
AND2x2_ASAP7_75t_L g409 ( .A(n_340), .B(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g413 ( .A(n_340), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g437 ( .A(n_340), .B(n_420), .Y(n_437) );
AND2x2_ASAP7_75t_L g461 ( .A(n_340), .B(n_410), .Y(n_461) );
AND2x4_ASAP7_75t_L g470 ( .A(n_340), .B(n_420), .Y(n_470) );
AND2x4_ASAP7_75t_L g553 ( .A(n_340), .B(n_402), .Y(n_553) );
AND2x4_ASAP7_75t_L g556 ( .A(n_340), .B(n_410), .Y(n_556) );
AND2x2_ASAP7_75t_L g580 ( .A(n_340), .B(n_349), .Y(n_580) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_348), .Y(n_340) );
INVx1_ASAP7_75t_L g377 ( .A(n_341), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_345), .Y(n_341) );
NAND2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx2_ASAP7_75t_L g347 ( .A(n_343), .Y(n_347) );
INVx3_ASAP7_75t_L g353 ( .A(n_343), .Y(n_353) );
NAND2xp33_ASAP7_75t_L g359 ( .A(n_343), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g372 ( .A(n_343), .Y(n_372) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_343), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_344), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g387 ( .A1(n_346), .A2(n_372), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g376 ( .A(n_348), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g386 ( .A(n_348), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g401 ( .A(n_348), .Y(n_401) );
AND2x4_ASAP7_75t_L g365 ( .A(n_349), .B(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_L g375 ( .A(n_349), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g425 ( .A(n_349), .B(n_400), .Y(n_425) );
AND2x2_ASAP7_75t_L g451 ( .A(n_349), .B(n_376), .Y(n_451) );
AND2x4_ASAP7_75t_L g468 ( .A(n_349), .B(n_366), .Y(n_468) );
AND2x4_ASAP7_75t_L g474 ( .A(n_349), .B(n_400), .Y(n_474) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_355), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g382 ( .A(n_351), .B(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g403 ( .A(n_351), .B(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g410 ( .A(n_351), .B(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g420 ( .A(n_351), .B(n_355), .Y(n_420) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_353), .B(n_358), .Y(n_357) );
INVxp67_ASAP7_75t_L g368 ( .A(n_353), .Y(n_368) );
NAND3xp33_ASAP7_75t_L g394 ( .A(n_354), .B(n_367), .C(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g404 ( .A(n_356), .Y(n_404) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx4_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx3_ASAP7_75t_L g600 ( .A(n_364), .Y(n_600) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_365), .Y(n_490) );
INVx3_ASAP7_75t_L g804 ( .A(n_365), .Y(n_804) );
AND2x4_ASAP7_75t_L g406 ( .A(n_366), .B(n_402), .Y(n_406) );
AND2x4_ASAP7_75t_L g432 ( .A(n_366), .B(n_410), .Y(n_432) );
AND2x4_ASAP7_75t_L g457 ( .A(n_366), .B(n_410), .Y(n_457) );
AND2x4_ASAP7_75t_L g465 ( .A(n_366), .B(n_402), .Y(n_465) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_371), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g707 ( .A(n_374), .Y(n_707) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_375), .Y(n_489) );
BUFx3_ASAP7_75t_L g577 ( .A(n_375), .Y(n_577) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_375), .Y(n_599) );
BUFx8_ASAP7_75t_SL g637 ( .A(n_375), .Y(n_637) );
AND2x4_ASAP7_75t_L g441 ( .A(n_376), .B(n_420), .Y(n_441) );
AND2x4_ASAP7_75t_L g467 ( .A(n_376), .B(n_420), .Y(n_467) );
AND2x4_ASAP7_75t_L g400 ( .A(n_377), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g485 ( .A(n_380), .Y(n_485) );
INVx4_ASAP7_75t_L g528 ( .A(n_380), .Y(n_528) );
INVx3_ASAP7_75t_L g609 ( .A(n_380), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g702 ( .A1(n_380), .A2(n_703), .B(n_704), .Y(n_702) );
INVx5_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx4f_ASAP7_75t_L g575 ( .A(n_381), .Y(n_575) );
BUFx2_ASAP7_75t_L g779 ( .A(n_381), .Y(n_779) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_386), .Y(n_381) );
AND2x2_ASAP7_75t_L g471 ( .A(n_382), .B(n_386), .Y(n_471) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_382), .B(n_386), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g393 ( .A(n_384), .Y(n_393) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_390), .B(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_390), .B(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_390), .B(n_677), .Y(n_676) );
INVx4_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx3_ASAP7_75t_L g583 ( .A(n_391), .Y(n_583) );
INVx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_392), .Y(n_496) );
AND4x1_ASAP7_75t_L g396 ( .A(n_397), .B(n_407), .C(n_415), .D(n_426), .Y(n_396) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_399), .Y(n_570) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_399), .Y(n_693) );
BUFx6f_ASAP7_75t_L g1061 ( .A(n_399), .Y(n_1061) );
AND2x4_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
AND2x4_ASAP7_75t_L g419 ( .A(n_400), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g429 ( .A(n_400), .B(n_410), .Y(n_429) );
AND2x4_ASAP7_75t_L g456 ( .A(n_400), .B(n_410), .Y(n_456) );
AND2x4_ASAP7_75t_L g464 ( .A(n_400), .B(n_414), .Y(n_464) );
AND2x4_ASAP7_75t_L g473 ( .A(n_400), .B(n_420), .Y(n_473) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g414 ( .A(n_403), .Y(n_414) );
INVx1_ASAP7_75t_L g411 ( .A(n_404), .Y(n_411) );
BUFx3_ASAP7_75t_L g796 ( .A(n_405), .Y(n_796) );
BUFx12f_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx6_ASAP7_75t_L g500 ( .A(n_406), .Y(n_500) );
BUFx8_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_409), .Y(n_522) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_412), .Y(n_793) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_413), .Y(n_459) );
BUFx12f_ASAP7_75t_L g523 ( .A(n_413), .Y(n_523) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_413), .Y(n_564) );
BUFx3_ASAP7_75t_L g612 ( .A(n_413), .Y(n_612) );
BUFx4f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g517 ( .A(n_418), .Y(n_517) );
INVx3_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx12f_ASAP7_75t_L g507 ( .A(n_419), .Y(n_507) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_419), .Y(n_651) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_423), .Y(n_618) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_425), .Y(n_508) );
BUFx5_ASAP7_75t_L g696 ( .A(n_425), .Y(n_696) );
BUFx3_ASAP7_75t_L g744 ( .A(n_425), .Y(n_744) );
BUFx12f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_428), .Y(n_615) );
BUFx12f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_429), .Y(n_504) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_429), .Y(n_653) );
INVx4_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g505 ( .A(n_431), .Y(n_505) );
INVx2_ASAP7_75t_L g525 ( .A(n_431), .Y(n_525) );
INVx4_ASAP7_75t_L g566 ( .A(n_431), .Y(n_566) );
INVx1_ASAP7_75t_L g698 ( .A(n_431), .Y(n_698) );
INVx1_ASAP7_75t_L g717 ( .A(n_431), .Y(n_717) );
INVx2_ASAP7_75t_SL g1058 ( .A(n_431), .Y(n_1058) );
INVx8_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g800 ( .A(n_436), .Y(n_800) );
BUFx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g604 ( .A(n_437), .Y(n_604) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_437), .Y(n_627) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_441), .Y(n_492) );
INVx1_ASAP7_75t_L g536 ( .A(n_441), .Y(n_536) );
BUFx3_ASAP7_75t_L g574 ( .A(n_441), .Y(n_574) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_445), .Y(n_475) );
NAND3x1_ASAP7_75t_L g446 ( .A(n_447), .B(n_454), .C(n_462), .Y(n_446) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_448), .Y(n_664) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g487 ( .A(n_449), .Y(n_487) );
INVx2_ASAP7_75t_L g777 ( .A(n_449), .Y(n_777) );
INVx2_ASAP7_75t_L g808 ( .A(n_449), .Y(n_808) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_458), .Y(n_454) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx4f_ASAP7_75t_L g502 ( .A(n_461), .Y(n_502) );
AND4x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_466), .C(n_469), .D(n_472), .Y(n_462) );
INVx2_ASAP7_75t_L g1089 ( .A(n_467), .Y(n_1089) );
INVx2_ASAP7_75t_L g1095 ( .A(n_468), .Y(n_1095) );
INVx1_ASAP7_75t_L g1093 ( .A(n_470), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_509), .B1(n_587), .B2(n_588), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_478), .Y(n_588) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
XNOR2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
NOR2xp67_ASAP7_75t_L g482 ( .A(n_483), .B(n_497), .Y(n_482) );
NAND4xp25_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .C(n_488), .D(n_491), .Y(n_483) );
BUFx3_ASAP7_75t_L g802 ( .A(n_489), .Y(n_802) );
BUFx3_ASAP7_75t_L g756 ( .A(n_490), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx2_ASAP7_75t_L g705 ( .A(n_495), .Y(n_705) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_496), .Y(n_539) );
INVx2_ASAP7_75t_L g751 ( .A(n_496), .Y(n_751) );
NAND4xp25_ASAP7_75t_SL g497 ( .A(n_498), .B(n_501), .C(n_503), .D(n_506), .Y(n_497) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx3_ASAP7_75t_L g519 ( .A(n_500), .Y(n_519) );
INVx1_ASAP7_75t_L g613 ( .A(n_500), .Y(n_613) );
INVx5_ASAP7_75t_L g767 ( .A(n_500), .Y(n_767) );
INVx2_ASAP7_75t_L g1056 ( .A(n_500), .Y(n_1056) );
BUFx2_ASAP7_75t_SL g788 ( .A(n_504), .Y(n_788) );
BUFx2_ASAP7_75t_SL g789 ( .A(n_505), .Y(n_789) );
INVx1_ASAP7_75t_L g587 ( .A(n_509), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B1(n_558), .B2(n_585), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
XOR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_541), .Y(n_511) );
INVx1_ASAP7_75t_L g540 ( .A(n_514), .Y(n_540) );
NAND4xp75_ASAP7_75t_L g514 ( .A(n_515), .B(n_520), .C(n_526), .D(n_530), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_518), .Y(n_515) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_524), .Y(n_520) );
BUFx3_ASAP7_75t_L g792 ( .A(n_522), .Y(n_792) );
BUFx3_ASAP7_75t_L g742 ( .A(n_523), .Y(n_742) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .Y(n_526) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_534), .Y(n_530) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_539), .B(n_723), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_539), .B(n_774), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g1067 ( .A(n_539), .B(n_1068), .Y(n_1067) );
NOR2xp33_ASAP7_75t_L g1099 ( .A(n_539), .B(n_1100), .Y(n_1099) );
OR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_551), .Y(n_542) );
NAND4xp25_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .C(n_547), .D(n_548), .Y(n_543) );
INVx1_ASAP7_75t_L g607 ( .A(n_545), .Y(n_607) );
BUFx3_ASAP7_75t_L g701 ( .A(n_545), .Y(n_701) );
NAND4xp25_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .C(n_555), .D(n_557), .Y(n_551) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx3_ASAP7_75t_L g586 ( .A(n_560), .Y(n_586) );
XNOR2x1_ASAP7_75t_L g560 ( .A(n_561), .B(n_584), .Y(n_560) );
NAND4xp75_ASAP7_75t_L g561 ( .A(n_562), .B(n_567), .C(n_571), .D(n_576), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
BUFx3_ASAP7_75t_L g616 ( .A(n_570), .Y(n_616) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
BUFx2_ASAP7_75t_L g799 ( .A(n_574), .Y(n_799) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g1098 ( .A(n_580), .Y(n_1098) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_583), .B(n_640), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_583), .B(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_583), .B(n_810), .Y(n_809) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_730), .B1(n_816), .B2(n_817), .Y(n_590) );
INVx1_ASAP7_75t_L g816 ( .A(n_591), .Y(n_816) );
XNOR2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_686), .Y(n_591) );
XNOR2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_643), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_621), .B1(n_622), .B2(n_642), .Y(n_593) );
INVx1_ASAP7_75t_L g642 ( .A(n_594), .Y(n_642) );
XOR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_620), .Y(n_594) );
NOR2x1_ASAP7_75t_L g595 ( .A(n_596), .B(n_610), .Y(n_595) );
NAND4xp25_ASAP7_75t_L g596 ( .A(n_597), .B(n_601), .C(n_605), .D(n_608), .Y(n_596) );
BUFx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g720 ( .A(n_599), .Y(n_720) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g666 ( .A(n_603), .Y(n_666) );
INVx1_ASAP7_75t_L g753 ( .A(n_603), .Y(n_753) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g709 ( .A(n_604), .Y(n_709) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND4xp25_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .C(n_617), .D(n_619), .Y(n_610) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
XOR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_641), .Y(n_622) );
NOR4xp75_ASAP7_75t_L g623 ( .A(n_624), .B(n_628), .C(n_631), .D(n_634), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_632), .B(n_633), .Y(n_631) );
OAI21x1_ASAP7_75t_SL g634 ( .A1(n_635), .A2(n_636), .B(n_638), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_667), .B(n_683), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_SL g685 ( .A(n_646), .Y(n_685) );
XNOR2x1_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NOR2x1_ASAP7_75t_L g648 ( .A(n_649), .B(n_656), .Y(n_648) );
NAND4xp25_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .C(n_654), .D(n_655), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_663), .C(n_665), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_662), .Y(n_658) );
BUFx3_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_668), .B(n_684), .Y(n_683) );
XNOR2x1_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_678), .Y(n_670) );
NAND4xp25_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .C(n_674), .D(n_675), .Y(n_671) );
NAND4xp25_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .C(n_681), .D(n_682), .Y(n_678) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
XNOR2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_711), .Y(n_688) );
XNOR2x1_ASAP7_75t_L g689 ( .A(n_690), .B(n_710), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_699), .Y(n_690) );
NAND4xp25_ASAP7_75t_SL g691 ( .A(n_692), .B(n_694), .C(n_695), .D(n_697), .Y(n_691) );
BUFx3_ASAP7_75t_L g795 ( .A(n_693), .Y(n_795) );
BUFx3_ASAP7_75t_L g786 ( .A(n_696), .Y(n_786) );
NAND3xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_706), .C(n_708), .Y(n_699) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NAND4xp75_ASAP7_75t_L g713 ( .A(n_714), .B(n_718), .C(n_724), .D(n_727), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
OA21x2_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B(n_721), .Y(n_718) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
AND2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_781), .B(n_811), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI22x1_ASAP7_75t_L g818 ( .A1(n_732), .A2(n_812), .B1(n_814), .B2(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g815 ( .A(n_735), .Y(n_815) );
OA22x2_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B1(n_761), .B2(n_780), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_746), .Y(n_738) );
INVxp67_ASAP7_75t_L g760 ( .A(n_739), .Y(n_760) );
NAND4xp25_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .C(n_743), .D(n_745), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_746), .B(n_759), .Y(n_758) );
NAND4xp25_ASAP7_75t_L g746 ( .A(n_747), .B(n_752), .C(n_754), .D(n_755), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx3_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_760), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_759), .A2(n_861), .B1(n_863), .B2(n_865), .Y(n_860) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_SL g780 ( .A(n_763), .Y(n_780) );
NOR2x1_ASAP7_75t_L g764 ( .A(n_765), .B(n_771), .Y(n_764) );
NAND4xp25_ASAP7_75t_L g765 ( .A(n_766), .B(n_768), .C(n_769), .D(n_770), .Y(n_765) );
NAND4xp25_ASAP7_75t_SL g771 ( .A(n_772), .B(n_775), .C(n_776), .D(n_778), .Y(n_771) );
INVx1_ASAP7_75t_L g819 ( .A(n_781), .Y(n_819) );
BUFx3_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_SL g813 ( .A(n_782), .Y(n_813) );
NAND4xp75_ASAP7_75t_L g783 ( .A(n_784), .B(n_790), .C(n_797), .D(n_805), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_787), .Y(n_784) );
AND2x2_ASAP7_75t_L g790 ( .A(n_791), .B(n_794), .Y(n_790) );
AND2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_801), .Y(n_797) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_814), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_1043), .B1(n_1046), .B2(n_1069), .C(n_1074), .Y(n_820) );
O2A1O1Ixp33_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_915), .B(n_956), .C(n_999), .Y(n_821) );
NAND3xp33_ASAP7_75t_L g822 ( .A(n_823), .B(n_885), .C(n_892), .Y(n_822) );
AOI222xp33_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_852), .B1(n_866), .B2(n_873), .C1(n_877), .C2(n_882), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_824), .B(n_874), .Y(n_1012) );
AND2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_839), .Y(n_824) );
INVx1_ASAP7_75t_L g867 ( .A(n_825), .Y(n_867) );
NAND2xp5_ASAP7_75t_SL g889 ( .A(n_825), .B(n_890), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_825), .B(n_902), .Y(n_901) );
INVx2_ASAP7_75t_L g906 ( .A(n_825), .Y(n_906) );
INVx2_ASAP7_75t_L g918 ( .A(n_825), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_825), .B(n_880), .Y(n_928) );
BUFx6f_ASAP7_75t_L g936 ( .A(n_825), .Y(n_936) );
AND2x2_ASAP7_75t_L g961 ( .A(n_825), .B(n_949), .Y(n_961) );
AND2x2_ASAP7_75t_L g991 ( .A(n_825), .B(n_853), .Y(n_991) );
NOR2x1_ASAP7_75t_L g1002 ( .A(n_825), .B(n_891), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_825), .B(n_854), .Y(n_1010) );
NAND2xp5_ASAP7_75t_SL g1030 ( .A(n_825), .B(n_1031), .Y(n_1030) );
INVx4_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_826), .B(n_869), .Y(n_878) );
OR2x2_ASAP7_75t_L g894 ( .A(n_826), .B(n_895), .Y(n_894) );
AND2x2_ASAP7_75t_L g900 ( .A(n_826), .B(n_854), .Y(n_900) );
AND2x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_835), .Y(n_826) );
INVx3_ASAP7_75t_L g856 ( .A(n_828), .Y(n_856) );
AND2x4_ASAP7_75t_L g828 ( .A(n_829), .B(n_831), .Y(n_828) );
AND2x2_ASAP7_75t_L g836 ( .A(n_829), .B(n_837), .Y(n_836) );
AND2x2_ASAP7_75t_L g847 ( .A(n_829), .B(n_837), .Y(n_847) );
AND2x4_ASAP7_75t_L g862 ( .A(n_829), .B(n_837), .Y(n_862) );
AND2x4_ASAP7_75t_L g833 ( .A(n_831), .B(n_834), .Y(n_833) );
AND2x4_ASAP7_75t_L g845 ( .A(n_831), .B(n_834), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_831), .B(n_834), .Y(n_858) );
AND2x2_ASAP7_75t_L g838 ( .A(n_834), .B(n_837), .Y(n_838) );
AND2x2_ASAP7_75t_L g848 ( .A(n_834), .B(n_837), .Y(n_848) );
AND2x4_ASAP7_75t_L g864 ( .A(n_834), .B(n_837), .Y(n_864) );
AND2x2_ASAP7_75t_L g907 ( .A(n_839), .B(n_895), .Y(n_907) );
AND2x2_ASAP7_75t_L g996 ( .A(n_839), .B(n_881), .Y(n_996) );
INVx1_ASAP7_75t_L g1035 ( .A(n_839), .Y(n_1035) );
AND2x2_ASAP7_75t_L g839 ( .A(n_840), .B(n_849), .Y(n_839) );
AND2x2_ASAP7_75t_L g873 ( .A(n_840), .B(n_874), .Y(n_873) );
AND2x2_ASAP7_75t_L g880 ( .A(n_840), .B(n_881), .Y(n_880) );
OR2x2_ASAP7_75t_L g891 ( .A(n_840), .B(n_849), .Y(n_891) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
OR2x2_ASAP7_75t_L g921 ( .A(n_841), .B(n_849), .Y(n_921) );
AND2x2_ASAP7_75t_L g927 ( .A(n_841), .B(n_849), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_841), .B(n_881), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_841), .B(n_874), .Y(n_985) );
AND2x2_ASAP7_75t_L g841 ( .A(n_842), .B(n_846), .Y(n_841) );
INVx1_ASAP7_75t_L g903 ( .A(n_849), .Y(n_903) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_849), .B(n_895), .Y(n_1040) );
AND2x2_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_852), .B(n_887), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_852), .B(n_909), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g1033 ( .A(n_852), .B(n_1034), .Y(n_1033) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g869 ( .A(n_854), .Y(n_869) );
AND2x2_ASAP7_75t_L g923 ( .A(n_854), .B(n_870), .Y(n_923) );
OR2x2_ASAP7_75t_L g933 ( .A(n_854), .B(n_870), .Y(n_933) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_854), .B(n_1018), .Y(n_1017) );
OR2x2_ASAP7_75t_L g854 ( .A(n_855), .B(n_860), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_855) );
OAI221xp5_ASAP7_75t_L g952 ( .A1(n_856), .A2(n_858), .B1(n_953), .B2(n_954), .C(n_955), .Y(n_952) );
INVx1_ASAP7_75t_L g1045 ( .A(n_856), .Y(n_1045) );
INVx3_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx2_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVxp67_ASAP7_75t_L g1008 ( .A(n_866), .Y(n_1008) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_867), .B(n_884), .Y(n_945) );
OAI322xp33_ASAP7_75t_L g893 ( .A1(n_868), .A2(n_890), .A3(n_894), .B1(n_897), .B2(n_898), .C1(n_899), .C2(n_901), .Y(n_893) );
OAI211xp5_ASAP7_75t_SL g915 ( .A1(n_868), .A2(n_916), .B(n_922), .C(n_939), .Y(n_915) );
INVx1_ASAP7_75t_L g982 ( .A(n_868), .Y(n_982) );
OR2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .Y(n_868) );
AND2x2_ASAP7_75t_L g942 ( .A(n_869), .B(n_931), .Y(n_942) );
AND2x2_ASAP7_75t_L g947 ( .A(n_869), .B(n_870), .Y(n_947) );
NOR2xp33_ASAP7_75t_L g1003 ( .A(n_869), .B(n_1004), .Y(n_1003) );
INVx2_ASAP7_75t_L g1021 ( .A(n_869), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_870), .Y(n_884) );
INVx2_ASAP7_75t_L g897 ( .A(n_870), .Y(n_897) );
OR2x2_ASAP7_75t_L g964 ( .A(n_870), .B(n_911), .Y(n_964) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_870), .B(n_912), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_870), .B(n_911), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_870), .B(n_910), .Y(n_1042) );
AND2x2_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g898 ( .A(n_873), .Y(n_898) );
NOR2xp33_ASAP7_75t_L g972 ( .A(n_873), .B(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g881 ( .A(n_874), .Y(n_881) );
INVx1_ASAP7_75t_SL g896 ( .A(n_874), .Y(n_896) );
OR2x2_ASAP7_75t_L g920 ( .A(n_874), .B(n_921), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_874), .B(n_890), .Y(n_941) );
AND2x2_ASAP7_75t_L g949 ( .A(n_874), .B(n_903), .Y(n_949) );
OR2x2_ASAP7_75t_L g974 ( .A(n_874), .B(n_891), .Y(n_974) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_874), .B(n_1002), .Y(n_1001) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g877 ( .A(n_878), .B(n_879), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g984 ( .A(n_878), .B(n_985), .Y(n_984) );
OAI221xp5_ASAP7_75t_L g977 ( .A1(n_879), .A2(n_889), .B1(n_978), .B2(n_980), .C(n_983), .Y(n_977) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
NOR2x1_ASAP7_75t_R g888 ( .A(n_881), .B(n_889), .Y(n_888) );
AND2x2_ASAP7_75t_L g902 ( .A(n_881), .B(n_903), .Y(n_902) );
AND2x2_ASAP7_75t_L g926 ( .A(n_881), .B(n_927), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_881), .B(n_1014), .Y(n_1013) );
OAI322xp33_ASAP7_75t_L g971 ( .A1(n_882), .A2(n_905), .A3(n_936), .B1(n_964), .B2(n_972), .C1(n_975), .C2(n_976), .Y(n_971) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_884), .B(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVxp67_ASAP7_75t_SL g887 ( .A(n_888), .Y(n_887) );
OAI21xp5_ASAP7_75t_SL g995 ( .A1(n_890), .A2(n_996), .B(n_997), .Y(n_995) );
INVx3_ASAP7_75t_SL g890 ( .A(n_891), .Y(n_890) );
OAI21xp5_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_904), .B(n_908), .Y(n_892) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_894), .B(n_1035), .Y(n_1034) );
AND2x2_ASAP7_75t_L g967 ( .A(n_895), .B(n_927), .Y(n_967) );
AND2x4_ASAP7_75t_L g987 ( .A(n_895), .B(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_897), .A2(n_898), .B1(n_959), .B2(n_960), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_897), .A2(n_962), .B1(n_1020), .B2(n_1022), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_897), .B(n_900), .Y(n_1038) );
O2A1O1Ixp33_ASAP7_75t_L g934 ( .A1(n_898), .A2(n_935), .B(n_937), .C(n_938), .Y(n_934) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
NOR2xp67_ASAP7_75t_SL g1020 ( .A(n_905), .B(n_1021), .Y(n_1020) );
NOR2xp33_ASAP7_75t_L g1022 ( .A(n_905), .B(n_1023), .Y(n_1022) );
NAND2xp67_ASAP7_75t_L g905 ( .A(n_906), .B(n_907), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_906), .B(n_927), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_906), .B(n_923), .Y(n_998) );
AOI221xp5_ASAP7_75t_L g922 ( .A1(n_907), .A2(n_923), .B1(n_924), .B2(n_929), .C(n_934), .Y(n_922) );
INVx1_ASAP7_75t_L g975 ( .A(n_907), .Y(n_975) );
NOR2xp33_ASAP7_75t_L g981 ( .A(n_908), .B(n_982), .Y(n_981) );
INVx1_ASAP7_75t_SL g908 ( .A(n_909), .Y(n_908) );
AOI221xp5_ASAP7_75t_L g1024 ( .A1(n_909), .A2(n_1018), .B1(n_1025), .B2(n_1026), .C(n_1036), .Y(n_1024) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g931 ( .A(n_912), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .Y(n_917) );
INVx1_ASAP7_75t_L g966 ( .A(n_918), .Y(n_966) );
NOR2xp33_ASAP7_75t_L g970 ( .A(n_918), .B(n_920), .Y(n_970) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g988 ( .A(n_921), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_921), .B(n_1015), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_925), .B(n_928), .Y(n_924) );
OAI221xp5_ASAP7_75t_L g1036 ( .A1(n_925), .A2(n_964), .B1(n_1037), .B2(n_1039), .C(n_1041), .Y(n_1036) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_926), .B(n_982), .Y(n_994) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_926), .B(n_935), .Y(n_1025) );
INVx1_ASAP7_75t_L g1015 ( .A(n_927), .Y(n_1015) );
INVx1_ASAP7_75t_L g976 ( .A(n_929), .Y(n_976) );
AND2x2_ASAP7_75t_L g929 ( .A(n_930), .B(n_932), .Y(n_929) );
AOI221xp5_ASAP7_75t_L g939 ( .A1(n_930), .A2(n_940), .B1(n_942), .B2(n_943), .C(n_950), .Y(n_939) );
INVx2_ASAP7_75t_L g962 ( .A(n_930), .Y(n_962) );
BUFx3_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_931), .B(n_933), .Y(n_979) );
INVx2_ASAP7_75t_L g992 ( .A(n_931), .Y(n_992) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx2_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_936), .B(n_947), .Y(n_959) );
INVx1_ASAP7_75t_L g969 ( .A(n_938), .Y(n_969) );
OAI21xp33_ASAP7_75t_L g1041 ( .A1(n_940), .A2(n_984), .B(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_944), .A2(n_945), .B1(n_946), .B2(n_948), .Y(n_943) );
A2O1A1Ixp33_ASAP7_75t_L g1026 ( .A1(n_946), .A2(n_1027), .B(n_1028), .C(n_1032), .Y(n_1026) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx2_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
AOI211xp5_ASAP7_75t_L g986 ( .A1(n_951), .A2(n_987), .B(n_989), .C(n_993), .Y(n_986) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
NAND4xp25_ASAP7_75t_L g956 ( .A(n_957), .B(n_968), .C(n_986), .D(n_995), .Y(n_956) );
AOI21xp5_ASAP7_75t_L g957 ( .A1(n_958), .A2(n_962), .B(n_963), .Y(n_957) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
NOR2xp33_ASAP7_75t_L g1028 ( .A(n_961), .B(n_1029), .Y(n_1028) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_964), .B(n_965), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_966), .B(n_967), .Y(n_965) );
NOR2xp33_ASAP7_75t_L g1006 ( .A(n_967), .B(n_996), .Y(n_1006) );
AOI211xp5_ASAP7_75t_L g968 ( .A1(n_969), .A2(n_970), .B(n_971), .C(n_977), .Y(n_968) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVxp67_ASAP7_75t_SL g980 ( .A(n_981), .Y(n_980) );
INVx1_ASAP7_75t_L g1031 ( .A(n_985), .Y(n_1031) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_991), .B(n_992), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_992), .B(n_1010), .Y(n_1009) );
INVxp67_ASAP7_75t_SL g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g1027 ( .A(n_996), .Y(n_1027) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
NAND3xp33_ASAP7_75t_SL g999 ( .A(n_1000), .B(n_1019), .C(n_1024), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1003), .B1(n_1005), .B2(n_1007), .C(n_1011), .Y(n_1000) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
NAND2xp5_ASAP7_75t_SL g1007 ( .A(n_1008), .B(n_1009), .Y(n_1007) );
AOI21xp33_ASAP7_75t_L g1011 ( .A1(n_1012), .A2(n_1013), .B(n_1016), .Y(n_1011) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
INVx2_ASAP7_75t_L g1023 ( .A(n_1021), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_1021), .B(n_1040), .Y(n_1039) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
CKINVDCx5p33_ASAP7_75t_R g1043 ( .A(n_1044), .Y(n_1043) );
HB1xp67_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
INVx2_ASAP7_75t_SL g1046 ( .A(n_1047), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
BUFx2_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
XNOR2x1_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1053), .Y(n_1050) );
CKINVDCx5p33_ASAP7_75t_R g1051 ( .A(n_1052), .Y(n_1051) );
NOR2x1_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1062), .Y(n_1053) );
NAND4xp25_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1057), .C(n_1059), .D(n_1060), .Y(n_1054) );
NAND4xp25_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .C(n_1065), .D(n_1066), .Y(n_1062) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
HB1xp67_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
HB1xp67_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
NAND4xp75_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1083), .C(n_1086), .D(n_1097), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1082), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1085), .Y(n_1083) );
NOR2xp33_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1092), .Y(n_1086) );
OAI21xp33_ASAP7_75t_L g1087 ( .A1(n_1088), .A2(n_1089), .B(n_1090), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_1093), .A2(n_1094), .B1(n_1095), .B2(n_1096), .Y(n_1092) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
endmodule