module fake_ariane_2388_n_411 (n_66, n_8, n_56, n_60, n_24, n_7, n_22, n_71, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_64, n_17, n_4, n_41, n_50, n_38, n_55, n_2, n_62, n_47, n_18, n_32, n_28, n_37, n_58, n_65, n_9, n_51, n_67, n_45, n_11, n_34, n_69, n_26, n_3, n_46, n_14, n_0, n_52, n_36, n_68, n_72, n_73, n_33, n_44, n_19, n_30, n_39, n_40, n_59, n_31, n_42, n_57, n_16, n_63, n_5, n_12, n_15, n_53, n_21, n_70, n_23, n_61, n_35, n_10, n_54, n_25, n_411);

input n_66;
input n_8;
input n_56;
input n_60;
input n_24;
input n_7;
input n_22;
input n_71;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_64;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_55;
input n_2;
input n_62;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_58;
input n_65;
input n_9;
input n_51;
input n_67;
input n_45;
input n_11;
input n_34;
input n_69;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_52;
input n_36;
input n_68;
input n_72;
input n_73;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_59;
input n_31;
input n_42;
input n_57;
input n_16;
input n_63;
input n_5;
input n_12;
input n_15;
input n_53;
input n_21;
input n_70;
input n_23;
input n_61;
input n_35;
input n_10;
input n_54;
input n_25;

output n_411;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_124;
wire n_119;
wire n_386;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_183;
wire n_373;
wire n_299;
wire n_133;
wire n_205;
wire n_341;
wire n_109;
wire n_245;
wire n_96;
wire n_319;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_103;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_387;
wire n_406;
wire n_117;
wire n_139;
wire n_85;
wire n_130;
wire n_391;
wire n_349;
wire n_346;
wire n_214;
wire n_348;
wire n_410;
wire n_379;
wire n_162;
wire n_138;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_385;
wire n_327;
wire n_77;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_87;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_167;
wire n_90;
wire n_153;
wire n_269;
wire n_75;
wire n_158;
wire n_259;
wire n_95;
wire n_143;
wire n_152;
wire n_405;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_320;
wire n_309;
wire n_115;
wire n_331;
wire n_401;
wire n_267;
wire n_335;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_398;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_79;
wire n_271;
wire n_247;
wire n_91;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_82;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_400;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_248;
wire n_301;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_93;
wire n_108;
wire n_303;
wire n_168;
wire n_81;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_88;
wire n_141;
wire n_390;
wire n_104;
wire n_314;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_392;
wire n_376;
wire n_221;
wire n_321;
wire n_86;
wire n_361;
wire n_89;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_74;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_84;
wire n_371;
wire n_199;
wire n_107;
wire n_217;
wire n_178;
wire n_308;
wire n_201;
wire n_343;
wire n_287;
wire n_302;
wire n_380;
wire n_94;
wire n_284;
wire n_249;
wire n_123;
wire n_212;
wire n_355;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_135;
wire n_409;
wire n_171;
wire n_384;
wire n_102;
wire n_182;
wire n_316;
wire n_196;
wire n_125;
wire n_407;
wire n_254;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_78;
wire n_99;
wire n_216;
wire n_223;
wire n_403;
wire n_83;
wire n_389;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_110;
wire n_304;
wire n_306;
wire n_313;
wire n_92;
wire n_203;
wire n_378;
wire n_150;
wire n_98;
wire n_375;
wire n_113;
wire n_114;
wire n_324;
wire n_337;
wire n_111;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_100;
wire n_132;
wire n_147;
wire n_204;
wire n_76;
wire n_342;
wire n_246;
wire n_159;
wire n_358;
wire n_105;
wire n_131;
wire n_263;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_101;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_112;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_121;
wire n_118;
wire n_353;
wire n_241;
wire n_357;
wire n_191;
wire n_382;
wire n_80;
wire n_211;
wire n_97;
wire n_408;
wire n_322;
wire n_251;
wire n_116;
wire n_397;
wire n_351;
wire n_393;
wire n_359;
wire n_155;
wire n_127;

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_10),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_8),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_32),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_1),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVxp33_ASAP7_75t_SL g83 ( 
.A(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_10),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVxp33_ASAP7_75t_SL g91 ( 
.A(n_58),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_66),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_1),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_5),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_13),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_9),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_68),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_11),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_12),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

INVxp33_ASAP7_75t_SL g110 ( 
.A(n_23),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_7),
.Y(n_111)
);

INVxp33_ASAP7_75t_SL g112 ( 
.A(n_48),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_29),
.Y(n_113)
);

INVxp67_ASAP7_75t_SL g114 ( 
.A(n_71),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_67),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_24),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_17),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_14),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_18),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_40),
.Y(n_120)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_46),
.Y(n_121)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_44),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_12),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_28),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_52),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_43),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_8),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_2),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_26),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_35),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_4),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_21),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_127),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_79),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_79),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_75),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_101),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_0),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_76),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_102),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_117),
.B(n_0),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

BUFx10_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_R g156 ( 
.A(n_116),
.B(n_113),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

NAND2xp33_ASAP7_75t_R g160 ( 
.A(n_115),
.B(n_31),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_77),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_124),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_115),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_131),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_R g170 ( 
.A(n_129),
.B(n_33),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_131),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_R g174 ( 
.A(n_129),
.B(n_27),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_133),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_100),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_88),
.B(n_3),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_89),
.A2(n_5),
.B(n_6),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_89),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_7),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_81),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_90),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_78),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_97),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_133),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_83),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_83),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_82),
.Y(n_192)
);

AO21x2_ASAP7_75t_L g193 ( 
.A1(n_84),
.A2(n_106),
.B(n_136),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_96),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_91),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_104),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

AOI211xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_153),
.B(n_147),
.C(n_191),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_194),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_120),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_134),
.Y(n_205)
);

AO22x1_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_91),
.B1(n_110),
.B2(n_112),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_188),
.B(n_139),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_139),
.B(n_103),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_140),
.B(n_146),
.Y(n_210)
);

AO22x2_ASAP7_75t_L g211 ( 
.A1(n_141),
.A2(n_103),
.B1(n_130),
.B2(n_126),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_108),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

AO22x2_ASAP7_75t_L g218 ( 
.A1(n_142),
.A2(n_130),
.B1(n_126),
.B2(n_137),
.Y(n_218)
);

AO22x2_ASAP7_75t_L g219 ( 
.A1(n_143),
.A2(n_128),
.B1(n_123),
.B2(n_109),
.Y(n_219)
);

AO22x1_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_110),
.B1(n_112),
.B2(n_94),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_157),
.B(n_122),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_184),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

OAI221xp5_ASAP7_75t_L g227 ( 
.A1(n_177),
.A2(n_121),
.B1(n_114),
.B2(n_80),
.C(n_119),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_181),
.A2(n_118),
.B(n_16),
.C(n_17),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_183),
.B(n_15),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_45),
.Y(n_234)
);

CKINVDCx11_ASAP7_75t_R g235 ( 
.A(n_144),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_138),
.A2(n_16),
.B1(n_18),
.B2(n_34),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_140),
.B(n_36),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_178),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_151),
.B(n_38),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_179),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_146),
.B(n_49),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_148),
.B(n_70),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_156),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_138),
.A2(n_62),
.B1(n_63),
.B2(n_195),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_145),
.B(n_168),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_203),
.B(n_148),
.Y(n_249)
);

AO32x1_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_179),
.A3(n_155),
.B1(n_170),
.B2(n_160),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_195),
.Y(n_252)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_150),
.C(n_168),
.Y(n_253)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_202),
.A2(n_179),
.B(n_155),
.C(n_174),
.Y(n_254)
);

BUFx4f_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_150),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_234),
.B(n_215),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_227),
.A2(n_190),
.B1(n_173),
.B2(n_169),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_190),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_152),
.B(n_144),
.C(n_163),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_163),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_202),
.A2(n_166),
.B(n_205),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_197),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_205),
.A2(n_198),
.B(n_199),
.C(n_200),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_201),
.B(n_224),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g270 ( 
.A1(n_238),
.A2(n_247),
.B1(n_246),
.B2(n_223),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_212),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_245),
.A2(n_244),
.B(n_240),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_236),
.A2(n_237),
.B(n_233),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_230),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_204),
.A2(n_207),
.B(n_230),
.C(n_245),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_222),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_219),
.B(n_208),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_206),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_220),
.B(n_218),
.Y(n_281)
);

O2A1O1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_219),
.A2(n_218),
.B(n_211),
.C(n_235),
.Y(n_282)
);

O2A1O1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_211),
.A2(n_147),
.B(n_202),
.C(n_228),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_203),
.B(n_139),
.Y(n_284)
);

O2A1O1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_202),
.A2(n_147),
.B(n_228),
.C(n_177),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_227),
.A2(n_75),
.B1(n_98),
.B2(n_77),
.Y(n_286)
);

AND2x4_ASAP7_75t_L g287 ( 
.A(n_221),
.B(n_224),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_227),
.A2(n_75),
.B1(n_98),
.B2(n_77),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_225),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_225),
.A2(n_234),
.B(n_215),
.Y(n_290)
);

O2A1O1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_260),
.A2(n_268),
.B(n_285),
.C(n_256),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_289),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_252),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_254),
.A2(n_274),
.B(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_289),
.B(n_283),
.Y(n_298)
);

AO21x2_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_276),
.B(n_281),
.Y(n_299)
);

AO21x2_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_266),
.B(n_269),
.Y(n_300)
);

OAI21xp33_ASAP7_75t_L g301 ( 
.A1(n_251),
.A2(n_258),
.B(n_267),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_255),
.A2(n_259),
.B1(n_288),
.B2(n_286),
.Y(n_303)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_249),
.A2(n_284),
.B(n_280),
.Y(n_304)
);

AO21x2_ASAP7_75t_L g305 ( 
.A1(n_250),
.A2(n_270),
.B(n_264),
.Y(n_305)
);

O2A1O1Ixp33_ASAP7_75t_SL g306 ( 
.A1(n_265),
.A2(n_262),
.B(n_271),
.C(n_287),
.Y(n_306)
);

OAI21x1_ASAP7_75t_SL g307 ( 
.A1(n_275),
.A2(n_285),
.B(n_245),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g309 ( 
.A1(n_275),
.A2(n_289),
.B(n_239),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_260),
.B(n_210),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_286),
.A2(n_288),
.B1(n_255),
.B2(n_242),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_257),
.A2(n_290),
.B(n_254),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_257),
.A2(n_290),
.B(n_254),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_261),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_257),
.A2(n_290),
.B(n_254),
.Y(n_315)
);

BUFx8_ASAP7_75t_L g316 ( 
.A(n_261),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

AOI21x1_ASAP7_75t_L g319 ( 
.A1(n_257),
.A2(n_234),
.B(n_290),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_260),
.B(n_210),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_260),
.B(n_285),
.C(n_268),
.Y(n_321)
);

OR2x6_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_281),
.Y(n_322)
);

NAND2x1p5_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_239),
.Y(n_323)
);

CKINVDCx11_ASAP7_75t_R g324 ( 
.A(n_261),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_261),
.Y(n_325)
);

AOI21xp33_ASAP7_75t_L g326 ( 
.A1(n_260),
.A2(n_259),
.B(n_285),
.Y(n_326)
);

CKINVDCx11_ASAP7_75t_R g327 ( 
.A(n_324),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_310),
.A2(n_320),
.B1(n_292),
.B2(n_293),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_300),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_316),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_295),
.Y(n_332)
);

OR2x6_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_304),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_295),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_311),
.A2(n_303),
.B1(n_302),
.B2(n_305),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_291),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_325),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_R g340 ( 
.A(n_314),
.B(n_308),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_303),
.B(n_309),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_322),
.Y(n_343)
);

NOR3xp33_ASAP7_75t_SL g344 ( 
.A(n_301),
.B(n_321),
.C(n_294),
.Y(n_344)
);

NOR3xp33_ASAP7_75t_SL g345 ( 
.A(n_313),
.B(n_315),
.C(n_312),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_322),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_328),
.A2(n_313),
.B1(n_318),
.B2(n_317),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_345),
.A2(n_318),
.B1(n_323),
.B2(n_319),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_298),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_305),
.Y(n_350)
);

AOI221xp5_ASAP7_75t_L g351 ( 
.A1(n_344),
.A2(n_306),
.B1(n_307),
.B2(n_305),
.C(n_300),
.Y(n_351)
);

CKINVDCx10_ASAP7_75t_R g352 ( 
.A(n_338),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_332),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_339),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_334),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_342),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_337),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_299),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_299),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_340),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_358),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_353),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_353),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_358),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_352),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_357),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_355),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_350),
.B(n_335),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_331),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_343),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_355),
.B(n_356),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_360),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_330),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_371),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_365),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_356),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_371),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_362),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_346),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_363),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_370),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_329),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_346),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_378),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_361),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_368),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_382),
.Y(n_388)
);

OAI222xp33_ASAP7_75t_L g389 ( 
.A1(n_382),
.A2(n_368),
.B1(n_343),
.B2(n_361),
.C1(n_364),
.C2(n_333),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_375),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_364),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_385),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_381),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_385),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_376),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_391),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_380),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_392),
.Y(n_398)
);

AOI221x1_ASAP7_75t_L g399 ( 
.A1(n_396),
.A2(n_384),
.B1(n_383),
.B2(n_348),
.C(n_347),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_395),
.A2(n_390),
.B1(n_384),
.B2(n_379),
.Y(n_400)
);

AND3x1_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_390),
.C(n_327),
.Y(n_401)
);

OAI211xp5_ASAP7_75t_L g402 ( 
.A1(n_394),
.A2(n_392),
.B(n_391),
.C(n_372),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_393),
.A2(n_348),
.B(n_349),
.Y(n_403)
);

NOR2x1_ASAP7_75t_L g404 ( 
.A(n_402),
.B(n_386),
.Y(n_404)
);

NAND3xp33_ASAP7_75t_SL g405 ( 
.A(n_400),
.B(n_397),
.C(n_386),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_405),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_406),
.A2(n_404),
.B(n_401),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_407),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_408),
.Y(n_409)
);

AOI222xp33_ASAP7_75t_L g410 ( 
.A1(n_409),
.A2(n_399),
.B1(n_327),
.B2(n_389),
.C1(n_351),
.C2(n_397),
.Y(n_410)
);

AOI221xp5_ASAP7_75t_L g411 ( 
.A1(n_410),
.A2(n_399),
.B1(n_403),
.B2(n_398),
.C(n_351),
.Y(n_411)
);


endmodule