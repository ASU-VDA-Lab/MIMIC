module fake_jpeg_4564_n_208 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_0),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_0),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_39),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_33),
.Y(n_38)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_17),
.B1(n_22),
.B2(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_17),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_58),
.B1(n_67),
.B2(n_68),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_34),
.A2(n_22),
.B1(n_32),
.B2(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_17),
.Y(n_63)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_28),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_18),
.B1(n_32),
.B2(n_29),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_44),
.B1(n_39),
.B2(n_24),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_52),
.C(n_59),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_19),
.C(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_27),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_40),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_91),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_44),
.B1(n_39),
.B2(n_24),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_23),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_23),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_62),
.A2(n_26),
.B1(n_33),
.B2(n_25),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_53),
.B1(n_51),
.B2(n_37),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_19),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_20),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_93),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_55),
.B1(n_60),
.B2(n_51),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_97),
.B1(n_108),
.B2(n_88),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_71),
.B1(n_79),
.B2(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_113),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_51),
.B1(n_54),
.B2(n_37),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_83),
.B1(n_106),
.B2(n_94),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_99),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_54),
.B1(n_46),
.B2(n_48),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_48),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_57),
.B(n_42),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_20),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_88),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_80),
.C(n_84),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_1),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_70),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_117),
.C(n_121),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_122),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_90),
.B(n_72),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_93),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_127),
.B1(n_111),
.B2(n_103),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_70),
.C(n_69),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_74),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_69),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_131),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_94),
.B(n_103),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_42),
.C(n_73),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_135),
.C(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_134),
.B(n_93),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_77),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_20),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_20),
.B(n_28),
.C(n_21),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_140),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_142),
.C(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_101),
.C(n_104),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_111),
.B(n_114),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_114),
.B1(n_101),
.B2(n_104),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_107),
.B(n_73),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_133),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_96),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_20),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_134),
.A2(n_74),
.B1(n_42),
.B2(n_28),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_153),
.A2(n_74),
.B1(n_28),
.B2(n_21),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_154),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_116),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_137),
.A3(n_142),
.B1(n_154),
.B2(n_117),
.C1(n_125),
.C2(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_162),
.B(n_143),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_166),
.C(n_139),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_169),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_126),
.C(n_130),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_145),
.B1(n_149),
.B2(n_141),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_174),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_150),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_147),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_140),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_177),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_158),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_168),
.B(n_151),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_186),
.B(n_167),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_175),
.A2(n_171),
.B1(n_170),
.B2(n_164),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_179),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_164),
.B(n_144),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_148),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_187),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_192),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_180),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_191),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_193),
.A2(n_194),
.B(n_184),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_197),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_188),
.A3(n_189),
.B1(n_178),
.B2(n_15),
.C1(n_14),
.C2(n_21),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_5),
.B(n_7),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_21),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_199),
.B(n_6),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_202),
.B(n_203),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_8),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_10),
.Y(n_205)
);

AOI322xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_12),
.A3(n_13),
.B1(n_191),
.B2(n_152),
.C1(n_177),
.C2(n_190),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_204),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_207),
.Y(n_208)
);


endmodule