module fake_ariane_1497_n_300 (n_8, n_56, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_55, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_52, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_57, n_16, n_5, n_12, n_15, n_53, n_21, n_23, n_35, n_10, n_54, n_25, n_300);

input n_8;
input n_56;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_55;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_52;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_57;
input n_16;
input n_5;
input n_12;
input n_15;
input n_53;
input n_21;
input n_23;
input n_35;
input n_10;
input n_54;
input n_25;

output n_300;

wire n_295;
wire n_83;
wire n_233;
wire n_170;
wire n_60;
wire n_190;
wire n_289;
wire n_288;
wire n_160;
wire n_64;
wire n_180;
wire n_179;
wire n_124;
wire n_119;
wire n_167;
wire n_90;
wire n_195;
wire n_213;
wire n_294;
wire n_110;
wire n_153;
wire n_221;
wire n_197;
wire n_86;
wire n_269;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_237;
wire n_172;
wire n_69;
wire n_259;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_181;
wire n_299;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_111;
wire n_260;
wire n_242;
wire n_274;
wire n_115;
wire n_133;
wire n_265;
wire n_66;
wire n_236;
wire n_205;
wire n_272;
wire n_71;
wire n_267;
wire n_109;
wire n_208;
wire n_245;
wire n_96;
wire n_156;
wire n_281;
wire n_209;
wire n_262;
wire n_292;
wire n_291;
wire n_174;
wire n_275;
wire n_100;
wire n_283;
wire n_187;
wire n_132;
wire n_62;
wire n_225;
wire n_147;
wire n_204;
wire n_235;
wire n_210;
wire n_200;
wire n_297;
wire n_166;
wire n_253;
wire n_76;
wire n_218;
wire n_103;
wire n_79;
wire n_244;
wire n_226;
wire n_246;
wire n_271;
wire n_290;
wire n_220;
wire n_84;
wire n_247;
wire n_261;
wire n_199;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_224;
wire n_217;
wire n_240;
wire n_82;
wire n_178;
wire n_286;
wire n_131;
wire n_263;
wire n_201;
wire n_229;
wire n_70;
wire n_250;
wire n_222;
wire n_117;
wire n_139;
wire n_165;
wire n_287;
wire n_85;
wire n_130;
wire n_144;
wire n_256;
wire n_214;
wire n_227;
wire n_94;
wire n_101;
wire n_243;
wire n_284;
wire n_134;
wire n_188;
wire n_185;
wire n_249;
wire n_58;
wire n_65;
wire n_123;
wire n_212;
wire n_138;
wire n_112;
wire n_162;
wire n_264;
wire n_129;
wire n_126;
wire n_137;
wire n_255;
wire n_278;
wire n_122;
wire n_268;
wire n_257;
wire n_266;
wire n_198;
wire n_282;
wire n_148;
wire n_232;
wire n_164;
wire n_277;
wire n_157;
wire n_248;
wire n_184;
wire n_177;
wire n_135;
wire n_258;
wire n_73;
wire n_77;
wire n_293;
wire n_171;
wire n_228;
wire n_121;
wire n_93;
wire n_118;
wire n_276;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_81;
wire n_87;
wire n_206;
wire n_279;
wire n_207;
wire n_241;
wire n_254;
wire n_238;
wire n_219;
wire n_140;
wire n_191;
wire n_151;
wire n_136;
wire n_231;
wire n_192;
wire n_80;
wire n_146;
wire n_234;
wire n_230;
wire n_211;
wire n_270;
wire n_194;
wire n_97;
wire n_154;
wire n_280;
wire n_215;
wire n_252;
wire n_142;
wire n_251;
wire n_161;
wire n_285;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_296;
wire n_298;
wire n_68;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_78;
wire n_193;
wire n_63;
wire n_59;
wire n_99;
wire n_216;
wire n_155;
wire n_127;
wire n_239;
wire n_223;
wire n_273;

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

INVxp33_ASAP7_75t_SL g73 ( 
.A(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_20),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_13),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_7),
.B(n_2),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

BUFx2_ASAP7_75t_SL g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_3),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_0),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_50),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_11),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_27),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_89),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_1),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_4),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_4),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_87),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_76),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_73),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_110),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_76),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_63),
.C(n_67),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_82),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_5),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_41),
.Y(n_135)
);

AND2x4_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_106),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_94),
.B1(n_98),
.B2(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_115),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_115),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_104),
.B1(n_105),
.B2(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_103),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_101),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_99),
.Y(n_147)
);

OAI221xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_97),
.B1(n_93),
.B2(n_92),
.C(n_107),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_151)
);

AND2x4_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_6),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_117),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_124),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_134),
.B(n_133),
.Y(n_158)
);

AOI222xp33_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_118),
.B1(n_119),
.B2(n_137),
.C1(n_152),
.C2(n_148),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_119),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_133),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_118),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_152),
.Y(n_166)
);

OR2x6_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_131),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_136),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_12),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_16),
.B(n_17),
.C(n_19),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_143),
.B(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

OAI21x1_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_151),
.B(n_140),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_166),
.A2(n_143),
.B(n_140),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_28),
.B(n_29),
.Y(n_190)
);

OR2x6_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_34),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

INVx4_ASAP7_75t_SL g193 ( 
.A(n_167),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_156),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

INVx5_ASAP7_75t_SL g197 ( 
.A(n_191),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g198 ( 
.A(n_196),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_170),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_159),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_169),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_163),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_156),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_172),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_175),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_175),
.B(n_178),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_204),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

NOR3xp33_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_190),
.C(n_177),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_185),
.B(n_182),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_191),
.B1(n_192),
.B2(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_198),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_199),
.Y(n_231)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_213),
.B(n_203),
.C(n_212),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_212),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_211),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_233),
.B(n_227),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_217),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_225),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_225),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_233),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_219),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_219),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_217),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_221),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_197),
.Y(n_256)
);

OR2x6_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_226),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_251),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

NAND2x1_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_248),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_243),
.B(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_253),
.Y(n_269)
);

BUFx4f_ASAP7_75t_SL g270 ( 
.A(n_269),
.Y(n_270)
);

AOI211x1_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_245),
.B(n_252),
.C(n_205),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_264),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_243),
.B1(n_242),
.B2(n_197),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_266),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_274),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_275),
.A2(n_263),
.B1(n_257),
.B2(n_268),
.Y(n_278)
);

NOR2x1_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_262),
.Y(n_279)
);

NOR3xp33_ASAP7_75t_SL g280 ( 
.A(n_279),
.B(n_256),
.C(n_272),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

NAND4xp25_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_271),
.C(n_267),
.D(n_265),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_276),
.Y(n_283)
);

AOI221xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_258),
.B1(n_176),
.B2(n_187),
.C(n_211),
.Y(n_284)
);

OAI221xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_257),
.B1(n_197),
.B2(n_187),
.C(n_210),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_281),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_257),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_286),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_285),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_179),
.C(n_210),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_287),
.A2(n_226),
.B(n_223),
.C(n_201),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_36),
.Y(n_292)
);

OAI322xp33_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_223),
.A3(n_174),
.B1(n_171),
.B2(n_178),
.C1(n_46),
.C2(n_48),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_290),
.Y(n_294)
);

NOR4xp25_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_174),
.C(n_42),
.D(n_44),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_292),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_296)
);

AOI31xp67_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_55),
.A3(n_56),
.B(n_57),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_295),
.A2(n_157),
.B1(n_291),
.B2(n_293),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_296),
.B(n_298),
.Y(n_300)
);


endmodule