module fake_jpeg_25016_n_198 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_198);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_18),
.Y(n_50)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_17),
.C(n_16),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_60),
.C(n_17),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_50),
.B(n_61),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_31),
.B1(n_28),
.B2(n_29),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_67),
.B1(n_46),
.B2(n_16),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_28),
.B1(n_31),
.B2(n_25),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_34),
.A2(n_18),
.B(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_19),
.B1(n_25),
.B2(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_33),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_45),
.B1(n_43),
.B2(n_47),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_63),
.B1(n_22),
.B2(n_26),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_76),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_54),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_84),
.Y(n_116)
);

AND2x4_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_91),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_90),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_69),
.B1(n_70),
.B2(n_48),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx11_ASAP7_75t_SL g85 ( 
.A(n_72),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_59),
.B(n_22),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_43),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_17),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_20),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_99),
.Y(n_117)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_69),
.B1(n_70),
.B2(n_48),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_106),
.B1(n_120),
.B2(n_97),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_63),
.C(n_57),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_112),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_78),
.B(n_91),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_21),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_21),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_78),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_76),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_20),
.B1(n_2),
.B2(n_4),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_129),
.B1(n_108),
.B2(n_110),
.Y(n_150)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_126),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_119),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_124),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_134),
.B(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_79),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_73),
.B1(n_77),
.B2(n_98),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_119),
.C(n_105),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_81),
.Y(n_133)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_85),
.B(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_102),
.B(n_92),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_137),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_100),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_87),
.C(n_10),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_0),
.C(n_4),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_142),
.C(n_6),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_112),
.C(n_102),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_107),
.B(n_115),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_103),
.B1(n_115),
.B2(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_74),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_147),
.A2(n_150),
.B(n_125),
.C(n_134),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_136),
.B(n_130),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_151),
.B(n_4),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_108),
.B1(n_84),
.B2(n_6),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

OAI321xp33_ASAP7_75t_L g157 ( 
.A1(n_155),
.A2(n_132),
.A3(n_127),
.B1(n_129),
.B2(n_139),
.C(n_128),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_155),
.Y(n_171)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_164),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_165),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_146),
.B(n_9),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_5),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_142),
.C(n_140),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_13),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_171),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_147),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_156),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_145),
.B1(n_143),
.B2(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_175),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_151),
.C(n_149),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_172),
.A2(n_162),
.B(n_156),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_183),
.B(n_168),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_179),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_174),
.A2(n_159),
.B1(n_158),
.B2(n_162),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_160),
.B1(n_145),
.B2(n_156),
.Y(n_181)
);

NOR2x1_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_177),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_149),
.B(n_176),
.C(n_168),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_187),
.B(n_188),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_178),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_13),
.B(n_14),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_190),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_185),
.A2(n_183),
.B1(n_14),
.B2(n_15),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_15),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_191),
.A2(n_6),
.B(n_8),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_195),
.A2(n_192),
.B(n_196),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_190),
.Y(n_198)
);


endmodule