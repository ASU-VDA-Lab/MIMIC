module fake_ibex_1583_n_4657 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_840, n_561, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_842, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_559, n_425, n_4657);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_840;
input n_561;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_842;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4657;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_4557;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4449;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_1930;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_4632;
wire n_1080;
wire n_909;
wire n_2290;
wire n_4607;
wire n_3750;
wire n_3838;
wire n_957;
wire n_4514;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_872;
wire n_2392;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_4343;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_4353;
wire n_2598;
wire n_3819;
wire n_4648;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4421;
wire n_4179;
wire n_4601;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3411;
wire n_3025;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_4360;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_4585;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_4378;
wire n_3904;
wire n_4169;
wire n_3175;
wire n_4239;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_4477;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_4654;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_4418;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4592;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_1307;
wire n_875;
wire n_4431;
wire n_1327;
wire n_2644;
wire n_4445;
wire n_876;
wire n_3479;
wire n_1840;
wire n_2837;
wire n_3211;
wire n_4652;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_4470;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_1636;
wire n_939;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3753;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4423;
wire n_4584;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_4578;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_4304;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_4382;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_4450;
wire n_3969;
wire n_4467;
wire n_1081;
wire n_4437;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4491;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_4569;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3949;
wire n_3507;
wire n_3884;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2436;
wire n_2333;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_3711;
wire n_1595;
wire n_2164;
wire n_4267;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_4389;
wire n_4510;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_4312;
wire n_1955;
wire n_3668;
wire n_3699;
wire n_4567;
wire n_917;
wire n_4556;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_4214;
wire n_1313;
wire n_3973;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_4430;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_4650;
wire n_1645;
wire n_3186;
wire n_4433;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_4428;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_4563;
wire n_3809;
wire n_979;
wire n_4503;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4517;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_4511;
wire n_1007;
wire n_2253;
wire n_4479;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_4422;
wire n_1219;
wire n_4513;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_4610;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_4481;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_971;
wire n_1326;
wire n_4444;
wire n_1350;
wire n_3627;
wire n_906;
wire n_4499;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1764;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_4595;
wire n_2541;
wire n_4598;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_4553;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_4533;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4455;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4518;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_4480;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_4548;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_4535;
wire n_1447;
wire n_2451;
wire n_2166;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_4252;
wire n_4505;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_4577;
wire n_2292;
wire n_3573;
wire n_4604;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_4398;
wire n_3516;
wire n_1298;
wire n_1844;
wire n_4522;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_4476;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_4615;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4103;
wire n_3583;
wire n_2019;
wire n_4126;
wire n_1407;
wire n_3282;
wire n_4435;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_4649;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_1543;
wire n_4653;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_4568;
wire n_4359;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4549;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_4623;
wire n_1041;
wire n_2766;
wire n_4156;
wire n_2828;
wire n_3754;
wire n_4411;
wire n_1964;
wire n_3756;
wire n_4523;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_4489;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_4419;
wire n_1583;
wire n_3520;
wire n_4404;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_4571;
wire n_959;
wire n_1106;
wire n_1312;
wire n_4655;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_4570;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_4494;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4122;
wire n_4542;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_4572;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_4374;
wire n_1140;
wire n_1985;
wire n_4375;
wire n_4501;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_4403;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_4230;
wire n_3849;
wire n_965;
wire n_1109;
wire n_4402;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4469;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_4558;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_4460;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4504;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_4527;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_4033;
wire n_3855;
wire n_4485;
wire n_4608;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_1236;
wire n_3364;
wire n_4384;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_4537;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4323;
wire n_4407;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_4646;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_4462;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_4540;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_4490;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_4362;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_4414;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_4409;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_4525;
wire n_3396;
wire n_4190;
wire n_4011;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_4443;
wire n_1682;
wire n_4151;
wire n_4625;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_4554;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_4424;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_4596;
wire n_4415;
wire n_1345;
wire n_4215;
wire n_4456;
wire n_4587;
wire n_4315;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_4492;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_4500;
wire n_4559;
wire n_1395;
wire n_1115;
wire n_998;
wire n_1729;
wire n_2551;
wire n_4641;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_882;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_3829;
wire n_4579;
wire n_1864;
wire n_4624;
wire n_943;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_2570;
wire n_4051;
wire n_4321;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_4552;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1400;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2842;
wire n_3070;
wire n_2711;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4416;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4640;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2612;
wire n_2193;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4561;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_4642;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_3557;
wire n_1746;
wire n_1439;
wire n_2263;
wire n_2352;
wire n_2212;
wire n_2716;
wire n_3495;
wire n_2185;
wire n_4141;
wire n_4614;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_4117;
wire n_3999;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3498;
wire n_2986;
wire n_3238;
wire n_4520;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_4496;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4566;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_4647;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4636;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1185;
wire n_1683;
wire n_4256;
wire n_3575;
wire n_4454;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_4278;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_4609;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_4458;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_4276;
wire n_4612;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3927;
wire n_3902;
wire n_2422;
wire n_4185;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_920;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_4441;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_991;
wire n_1331;
wire n_1223;
wire n_961;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_4536;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_4633;
wire n_1950;
wire n_4497;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_996;
wire n_4593;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_2619;
wire n_3289;
wire n_1174;
wire n_4512;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_4483;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4488;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4142;
wire n_4183;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1458;
wire n_1694;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_4621;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_4123;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_4619;
wire n_4645;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3908;
wire n_3616;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_4286;
wire n_4429;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_4438;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_4638;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_4498;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_4001;
wire n_3427;
wire n_3669;
wire n_1348;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4377;
wire n_4099;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_3899;
wire n_1617;
wire n_1839;
wire n_3930;
wire n_4149;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_4118;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_4319;
wire n_4637;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_4543;
wire n_4466;
wire n_2688;
wire n_2881;
wire n_4643;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_4603;
wire n_2268;
wire n_2320;
wire n_2237;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_4417;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4212;
wire n_4022;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_3162;
wire n_2984;
wire n_4436;
wire n_4599;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_4538;
wire n_3096;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_4616;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4288;
wire n_4068;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_4434;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_4586;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_4622;
wire n_3273;
wire n_4367;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_4282;
wire n_1630;
wire n_3408;
wire n_4475;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_4588;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3647;
wire n_3623;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_4410;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_4440;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3649;
wire n_1838;
wire n_3604;
wire n_3540;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_4529;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2576;
wire n_2348;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4162;
wire n_4200;
wire n_4408;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_4575;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_4620;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_4439;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_885;
wire n_1530;
wire n_4111;
wire n_3215;
wire n_3413;
wire n_877;
wire n_4580;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_4565;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_4581;
wire n_1288;
wire n_4058;
wire n_4487;
wire n_4618;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4519;
wire n_4148;
wire n_897;
wire n_1622;
wire n_2757;
wire n_4611;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_4541;
wire n_4515;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_4530;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_4463;
wire n_4591;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1809;
wire n_1206;
wire n_2367;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_4265;
wire n_3062;
wire n_4524;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4628;
wire n_4017;
wire n_1547;
wire n_1542;
wire n_1586;
wire n_1362;
wire n_946;
wire n_3497;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4597;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_4574;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1887;
wire n_1212;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_4555;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_4562;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_4453;
wire n_1098;
wire n_4474;
wire n_1366;
wire n_1518;
wire n_4350;
wire n_4380;
wire n_1361;
wire n_1187;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2653;
wire n_3102;
wire n_2872;
wire n_3173;
wire n_4281;
wire n_4345;
wire n_2411;
wire n_4478;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_4473;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_4464;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_4605;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_4546;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1572;
wire n_1635;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2929;
wire n_2701;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_4045;
wire n_4432;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_4405;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3791;
wire n_3742;
wire n_3655;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4461;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_4516;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_4528;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_4502;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_914;
wire n_3992;
wire n_4147;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_4471;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3547;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4386;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_4547;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3831;
wire n_3296;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_2005;
wire n_1284;
wire n_4482;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_4406;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3430;
wire n_3200;
wire n_4493;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1488;
wire n_1193;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3483;
wire n_1074;
wire n_3380;
wire n_3225;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3823;
wire n_3369;
wire n_3606;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_4634;
wire n_4644;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_1022;
wire n_4412;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_4560;
wire n_3285;
wire n_3160;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3124;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3286;
wire n_4038;
wire n_1092;
wire n_4472;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_4639;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_4635;
wire n_4521;
wire n_1230;
wire n_4459;
wire n_1516;
wire n_1027;
wire n_4551;
wire n_3893;
wire n_4484;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2357;
wire n_2303;
wire n_2618;
wire n_2855;
wire n_4448;
wire n_3938;
wire n_4354;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_4401;
wire n_4532;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_4413;
wire n_1757;
wire n_4627;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2560;
wire n_2302;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_2802;
wire n_3189;
wire n_4544;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1158;
wire n_1974;
wire n_2988;
wire n_3945;
wire n_4275;
wire n_1882;
wire n_4046;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_4589;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_4468;
wire n_1736;
wire n_4617;
wire n_4442;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_4594;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_4613;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_4629;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_4539;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_4486;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3933;
wire n_2262;
wire n_3562;
wire n_4188;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2917;
wire n_2726;
wire n_3873;
wire n_4506;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4226;
wire n_1551;
wire n_4153;
wire n_3793;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_4327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4251;
wire n_4106;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_4465;
wire n_1355;
wire n_4452;
wire n_3691;
wire n_2544;
wire n_3193;
wire n_4534;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_4590;
wire n_2915;
wire n_1579;
wire n_4446;
wire n_1280;
wire n_4602;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_4576;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_4606;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_4508;
wire n_3851;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_4425;
wire n_3980;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_1655;
wire n_984;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_196),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_538),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_172),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_759),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_406),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_861),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_125),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_570),
.Y(n_871)
);

CKINVDCx16_ASAP7_75t_R g872 ( 
.A(n_111),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_525),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_795),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_721),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_455),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_709),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_588),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_56),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_792),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_176),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_399),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_118),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_758),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_539),
.B(n_415),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_838),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_29),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_183),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_784),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_433),
.Y(n_890)
);

BUFx8_ASAP7_75t_SL g891 ( 
.A(n_139),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_258),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_506),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_341),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_313),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_162),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_831),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_206),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_143),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_141),
.Y(n_900)
);

BUFx5_ASAP7_75t_L g901 ( 
.A(n_38),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_744),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_800),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_290),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_653),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_188),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_737),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_468),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_837),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_370),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_438),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_680),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_526),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_751),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_803),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_195),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_176),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_737),
.Y(n_918)
);

CKINVDCx14_ASAP7_75t_R g919 ( 
.A(n_513),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_788),
.B(n_193),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_179),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_366),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_191),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_658),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_526),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_814),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_328),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_760),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_598),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_54),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_364),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_678),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_328),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_825),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_485),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_717),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_292),
.Y(n_937)
);

BUFx5_ASAP7_75t_L g938 ( 
.A(n_273),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_476),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_396),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_478),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_468),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_279),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_522),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_357),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_442),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_318),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_853),
.Y(n_948)
);

BUFx10_ASAP7_75t_L g949 ( 
.A(n_310),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_796),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_367),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_441),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_824),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_840),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_432),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_820),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_859),
.Y(n_957)
);

CKINVDCx16_ASAP7_75t_R g958 ( 
.A(n_242),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_295),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_112),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_214),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_177),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_718),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_613),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_618),
.Y(n_965)
);

BUFx5_ASAP7_75t_L g966 ( 
.A(n_840),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_713),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_727),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_813),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_704),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_610),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_298),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_773),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_624),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_815),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_346),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_677),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_694),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_498),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_69),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_839),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_97),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_34),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_832),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_785),
.Y(n_985)
);

BUFx2_ASAP7_75t_SL g986 ( 
.A(n_535),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_246),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_191),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_361),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_509),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_793),
.Y(n_991)
);

CKINVDCx16_ASAP7_75t_R g992 ( 
.A(n_99),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_674),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_716),
.Y(n_994)
);

CKINVDCx20_ASAP7_75t_R g995 ( 
.A(n_549),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_373),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_639),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_219),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_218),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_175),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_365),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_792),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_630),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_81),
.Y(n_1004)
);

BUFx10_ASAP7_75t_L g1005 ( 
.A(n_143),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_95),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_509),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_471),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_110),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_599),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_338),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_514),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_811),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_558),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_332),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_832),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_224),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_608),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_835),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_241),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_385),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_772),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_29),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_8),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_63),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_166),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_279),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_820),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_349),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_507),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_64),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_266),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_281),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_326),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_38),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_171),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_454),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_611),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_856),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_834),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_836),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_583),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_482),
.Y(n_1043)
);

BUFx10_ASAP7_75t_L g1044 ( 
.A(n_662),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_182),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_582),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_475),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_704),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_789),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_692),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_431),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_134),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_182),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_102),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_31),
.B(n_812),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_698),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_493),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_539),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_657),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_296),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_753),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_188),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_522),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_18),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_140),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_401),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_536),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_297),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_45),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_800),
.Y(n_1070)
);

BUFx10_ASAP7_75t_L g1071 ( 
.A(n_364),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_578),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_394),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_629),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_149),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_495),
.Y(n_1076)
);

BUFx8_ASAP7_75t_SL g1077 ( 
.A(n_782),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_667),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_781),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_447),
.Y(n_1080)
);

CKINVDCx16_ASAP7_75t_R g1081 ( 
.A(n_834),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_829),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_257),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_766),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_549),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_313),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_58),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_714),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_794),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_649),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_49),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_310),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_190),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_236),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_283),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_360),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_586),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_265),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_717),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_351),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_322),
.Y(n_1101)
);

CKINVDCx16_ASAP7_75t_R g1102 ( 
.A(n_390),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_559),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_149),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_130),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_186),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_200),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_288),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_305),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_288),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_844),
.Y(n_1111)
);

CKINVDCx16_ASAP7_75t_R g1112 ( 
.A(n_686),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_28),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_590),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_818),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_846),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_754),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_412),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_512),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_99),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_808),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_157),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_42),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_530),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_98),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_32),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_476),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_773),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_69),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_9),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_360),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_265),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_826),
.Y(n_1133)
);

NOR2xp67_ASAP7_75t_L g1134 ( 
.A(n_260),
.B(n_63),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_561),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_845),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_797),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_485),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_448),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_569),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_348),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_625),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_44),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_489),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_379),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_216),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_103),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_64),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_776),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_828),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_62),
.Y(n_1151)
);

CKINVDCx16_ASAP7_75t_R g1152 ( 
.A(n_504),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_329),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_659),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_657),
.Y(n_1155)
);

INVxp67_ASAP7_75t_SL g1156 ( 
.A(n_710),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_603),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_453),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_693),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_557),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_30),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_64),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_495),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_658),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_293),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_204),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_124),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_471),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_757),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_76),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_745),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_33),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_806),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_78),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_249),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_828),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_701),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_660),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_786),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_685),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_807),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_801),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_706),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_788),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_98),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_367),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_683),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_780),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_375),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_789),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_96),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_822),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_165),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_506),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_777),
.Y(n_1195)
);

BUFx10_ASAP7_75t_L g1196 ( 
.A(n_290),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_309),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_432),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_612),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_696),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_453),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_247),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_554),
.Y(n_1203)
);

BUFx10_ASAP7_75t_L g1204 ( 
.A(n_635),
.Y(n_1204)
);

CKINVDCx20_ASAP7_75t_R g1205 ( 
.A(n_237),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_298),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_825),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_799),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_173),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_285),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_716),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_823),
.Y(n_1212)
);

INVxp67_ASAP7_75t_L g1213 ( 
.A(n_601),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_119),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_88),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_842),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_830),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_33),
.Y(n_1218)
);

BUFx10_ASAP7_75t_L g1219 ( 
.A(n_546),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_819),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_804),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_390),
.B(n_441),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_847),
.Y(n_1223)
);

NOR2xp67_ASAP7_75t_L g1224 ( 
.A(n_11),
.B(n_161),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_119),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_600),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_821),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_31),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_190),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_150),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_220),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_349),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_735),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_841),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_791),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_482),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_L g1237 ( 
.A(n_100),
.B(n_409),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_402),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_13),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_464),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_738),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_541),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_805),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_356),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_639),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_129),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_492),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_27),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_816),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_616),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_707),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_122),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_643),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_350),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_325),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_465),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_153),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_632),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_455),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_490),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_283),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_843),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_548),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_101),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_266),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_280),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_602),
.Y(n_1267)
);

CKINVDCx16_ASAP7_75t_R g1268 ( 
.A(n_748),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_319),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_802),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_493),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_96),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_778),
.Y(n_1273)
);

CKINVDCx14_ASAP7_75t_R g1274 ( 
.A(n_417),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_32),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_95),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_779),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_538),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_745),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_60),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_51),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_809),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_809),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_761),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_263),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_253),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_726),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_584),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_827),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_484),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_568),
.Y(n_1291)
);

BUFx5_ASAP7_75t_L g1292 ( 
.A(n_589),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_641),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_833),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_781),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_790),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_786),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_155),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_420),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_49),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_805),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_41),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_561),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_725),
.Y(n_1304)
);

NOR2xp67_ASAP7_75t_L g1305 ( 
.A(n_531),
.B(n_796),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_334),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_39),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_817),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_0),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_232),
.Y(n_1310)
);

BUFx10_ASAP7_75t_L g1311 ( 
.A(n_300),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_783),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_92),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_363),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_798),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_231),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_810),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_667),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_489),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_604),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_167),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_52),
.Y(n_1322)
);

BUFx5_ASAP7_75t_L g1323 ( 
.A(n_187),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_787),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_41),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_267),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_736),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_524),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_775),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_118),
.Y(n_1330)
);

INVxp67_ASAP7_75t_SL g1331 ( 
.A(n_345),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_171),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_498),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_3),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_403),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_408),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_309),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_130),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_28),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_553),
.Y(n_1340)
);

INVx5_ASAP7_75t_L g1341 ( 
.A(n_1064),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1004),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_919),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1006),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_864),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_864),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_864),
.Y(n_1347)
);

BUFx12f_ASAP7_75t_L g1348 ( 
.A(n_949),
.Y(n_1348)
);

AND2x6_ASAP7_75t_L g1349 ( 
.A(n_1129),
.B(n_0),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_938),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1087),
.B(n_0),
.Y(n_1351)
);

BUFx12f_ASAP7_75t_L g1352 ( 
.A(n_949),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1280),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_864),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1129),
.B(n_1),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_938),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_904),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_906),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1022),
.B(n_1),
.Y(n_1359)
);

OAI22x1_ASAP7_75t_SL g1360 ( 
.A1(n_1035),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_1360)
);

AND2x2_ASAP7_75t_SL g1361 ( 
.A(n_958),
.B(n_2),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_949),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1075),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_980),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_919),
.Y(n_1365)
);

BUFx8_ASAP7_75t_L g1366 ( 
.A(n_1033),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_904),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_904),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1133),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1069),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1274),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_938),
.Y(n_1372)
);

INVx6_ASAP7_75t_L g1373 ( 
.A(n_1005),
.Y(n_1373)
);

AOI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1274),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1005),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1163),
.B(n_4),
.Y(n_1376)
);

CKINVDCx6p67_ASAP7_75t_R g1377 ( 
.A(n_1005),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1223),
.B(n_4),
.Y(n_1378)
);

AOI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1339),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_1379)
);

NOR2xp67_ASAP7_75t_L g1380 ( 
.A(n_918),
.B(n_5),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1130),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1247),
.B(n_5),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1279),
.B(n_6),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_909),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_879),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1143),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1148),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1162),
.Y(n_1388)
);

OAI22x1_ASAP7_75t_SL g1389 ( 
.A1(n_1061),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1389)
);

BUFx12f_ASAP7_75t_L g1390 ( 
.A(n_1044),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_887),
.A2(n_7),
.B(n_8),
.Y(n_1391)
);

INVx6_ASAP7_75t_L g1392 ( 
.A(n_1044),
.Y(n_1392)
);

BUFx12f_ASAP7_75t_L g1393 ( 
.A(n_1044),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1191),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1215),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_938),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1248),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_887),
.A2(n_9),
.B(n_10),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1075),
.B(n_9),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1309),
.A2(n_10),
.B(n_11),
.Y(n_1400)
);

BUFx12f_ASAP7_75t_L g1401 ( 
.A(n_1071),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1071),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1061),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_1403)
);

INVx6_ASAP7_75t_L g1404 ( 
.A(n_1071),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_922),
.B(n_12),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_891),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_904),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_938),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_872),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_938),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1125),
.B(n_14),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1196),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_975),
.B(n_14),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1196),
.Y(n_1414)
);

OAI22x1_ASAP7_75t_SL g1415 ( 
.A1(n_1231),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_914),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1171),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1196),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1272),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_901),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1185),
.B(n_15),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_948),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_891),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_992),
.B(n_15),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1275),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_914),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1302),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_930),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1077),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1125),
.B(n_19),
.Y(n_1430)
);

INVx5_ASAP7_75t_L g1431 ( 
.A(n_1064),
.Y(n_1431)
);

CKINVDCx16_ASAP7_75t_R g1432 ( 
.A(n_1081),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1309),
.A2(n_19),
.B(n_20),
.Y(n_1433)
);

INVx5_ASAP7_75t_L g1434 ( 
.A(n_1064),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1307),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1201),
.B(n_20),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1201),
.B(n_21),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1322),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1064),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_901),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_966),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1371),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1371),
.B(n_1102),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1406),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1344),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1385),
.B(n_1353),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1423),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1429),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1342),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1343),
.B(n_901),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1432),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1363),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1355),
.Y(n_1453)
);

NAND2xp33_ASAP7_75t_R g1454 ( 
.A(n_1365),
.B(n_983),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1345),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1377),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1409),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1358),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1348),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1411),
.Y(n_1460)
);

BUFx10_ASAP7_75t_L g1461 ( 
.A(n_1373),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1430),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1352),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1375),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1436),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1390),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1393),
.Y(n_1467)
);

XNOR2xp5_ASAP7_75t_L g1468 ( 
.A(n_1361),
.B(n_1231),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1437),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1384),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1422),
.B(n_925),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1417),
.B(n_1112),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1401),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1439),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1345),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1350),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1369),
.B(n_1152),
.Y(n_1477)
);

INVx2_ASAP7_75t_SL g1478 ( 
.A(n_1373),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1366),
.Y(n_1479)
);

INVxp33_ASAP7_75t_L g1480 ( 
.A(n_1424),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1392),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1392),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1356),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_R g1484 ( 
.A(n_1362),
.B(n_1268),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1372),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1364),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1404),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1389),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1402),
.B(n_901),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1415),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1360),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1414),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1418),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_R g1494 ( 
.A(n_1349),
.B(n_1023),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1396),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_1378),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1408),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1351),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1346),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1374),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1376),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1412),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1346),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1370),
.Y(n_1504)
);

CKINVDCx16_ASAP7_75t_R g1505 ( 
.A(n_1359),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1381),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1398),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1410),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1386),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1383),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1387),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1388),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1394),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1403),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1395),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1382),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1397),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1349),
.Y(n_1518)
);

NAND2xp33_ASAP7_75t_R g1519 ( 
.A(n_1391),
.B(n_1024),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1419),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1349),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1405),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1425),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1413),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1347),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1400),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1433),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1379),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1428),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_R g1530 ( 
.A(n_1427),
.B(n_1025),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1435),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1421),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1438),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1441),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_1391),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1420),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1440),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1380),
.B(n_1204),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1440),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1341),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_R g1541 ( 
.A(n_1431),
.B(n_1031),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1431),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1347),
.B(n_1313),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_R g1544 ( 
.A(n_1434),
.B(n_1091),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1434),
.B(n_1354),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1434),
.Y(n_1546)
);

NAND2xp33_ASAP7_75t_SL g1547 ( 
.A(n_1354),
.B(n_1055),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1357),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1357),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1367),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1367),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1368),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1407),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1407),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1416),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1416),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1426),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1426),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1406),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1406),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1371),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1406),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1406),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1385),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1371),
.B(n_1204),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1342),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1344),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1344),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1363),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1406),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1345),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1399),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1363),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1406),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1399),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1344),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1344),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1406),
.Y(n_1578)
);

CKINVDCx16_ASAP7_75t_R g1579 ( 
.A(n_1432),
.Y(n_1579)
);

INVxp67_ASAP7_75t_SL g1580 ( 
.A(n_1371),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1406),
.Y(n_1581)
);

BUFx10_ASAP7_75t_L g1582 ( 
.A(n_1373),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1385),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1406),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1406),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1406),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1371),
.B(n_1204),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1371),
.B(n_1113),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1345),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_1342),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_1342),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1406),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_R g1593 ( 
.A(n_1406),
.B(n_1123),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1344),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1363),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1406),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_R g1597 ( 
.A(n_1406),
.B(n_1126),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1344),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1406),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1406),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1406),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1344),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1385),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1399),
.Y(n_1604)
);

CKINVDCx16_ASAP7_75t_R g1605 ( 
.A(n_1432),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1406),
.Y(n_1606)
);

AND3x2_ASAP7_75t_L g1607 ( 
.A(n_1385),
.B(n_1331),
.C(n_1156),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1406),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1406),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1406),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1406),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1344),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_R g1613 ( 
.A(n_1406),
.B(n_1151),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1364),
.B(n_966),
.Y(n_1614)
);

INVxp67_ASAP7_75t_SL g1615 ( 
.A(n_1371),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1458),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1543),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1530),
.B(n_1161),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1531),
.B(n_1170),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1507),
.Y(n_1620)
);

BUFx2_ASAP7_75t_R g1621 ( 
.A(n_1479),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1518),
.B(n_1325),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1452),
.Y(n_1623)
);

NAND2xp33_ASAP7_75t_L g1624 ( 
.A(n_1521),
.B(n_966),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1526),
.Y(n_1625)
);

NAND2xp33_ASAP7_75t_SL g1626 ( 
.A(n_1484),
.B(n_1334),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1493),
.B(n_972),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1445),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1493),
.B(n_1213),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1522),
.B(n_1172),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1535),
.A2(n_1281),
.B1(n_1218),
.B2(n_1228),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1588),
.B(n_970),
.Y(n_1632)
);

NOR3xp33_ASAP7_75t_L g1633 ( 
.A(n_1579),
.B(n_997),
.C(n_865),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1472),
.B(n_1219),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1478),
.B(n_1013),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1532),
.B(n_1174),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1567),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_SL g1638 ( 
.A(n_1583),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1568),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1576),
.Y(n_1640)
);

NAND2x1_ASAP7_75t_L g1641 ( 
.A(n_1486),
.B(n_1281),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1524),
.B(n_1239),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1453),
.B(n_1276),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1569),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1501),
.B(n_1300),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1461),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1577),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1516),
.B(n_966),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1594),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1461),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1598),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1602),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1460),
.B(n_1281),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1446),
.B(n_1100),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1612),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1572),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1504),
.B(n_966),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_SL g1658 ( 
.A(n_1564),
.B(n_1077),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1462),
.B(n_1465),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1506),
.B(n_966),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1469),
.B(n_1281),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1509),
.B(n_1511),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1572),
.Y(n_1663)
);

BUFx6f_ASAP7_75t_L g1664 ( 
.A(n_1546),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1573),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1545),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1575),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1512),
.B(n_1292),
.Y(n_1668)
);

OR2x6_ASAP7_75t_L g1669 ( 
.A(n_1442),
.B(n_1561),
.Y(n_1669)
);

NOR3xp33_ASAP7_75t_L g1670 ( 
.A(n_1605),
.B(n_1094),
.C(n_1003),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1536),
.B(n_914),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1575),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1513),
.B(n_1292),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1502),
.B(n_867),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1515),
.B(n_1292),
.Y(n_1675)
);

AND2x6_ASAP7_75t_L g1676 ( 
.A(n_1519),
.B(n_1565),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1604),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1517),
.B(n_1292),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1595),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1604),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1614),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1614),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1537),
.B(n_957),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1498),
.B(n_869),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1520),
.B(n_1292),
.Y(n_1685)
);

OR2x6_ASAP7_75t_L g1686 ( 
.A(n_1603),
.B(n_1443),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1587),
.B(n_870),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1523),
.B(n_1292),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1538),
.B(n_1134),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1580),
.B(n_1323),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1615),
.B(n_1539),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1471),
.B(n_1323),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1489),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1477),
.B(n_1219),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1480),
.B(n_1219),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1450),
.B(n_1323),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_SL g1697 ( 
.A(n_1456),
.B(n_1459),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1481),
.B(n_1582),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1582),
.B(n_1505),
.Y(n_1699)
);

NAND2x1p5_ASAP7_75t_L g1700 ( 
.A(n_1463),
.B(n_920),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1547),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1474),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1476),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1483),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1482),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1485),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1495),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1497),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1510),
.B(n_1323),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1545),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1492),
.B(n_957),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1508),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1534),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1487),
.B(n_1541),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1544),
.B(n_1233),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1496),
.B(n_1233),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1555),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1470),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1607),
.B(n_1314),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1556),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1557),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1540),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1542),
.B(n_1328),
.Y(n_1723)
);

NOR3xp33_ASAP7_75t_L g1724 ( 
.A(n_1528),
.B(n_1199),
.C(n_1187),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1593),
.B(n_957),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1550),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_SL g1727 ( 
.A(n_1451),
.Y(n_1727)
);

NOR2x1_ASAP7_75t_L g1728 ( 
.A(n_1549),
.B(n_1558),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1464),
.B(n_1466),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1551),
.Y(n_1730)
);

NAND2xp33_ASAP7_75t_L g1731 ( 
.A(n_1467),
.B(n_957),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1597),
.B(n_988),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1552),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1613),
.B(n_988),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1473),
.B(n_988),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1529),
.B(n_876),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_SL g1737 ( 
.A(n_1444),
.B(n_988),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1514),
.B(n_881),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1533),
.A2(n_868),
.B1(n_873),
.B2(n_866),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1554),
.B(n_882),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1500),
.B(n_886),
.Y(n_1741)
);

NOR2xp67_ASAP7_75t_L g1742 ( 
.A(n_1447),
.B(n_21),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1468),
.B(n_1311),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1548),
.B(n_888),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1553),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1454),
.B(n_889),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1448),
.B(n_890),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1455),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1559),
.B(n_893),
.Y(n_1749)
);

INVx2_ASAP7_75t_SL g1750 ( 
.A(n_1449),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1560),
.B(n_895),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1455),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1475),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1562),
.B(n_898),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1563),
.B(n_1021),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1570),
.B(n_899),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1574),
.B(n_902),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1475),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1578),
.B(n_905),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1475),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1499),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1499),
.Y(n_1762)
);

NAND2xp33_ASAP7_75t_L g1763 ( 
.A(n_1581),
.B(n_1021),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1503),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1503),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1584),
.B(n_907),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1585),
.B(n_911),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1586),
.B(n_912),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1457),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1592),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1503),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1596),
.B(n_913),
.Y(n_1772)
);

INVx4_ASAP7_75t_L g1773 ( 
.A(n_1599),
.Y(n_1773)
);

NOR2xp67_ASAP7_75t_L g1774 ( 
.A(n_1600),
.B(n_22),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1525),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1601),
.B(n_916),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1571),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1611),
.B(n_917),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1606),
.B(n_923),
.Y(n_1779)
);

NAND2xp33_ASAP7_75t_L g1780 ( 
.A(n_1608),
.B(n_1021),
.Y(n_1780)
);

NOR3xp33_ASAP7_75t_L g1781 ( 
.A(n_1488),
.B(n_1225),
.C(n_1211),
.Y(n_1781)
);

OA21x2_ASAP7_75t_L g1782 ( 
.A1(n_1609),
.A2(n_875),
.B(n_874),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1571),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1589),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1610),
.B(n_1021),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_SL g1786 ( 
.A(n_1490),
.Y(n_1786)
);

INVx4_ASAP7_75t_L g1787 ( 
.A(n_1589),
.Y(n_1787)
);

NOR2xp67_ASAP7_75t_L g1788 ( 
.A(n_1491),
.B(n_22),
.Y(n_1788)
);

NOR3xp33_ASAP7_75t_L g1789 ( 
.A(n_1566),
.B(n_1277),
.C(n_1245),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1589),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1590),
.A2(n_883),
.B1(n_884),
.B2(n_878),
.Y(n_1791)
);

INVx2_ASAP7_75t_SL g1792 ( 
.A(n_1591),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_SL g1793 ( 
.A(n_1583),
.Y(n_1793)
);

BUFx5_ASAP7_75t_L g1794 ( 
.A(n_1507),
.Y(n_1794)
);

NAND2xp33_ASAP7_75t_L g1795 ( 
.A(n_1494),
.B(n_1115),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1543),
.Y(n_1796)
);

NAND3xp33_ASAP7_75t_L g1797 ( 
.A(n_1532),
.B(n_926),
.C(n_924),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1522),
.B(n_929),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1458),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1493),
.B(n_933),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1522),
.B(n_934),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1522),
.B(n_935),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1527),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1543),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_SL g1805 ( 
.A(n_1494),
.B(n_1115),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1493),
.B(n_936),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1522),
.B(n_940),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1522),
.B(n_946),
.Y(n_1808)
);

INVx2_ASAP7_75t_SL g1809 ( 
.A(n_1461),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1458),
.B(n_1311),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1493),
.B(n_947),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1543),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1493),
.B(n_950),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1522),
.B(n_951),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1493),
.B(n_952),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1543),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1522),
.B(n_959),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1543),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1522),
.B(n_962),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1522),
.B(n_964),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1522),
.B(n_968),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1493),
.B(n_969),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1522),
.B(n_971),
.Y(n_1823)
);

NOR2xp67_ASAP7_75t_L g1824 ( 
.A(n_1459),
.B(n_23),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1522),
.B(n_976),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1522),
.B(n_978),
.Y(n_1826)
);

NAND2xp33_ASAP7_75t_L g1827 ( 
.A(n_1494),
.B(n_1115),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1522),
.B(n_982),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1494),
.B(n_1115),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1522),
.B(n_985),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1494),
.B(n_1120),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1543),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1522),
.B(n_987),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1494),
.B(n_1120),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1522),
.B(n_990),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1493),
.B(n_991),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1522),
.B(n_993),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_SL g1838 ( 
.A(n_1494),
.B(n_1120),
.Y(n_1838)
);

NOR2xp67_ASAP7_75t_SL g1839 ( 
.A(n_1518),
.B(n_1330),
.Y(n_1839)
);

CKINVDCx20_ASAP7_75t_R g1840 ( 
.A(n_1470),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_1493),
.B(n_998),
.Y(n_1841)
);

OR2x6_ASAP7_75t_L g1842 ( 
.A(n_1583),
.B(n_986),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_SL g1843 ( 
.A(n_1518),
.B(n_1263),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1543),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_SL g1845 ( 
.A(n_1518),
.B(n_1263),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1522),
.B(n_1000),
.Y(n_1846)
);

BUFx3_ASAP7_75t_L g1847 ( 
.A(n_1583),
.Y(n_1847)
);

NAND2xp33_ASAP7_75t_L g1848 ( 
.A(n_1494),
.B(n_1140),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1527),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1630),
.B(n_1001),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1616),
.B(n_871),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1620),
.B(n_1002),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1628),
.Y(n_1853)
);

NOR2xp67_ASAP7_75t_L g1854 ( 
.A(n_1773),
.B(n_23),
.Y(n_1854)
);

BUFx3_ASAP7_75t_L g1855 ( 
.A(n_1840),
.Y(n_1855)
);

INVx4_ASAP7_75t_L g1856 ( 
.A(n_1620),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1620),
.B(n_1007),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1637),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1639),
.Y(n_1859)
);

NAND2xp33_ASAP7_75t_L g1860 ( 
.A(n_1625),
.B(n_1008),
.Y(n_1860)
);

BUFx4f_ASAP7_75t_L g1861 ( 
.A(n_1842),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1642),
.B(n_1010),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1645),
.B(n_1012),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1640),
.Y(n_1864)
);

NAND2xp33_ASAP7_75t_SL g1865 ( 
.A(n_1625),
.B(n_1329),
.Y(n_1865)
);

NAND3xp33_ASAP7_75t_L g1866 ( 
.A(n_1789),
.B(n_1016),
.C(n_1014),
.Y(n_1866)
);

AND2x4_ASAP7_75t_SL g1867 ( 
.A(n_1669),
.B(n_877),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1681),
.B(n_1017),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1682),
.B(n_1020),
.Y(n_1869)
);

A2O1A1Ixp33_ASAP7_75t_L g1870 ( 
.A1(n_1647),
.A2(n_1224),
.B(n_885),
.C(n_1222),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1676),
.A2(n_896),
.B1(n_897),
.B2(n_894),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1662),
.B(n_1028),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1799),
.B(n_1694),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1649),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1625),
.B(n_1029),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1794),
.B(n_1030),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1651),
.B(n_1652),
.Y(n_1877)
);

INVx4_ASAP7_75t_L g1878 ( 
.A(n_1669),
.Y(n_1878)
);

NAND2x1p5_ASAP7_75t_L g1879 ( 
.A(n_1847),
.B(n_1237),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1803),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1794),
.B(n_1032),
.Y(n_1881)
);

BUFx2_ASAP7_75t_L g1882 ( 
.A(n_1718),
.Y(n_1882)
);

OR2x6_ASAP7_75t_L g1883 ( 
.A(n_1842),
.B(n_1305),
.Y(n_1883)
);

BUFx3_ASAP7_75t_L g1884 ( 
.A(n_1699),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1655),
.B(n_1034),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1798),
.B(n_1037),
.Y(n_1886)
);

BUFx8_ASAP7_75t_L g1887 ( 
.A(n_1727),
.Y(n_1887)
);

NAND2xp33_ASAP7_75t_L g1888 ( 
.A(n_1794),
.B(n_1040),
.Y(n_1888)
);

AND2x6_ASAP7_75t_SL g1889 ( 
.A(n_1729),
.B(n_885),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1686),
.B(n_927),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1801),
.B(n_1041),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1802),
.B(n_1043),
.Y(n_1892)
);

INVx2_ASAP7_75t_SL g1893 ( 
.A(n_1698),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1686),
.B(n_953),
.Y(n_1894)
);

INVx3_ASAP7_75t_L g1895 ( 
.A(n_1638),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1807),
.B(n_1047),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1794),
.B(n_1048),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1646),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1808),
.B(n_1054),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1634),
.B(n_960),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1814),
.B(n_1057),
.Y(n_1901)
);

INVx3_ASAP7_75t_L g1902 ( 
.A(n_1638),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1656),
.Y(n_1903)
);

OR2x6_ASAP7_75t_L g1904 ( 
.A(n_1750),
.B(n_880),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1817),
.B(n_1058),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1663),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1849),
.A2(n_908),
.B(n_900),
.Y(n_1907)
);

OR2x6_ASAP7_75t_L g1908 ( 
.A(n_1792),
.B(n_880),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1728),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1667),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1793),
.Y(n_1911)
);

HB1xp67_ASAP7_75t_L g1912 ( 
.A(n_1793),
.Y(n_1912)
);

INVx3_ASAP7_75t_L g1913 ( 
.A(n_1722),
.Y(n_1913)
);

INVxp67_ASAP7_75t_L g1914 ( 
.A(n_1658),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1672),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1617),
.B(n_910),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1677),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1794),
.B(n_1060),
.Y(n_1918)
);

CKINVDCx11_ASAP7_75t_R g1919 ( 
.A(n_1621),
.Y(n_1919)
);

INVx3_ASAP7_75t_L g1920 ( 
.A(n_1722),
.Y(n_1920)
);

AOI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1687),
.A2(n_1063),
.B1(n_1068),
.B2(n_1062),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1727),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1636),
.B(n_963),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1676),
.A2(n_1072),
.B1(n_1076),
.B2(n_1070),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_1786),
.Y(n_1925)
);

BUFx6f_ASAP7_75t_L g1926 ( 
.A(n_1666),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1819),
.B(n_1080),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1796),
.B(n_915),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1820),
.B(n_1082),
.Y(n_1929)
);

OR2x6_ASAP7_75t_L g1930 ( 
.A(n_1650),
.B(n_892),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1680),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1657),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1691),
.B(n_1084),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1660),
.Y(n_1934)
);

BUFx3_ASAP7_75t_L g1935 ( 
.A(n_1809),
.Y(n_1935)
);

INVx6_ASAP7_75t_L g1936 ( 
.A(n_1689),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1676),
.A2(n_932),
.B1(n_937),
.B2(n_921),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_1769),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1626),
.B(n_1090),
.Y(n_1939)
);

AO22x1_ASAP7_75t_L g1940 ( 
.A1(n_1676),
.A2(n_1222),
.B1(n_941),
.B2(n_942),
.Y(n_1940)
);

AOI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1782),
.A2(n_943),
.B1(n_944),
.B2(n_939),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1821),
.B(n_1092),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1823),
.B(n_1825),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1668),
.Y(n_1944)
);

NOR2x2_ASAP7_75t_L g1945 ( 
.A(n_1843),
.B(n_967),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1673),
.Y(n_1946)
);

BUFx3_ASAP7_75t_L g1947 ( 
.A(n_1666),
.Y(n_1947)
);

BUFx2_ASAP7_75t_L g1948 ( 
.A(n_1700),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1741),
.B(n_1095),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1770),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_SL g1951 ( 
.A(n_1826),
.B(n_1097),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1828),
.B(n_1846),
.Y(n_1952)
);

INVx5_ASAP7_75t_L g1953 ( 
.A(n_1666),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1830),
.B(n_1098),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_L g1955 ( 
.A(n_1710),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1833),
.B(n_1101),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1675),
.Y(n_1957)
);

A2O1A1Ixp33_ASAP7_75t_L g1958 ( 
.A1(n_1654),
.A2(n_955),
.B(n_956),
.C(n_954),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1678),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1685),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1810),
.B(n_973),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1835),
.B(n_1104),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1688),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1837),
.B(n_1108),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1648),
.B(n_1110),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1623),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1631),
.B(n_1111),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1644),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1804),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1705),
.Y(n_1970)
);

OAI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1845),
.A2(n_979),
.B1(n_989),
.B2(n_977),
.Y(n_1971)
);

INVx2_ASAP7_75t_SL g1972 ( 
.A(n_1695),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1619),
.B(n_995),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1736),
.B(n_996),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1812),
.Y(n_1975)
);

BUFx10_ASAP7_75t_L g1976 ( 
.A(n_1759),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1816),
.B(n_961),
.Y(n_1977)
);

AOI22xp33_ASAP7_75t_L g1978 ( 
.A1(n_1782),
.A2(n_974),
.B1(n_981),
.B2(n_965),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1818),
.Y(n_1979)
);

INVx2_ASAP7_75t_SL g1980 ( 
.A(n_1689),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1710),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1832),
.Y(n_1982)
);

BUFx8_ASAP7_75t_L g1983 ( 
.A(n_1743),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1797),
.B(n_1114),
.Y(n_1984)
);

BUFx2_ASAP7_75t_L g1985 ( 
.A(n_1716),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1844),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_1710),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1739),
.A2(n_1332),
.B1(n_1011),
.B2(n_1036),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1632),
.B(n_1116),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1659),
.B(n_1119),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1702),
.Y(n_1991)
);

NAND2x1p5_ASAP7_75t_L g1992 ( 
.A(n_1714),
.B(n_984),
.Y(n_1992)
);

INVx2_ASAP7_75t_SL g1993 ( 
.A(n_1725),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1776),
.Y(n_1994)
);

A2O1A1Ixp33_ASAP7_75t_L g1995 ( 
.A1(n_1627),
.A2(n_999),
.B(n_1015),
.C(n_994),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1738),
.B(n_1009),
.Y(n_1996)
);

AND2x6_ASAP7_75t_SL g1997 ( 
.A(n_1778),
.B(n_1019),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1665),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1746),
.B(n_1050),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1643),
.B(n_1053),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1690),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1684),
.B(n_1066),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1708),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1674),
.B(n_1122),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_R g2005 ( 
.A(n_1697),
.B(n_1073),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1800),
.B(n_1124),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1679),
.Y(n_2007)
);

AOI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1724),
.A2(n_1027),
.B1(n_1038),
.B2(n_1026),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1779),
.B(n_1083),
.Y(n_2009)
);

NAND2x1p5_ASAP7_75t_L g2010 ( 
.A(n_1839),
.B(n_1042),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1709),
.B(n_1715),
.Y(n_2011)
);

NOR2xp67_ASAP7_75t_L g2012 ( 
.A(n_1747),
.B(n_24),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1744),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1791),
.B(n_1178),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1806),
.B(n_1128),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1703),
.Y(n_2016)
);

NAND2x1p5_ASAP7_75t_L g2017 ( 
.A(n_1824),
.B(n_1045),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1749),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1811),
.B(n_1131),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1701),
.Y(n_2020)
);

NOR2x2_ASAP7_75t_L g2021 ( 
.A(n_1633),
.B(n_1200),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1726),
.B(n_1046),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1664),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1704),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_1742),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_L g2026 ( 
.A(n_1618),
.B(n_1203),
.Y(n_2026)
);

INVx4_ASAP7_75t_L g2027 ( 
.A(n_1706),
.Y(n_2027)
);

AND2x4_ASAP7_75t_L g2028 ( 
.A(n_1730),
.B(n_1049),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1707),
.Y(n_2029)
);

AOI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_1629),
.A2(n_1135),
.B1(n_1136),
.B2(n_1132),
.Y(n_2030)
);

AO22x1_ASAP7_75t_L g2031 ( 
.A1(n_1670),
.A2(n_1138),
.B1(n_1141),
.B2(n_1137),
.Y(n_2031)
);

INVx2_ASAP7_75t_SL g2032 ( 
.A(n_1732),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1813),
.B(n_1142),
.Y(n_2033)
);

BUFx12f_ASAP7_75t_L g2034 ( 
.A(n_1787),
.Y(n_2034)
);

AOI22xp33_ASAP7_75t_L g2035 ( 
.A1(n_1712),
.A2(n_1056),
.B1(n_1059),
.B2(n_1052),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1815),
.B(n_1144),
.Y(n_2036)
);

OAI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_1751),
.A2(n_1226),
.B1(n_1229),
.B2(n_1205),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1713),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_L g2039 ( 
.A(n_1754),
.B(n_1230),
.Y(n_2039)
);

INVx6_ASAP7_75t_L g2040 ( 
.A(n_1787),
.Y(n_2040)
);

INVxp67_ASAP7_75t_L g2041 ( 
.A(n_1822),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1836),
.B(n_1147),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1723),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1841),
.B(n_1692),
.Y(n_2044)
);

AND2x4_ASAP7_75t_L g2045 ( 
.A(n_1733),
.B(n_1622),
.Y(n_2045)
);

BUFx6f_ASAP7_75t_L g2046 ( 
.A(n_1641),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_1671),
.Y(n_2047)
);

INVx3_ASAP7_75t_L g2048 ( 
.A(n_1693),
.Y(n_2048)
);

AND2x6_ASAP7_75t_SL g2049 ( 
.A(n_1719),
.B(n_1065),
.Y(n_2049)
);

NOR2xp33_ASAP7_75t_L g2050 ( 
.A(n_1756),
.B(n_1236),
.Y(n_2050)
);

OR2x6_ASAP7_75t_L g2051 ( 
.A(n_1774),
.B(n_892),
.Y(n_2051)
);

BUFx2_ASAP7_75t_L g2052 ( 
.A(n_1757),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1740),
.B(n_1153),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1653),
.Y(n_2054)
);

INVx2_ASAP7_75t_SL g2055 ( 
.A(n_1734),
.Y(n_2055)
);

CKINVDCx5p33_ASAP7_75t_R g2056 ( 
.A(n_1766),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_1767),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1683),
.B(n_1159),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1768),
.B(n_1160),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1721),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1661),
.Y(n_2061)
);

AND2x6_ASAP7_75t_SL g2062 ( 
.A(n_1772),
.B(n_1067),
.Y(n_2062)
);

INVx5_ASAP7_75t_L g2063 ( 
.A(n_1717),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1635),
.B(n_1166),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1711),
.B(n_1167),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_1805),
.A2(n_1078),
.B1(n_1079),
.B2(n_1074),
.Y(n_2066)
);

INVx4_ASAP7_75t_L g2067 ( 
.A(n_1720),
.Y(n_2067)
);

INVx3_ASAP7_75t_L g2068 ( 
.A(n_1745),
.Y(n_2068)
);

BUFx2_ASAP7_75t_L g2069 ( 
.A(n_1696),
.Y(n_2069)
);

AND2x6_ASAP7_75t_L g2070 ( 
.A(n_1748),
.B(n_903),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1829),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1737),
.B(n_1238),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1831),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1834),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1760),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1755),
.B(n_1169),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1838),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1785),
.Y(n_2078)
);

INVx2_ASAP7_75t_SL g2079 ( 
.A(n_1735),
.Y(n_2079)
);

OAI22xp33_ASAP7_75t_L g2080 ( 
.A1(n_1788),
.A2(n_1250),
.B1(n_1273),
.B2(n_1240),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1624),
.B(n_1173),
.Y(n_2081)
);

OR2x6_ASAP7_75t_L g2082 ( 
.A(n_1763),
.B(n_903),
.Y(n_2082)
);

AND2x6_ASAP7_75t_SL g2083 ( 
.A(n_1781),
.B(n_1085),
.Y(n_2083)
);

INVxp67_ASAP7_75t_L g2084 ( 
.A(n_1731),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1795),
.B(n_1177),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1827),
.B(n_1180),
.Y(n_2086)
);

INVx2_ASAP7_75t_SL g2087 ( 
.A(n_1777),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1790),
.Y(n_2088)
);

AND2x6_ASAP7_75t_L g2089 ( 
.A(n_1752),
.B(n_928),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1848),
.B(n_1181),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1753),
.B(n_1182),
.Y(n_2091)
);

BUFx6f_ASAP7_75t_L g2092 ( 
.A(n_1758),
.Y(n_2092)
);

BUFx3_ASAP7_75t_L g2093 ( 
.A(n_1761),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_1762),
.B(n_1183),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1780),
.B(n_1186),
.Y(n_2095)
);

INVx2_ASAP7_75t_SL g2096 ( 
.A(n_1764),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1765),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1771),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1775),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1783),
.B(n_1188),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1784),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1620),
.B(n_1189),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1628),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1630),
.B(n_1190),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_SL g2105 ( 
.A(n_1620),
.B(n_1192),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_1617),
.B(n_1086),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_L g2107 ( 
.A(n_1620),
.Y(n_2107)
);

INVx5_ASAP7_75t_L g2108 ( 
.A(n_1620),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1630),
.B(n_1195),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1620),
.B(n_1197),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1628),
.Y(n_2111)
);

AOI22xp33_ASAP7_75t_L g2112 ( 
.A1(n_1676),
.A2(n_1089),
.B1(n_1099),
.B2(n_1088),
.Y(n_2112)
);

AOI21xp5_ASAP7_75t_L g2113 ( 
.A1(n_1849),
.A2(n_1105),
.B(n_1103),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1620),
.B(n_1198),
.Y(n_2114)
);

BUFx3_ASAP7_75t_L g2115 ( 
.A(n_1840),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1628),
.Y(n_2116)
);

HB1xp67_ASAP7_75t_L g2117 ( 
.A(n_1840),
.Y(n_2117)
);

BUFx6f_ASAP7_75t_L g2118 ( 
.A(n_1620),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1630),
.B(n_1202),
.Y(n_2119)
);

OR2x6_ASAP7_75t_L g2120 ( 
.A(n_1669),
.B(n_928),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1628),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1630),
.B(n_1207),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_1676),
.A2(n_1107),
.B1(n_1109),
.B2(n_1106),
.Y(n_2123)
);

INVxp67_ASAP7_75t_SL g2124 ( 
.A(n_1620),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1628),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_1616),
.B(n_1285),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1630),
.B(n_1208),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_1849),
.A2(n_1118),
.B(n_1117),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1628),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_SL g2130 ( 
.A(n_1620),
.B(n_1209),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1628),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1628),
.Y(n_2132)
);

BUFx6f_ASAP7_75t_L g2133 ( 
.A(n_1620),
.Y(n_2133)
);

AOI22xp33_ASAP7_75t_L g2134 ( 
.A1(n_1676),
.A2(n_1127),
.B1(n_1139),
.B2(n_1121),
.Y(n_2134)
);

BUFx3_ASAP7_75t_L g2135 ( 
.A(n_1840),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1628),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1943),
.B(n_1210),
.Y(n_2137)
);

OAI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_1877),
.A2(n_1301),
.B1(n_1310),
.B2(n_1297),
.Y(n_2138)
);

AOI21xp5_ASAP7_75t_L g2139 ( 
.A1(n_1952),
.A2(n_1146),
.B(n_1145),
.Y(n_2139)
);

O2A1O1Ixp33_ASAP7_75t_L g2140 ( 
.A1(n_1958),
.A2(n_1150),
.B(n_1154),
.C(n_1149),
.Y(n_2140)
);

OAI22xp5_ASAP7_75t_SL g2141 ( 
.A1(n_2120),
.A2(n_1217),
.B1(n_1220),
.B2(n_1216),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1969),
.B(n_1227),
.Y(n_2142)
);

AOI22xp5_ASAP7_75t_L g2143 ( 
.A1(n_2126),
.A2(n_1235),
.B1(n_1241),
.B2(n_1232),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1853),
.Y(n_2144)
);

BUFx3_ASAP7_75t_L g2145 ( 
.A(n_1887),
.Y(n_2145)
);

NAND3xp33_ASAP7_75t_SL g2146 ( 
.A(n_2005),
.B(n_1243),
.C(n_1242),
.Y(n_2146)
);

A2O1A1Ixp33_ASAP7_75t_L g2147 ( 
.A1(n_2044),
.A2(n_1157),
.B(n_1158),
.C(n_1155),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1975),
.Y(n_2148)
);

A2O1A1Ixp33_ASAP7_75t_L g2149 ( 
.A1(n_2001),
.A2(n_1165),
.B(n_1168),
.C(n_1164),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1979),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1858),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_1878),
.B(n_1320),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1982),
.Y(n_2153)
);

AOI33xp33_ASAP7_75t_L g2154 ( 
.A1(n_2008),
.A2(n_1193),
.A3(n_1179),
.B1(n_1194),
.B2(n_1184),
.B3(n_1175),
.Y(n_2154)
);

BUFx3_ASAP7_75t_L g2155 ( 
.A(n_1887),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1986),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1859),
.Y(n_2157)
);

HB1xp67_ASAP7_75t_L g2158 ( 
.A(n_2120),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1864),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1874),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2103),
.Y(n_2161)
);

OR2x2_ASAP7_75t_L g2162 ( 
.A(n_1988),
.B(n_1244),
.Y(n_2162)
);

O2A1O1Ixp33_ASAP7_75t_L g2163 ( 
.A1(n_1995),
.A2(n_1214),
.B(n_1221),
.C(n_1212),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_R g2164 ( 
.A(n_1865),
.B(n_1249),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_1878),
.B(n_1251),
.Y(n_2165)
);

AND2x4_ASAP7_75t_L g2166 ( 
.A(n_2057),
.B(n_1234),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_1882),
.Y(n_2167)
);

INVx4_ASAP7_75t_L g2168 ( 
.A(n_1953),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2111),
.B(n_1252),
.Y(n_2169)
);

OR2x6_ASAP7_75t_L g2170 ( 
.A(n_1948),
.B(n_931),
.Y(n_2170)
);

O2A1O1Ixp5_ASAP7_75t_L g2171 ( 
.A1(n_1876),
.A2(n_1897),
.B(n_1918),
.C(n_1881),
.Y(n_2171)
);

OAI22xp5_ASAP7_75t_L g2172 ( 
.A1(n_2041),
.A2(n_1978),
.B1(n_1941),
.B2(n_1937),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2014),
.B(n_1254),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2116),
.Y(n_2174)
);

INVx3_ASAP7_75t_L g2175 ( 
.A(n_1953),
.Y(n_2175)
);

NAND2x1p5_ASAP7_75t_L g2176 ( 
.A(n_1861),
.B(n_1140),
.Y(n_2176)
);

AOI22xp5_ASAP7_75t_L g2177 ( 
.A1(n_1851),
.A2(n_1258),
.B1(n_1259),
.B2(n_1255),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1950),
.B(n_1333),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2121),
.B(n_1260),
.Y(n_2179)
);

NOR2xp33_ASAP7_75t_L g2180 ( 
.A(n_2039),
.B(n_1261),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_1953),
.B(n_1340),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2125),
.Y(n_2182)
);

O2A1O1Ixp33_ASAP7_75t_L g2183 ( 
.A1(n_1870),
.A2(n_1256),
.B(n_1257),
.C(n_1253),
.Y(n_2183)
);

AO22x1_ASAP7_75t_L g2184 ( 
.A1(n_1945),
.A2(n_1264),
.B1(n_1265),
.B2(n_1262),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2129),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2131),
.B(n_1266),
.Y(n_2186)
);

BUFx3_ASAP7_75t_L g2187 ( 
.A(n_2034),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2132),
.Y(n_2188)
);

A2O1A1Ixp33_ASAP7_75t_L g2189 ( 
.A1(n_1907),
.A2(n_1282),
.B(n_1284),
.C(n_1267),
.Y(n_2189)
);

OAI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_1871),
.A2(n_1270),
.B1(n_1271),
.B2(n_1269),
.Y(n_2190)
);

INVx2_ASAP7_75t_SL g2191 ( 
.A(n_1867),
.Y(n_2191)
);

BUFx2_ASAP7_75t_L g2192 ( 
.A(n_1855),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_2018),
.B(n_1321),
.Y(n_2193)
);

AOI21xp5_ASAP7_75t_L g2194 ( 
.A1(n_1880),
.A2(n_1296),
.B(n_1293),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_2045),
.B(n_2013),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2136),
.B(n_1873),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1872),
.B(n_1278),
.Y(n_2197)
);

OR2x6_ASAP7_75t_L g2198 ( 
.A(n_2115),
.B(n_945),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_R g2199 ( 
.A(n_1919),
.B(n_1283),
.Y(n_2199)
);

OAI22xp5_ASAP7_75t_SL g2200 ( 
.A1(n_1904),
.A2(n_1287),
.B1(n_1288),
.B2(n_1286),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_2112),
.A2(n_1290),
.B1(n_1291),
.B2(n_1289),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1991),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_2107),
.Y(n_2203)
);

BUFx8_ASAP7_75t_SL g2204 ( 
.A(n_2135),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1916),
.B(n_1294),
.Y(n_2205)
);

OAI21xp33_ASAP7_75t_SL g2206 ( 
.A1(n_2060),
.A2(n_1318),
.B(n_1316),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_R g2207 ( 
.A(n_1925),
.B(n_1295),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_1970),
.Y(n_2208)
);

INVx2_ASAP7_75t_SL g2209 ( 
.A(n_1935),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1916),
.B(n_1303),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1928),
.B(n_1304),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_SL g2212 ( 
.A(n_2056),
.B(n_1312),
.Y(n_2212)
);

AO32x2_ASAP7_75t_L g2213 ( 
.A1(n_1856),
.A2(n_1206),
.A3(n_1140),
.B1(n_1039),
.B2(n_1051),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_2050),
.B(n_1306),
.Y(n_2214)
);

BUFx2_ASAP7_75t_L g2215 ( 
.A(n_1904),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2003),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1928),
.B(n_1308),
.Y(n_2217)
);

BUFx6f_ASAP7_75t_L g2218 ( 
.A(n_2107),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_1955),
.B(n_1319),
.Y(n_2219)
);

A2O1A1Ixp33_ASAP7_75t_L g2220 ( 
.A1(n_2113),
.A2(n_1338),
.B(n_1018),
.C(n_1039),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1955),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_1996),
.B(n_1315),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_1955),
.B(n_1326),
.Y(n_2223)
);

NOR2xp33_ASAP7_75t_L g2224 ( 
.A(n_1999),
.B(n_1317),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1987),
.Y(n_2225)
);

NOR2x1_ASAP7_75t_L g2226 ( 
.A(n_1856),
.B(n_2027),
.Y(n_2226)
);

BUFx8_ASAP7_75t_L g2227 ( 
.A(n_1884),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1977),
.B(n_1324),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2024),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_1977),
.B(n_1327),
.Y(n_2230)
);

OA22x2_ASAP7_75t_L g2231 ( 
.A1(n_1908),
.A2(n_1336),
.B1(n_1337),
.B2(n_1335),
.Y(n_2231)
);

A2O1A1Ixp33_ASAP7_75t_L g2232 ( 
.A1(n_2128),
.A2(n_1096),
.B(n_1176),
.C(n_1093),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_1987),
.Y(n_2233)
);

INVx4_ASAP7_75t_L g2234 ( 
.A(n_2108),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2106),
.B(n_1868),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2106),
.B(n_1096),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_SL g2237 ( 
.A(n_1938),
.B(n_1206),
.Y(n_2237)
);

A2O1A1Ixp33_ASAP7_75t_L g2238 ( 
.A1(n_1932),
.A2(n_1246),
.B(n_1299),
.C(n_1298),
.Y(n_2238)
);

AOI22xp33_ASAP7_75t_L g2239 ( 
.A1(n_1900),
.A2(n_1206),
.B1(n_1299),
.B2(n_1298),
.Y(n_2239)
);

OAI22xp5_ASAP7_75t_L g2240 ( 
.A1(n_2123),
.A2(n_2134),
.B1(n_1944),
.B2(n_1946),
.Y(n_2240)
);

AO22x1_ASAP7_75t_L g2241 ( 
.A1(n_1983),
.A2(n_26),
.B1(n_27),
.B2(n_25),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1869),
.B(n_24),
.Y(n_2242)
);

NOR2xp33_ASAP7_75t_L g2243 ( 
.A(n_1961),
.B(n_25),
.Y(n_2243)
);

INVx5_ASAP7_75t_L g2244 ( 
.A(n_2107),
.Y(n_2244)
);

INVx1_ASAP7_75t_SL g2245 ( 
.A(n_1890),
.Y(n_2245)
);

AOI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2037),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_2246)
);

AOI21xp5_ASAP7_75t_L g2247 ( 
.A1(n_1934),
.A2(n_29),
.B(n_30),
.Y(n_2247)
);

A2O1A1Ixp33_ASAP7_75t_SL g2248 ( 
.A1(n_1895),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_2248)
);

BUFx3_ASAP7_75t_L g2249 ( 
.A(n_1902),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_L g2250 ( 
.A(n_2118),
.Y(n_2250)
);

CKINVDCx11_ASAP7_75t_R g2251 ( 
.A(n_2083),
.Y(n_2251)
);

CKINVDCx20_ASAP7_75t_R g2252 ( 
.A(n_2117),
.Y(n_2252)
);

OAI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_1971),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2253)
);

AND2x4_ASAP7_75t_L g2254 ( 
.A(n_2043),
.B(n_35),
.Y(n_2254)
);

AOI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_1957),
.A2(n_35),
.B(n_36),
.Y(n_2255)
);

AOI21xp5_ASAP7_75t_L g2256 ( 
.A1(n_1959),
.A2(n_36),
.B(n_37),
.Y(n_2256)
);

A2O1A1Ixp33_ASAP7_75t_L g2257 ( 
.A1(n_1960),
.A2(n_40),
.B(n_37),
.C(n_39),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_2062),
.Y(n_2258)
);

OAI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_1963),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_2259)
);

NOR3xp33_ASAP7_75t_SL g2260 ( 
.A(n_1994),
.B(n_40),
.C(n_41),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2052),
.B(n_42),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_2108),
.B(n_43),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_1983),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_2108),
.B(n_43),
.Y(n_2264)
);

A2O1A1Ixp33_ASAP7_75t_L g2265 ( 
.A1(n_2012),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_2265)
);

OAI22xp33_ASAP7_75t_L g2266 ( 
.A1(n_1908),
.A2(n_1930),
.B1(n_2080),
.B2(n_1949),
.Y(n_2266)
);

INVx3_ASAP7_75t_SL g2267 ( 
.A(n_1922),
.Y(n_2267)
);

AND2x4_ASAP7_75t_L g2268 ( 
.A(n_1913),
.B(n_45),
.Y(n_2268)
);

NOR3xp33_ASAP7_75t_SL g2269 ( 
.A(n_1866),
.B(n_1923),
.C(n_2026),
.Y(n_2269)
);

INVx3_ASAP7_75t_L g2270 ( 
.A(n_1947),
.Y(n_2270)
);

BUFx3_ASAP7_75t_L g2271 ( 
.A(n_1911),
.Y(n_2271)
);

INVx2_ASAP7_75t_SL g2272 ( 
.A(n_1930),
.Y(n_2272)
);

OAI22xp5_ASAP7_75t_L g2273 ( 
.A1(n_2027),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2273)
);

AOI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_2011),
.A2(n_46),
.B(n_47),
.Y(n_2274)
);

INVx1_ASAP7_75t_SL g2275 ( 
.A(n_1894),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_2063),
.A2(n_51),
.B1(n_48),
.B2(n_50),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_R g2277 ( 
.A(n_1912),
.B(n_50),
.Y(n_2277)
);

INVx2_ASAP7_75t_SL g2278 ( 
.A(n_1936),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1985),
.B(n_50),
.Y(n_2279)
);

AOI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_2002),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_2280)
);

AOI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_1888),
.A2(n_52),
.B(n_53),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2009),
.B(n_53),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_2000),
.B(n_54),
.Y(n_2283)
);

OAI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_2063),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_2284)
);

AOI21xp5_ASAP7_75t_L g2285 ( 
.A1(n_1885),
.A2(n_55),
.B(n_56),
.Y(n_2285)
);

NOR2xp67_ASAP7_75t_L g2286 ( 
.A(n_2063),
.B(n_55),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_2049),
.Y(n_2287)
);

INVx5_ASAP7_75t_L g2288 ( 
.A(n_2118),
.Y(n_2288)
);

NOR3xp33_ASAP7_75t_SL g2289 ( 
.A(n_1973),
.B(n_57),
.C(n_58),
.Y(n_2289)
);

BUFx2_ASAP7_75t_L g2290 ( 
.A(n_1893),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2022),
.B(n_2028),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2029),
.Y(n_2292)
);

BUFx6f_ASAP7_75t_L g2293 ( 
.A(n_2133),
.Y(n_2293)
);

O2A1O1Ixp33_ASAP7_75t_L g2294 ( 
.A1(n_1967),
.A2(n_1862),
.B(n_1863),
.C(n_1850),
.Y(n_2294)
);

CKINVDCx20_ASAP7_75t_R g2295 ( 
.A(n_1914),
.Y(n_2295)
);

OAI22x1_ASAP7_75t_L g2296 ( 
.A1(n_2017),
.A2(n_2021),
.B1(n_1924),
.B2(n_2022),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2038),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1903),
.Y(n_2298)
);

O2A1O1Ixp33_ASAP7_75t_L g2299 ( 
.A1(n_2104),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_2299)
);

BUFx2_ASAP7_75t_L g2300 ( 
.A(n_2070),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2028),
.B(n_1972),
.Y(n_2301)
);

OAI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_2067),
.A2(n_60),
.B1(n_57),
.B2(n_59),
.Y(n_2302)
);

INVx3_ASAP7_75t_L g2303 ( 
.A(n_2040),
.Y(n_2303)
);

NAND2x1p5_ASAP7_75t_L g2304 ( 
.A(n_1898),
.B(n_59),
.Y(n_2304)
);

OAI22xp5_ASAP7_75t_L g2305 ( 
.A1(n_2067),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_SL g2306 ( 
.A(n_1854),
.B(n_62),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2109),
.B(n_61),
.Y(n_2307)
);

NOR2xp33_ASAP7_75t_L g2308 ( 
.A(n_1936),
.B(n_61),
.Y(n_2308)
);

AOI21xp5_ASAP7_75t_L g2309 ( 
.A1(n_1965),
.A2(n_63),
.B(n_65),
.Y(n_2309)
);

BUFx3_ASAP7_75t_L g2310 ( 
.A(n_1920),
.Y(n_2310)
);

INVx3_ASAP7_75t_L g2311 ( 
.A(n_2040),
.Y(n_2311)
);

NOR2x1_ASAP7_75t_SL g2312 ( 
.A(n_2051),
.B(n_66),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_2133),
.B(n_66),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_1921),
.B(n_65),
.Y(n_2314)
);

BUFx6f_ASAP7_75t_L g2315 ( 
.A(n_2133),
.Y(n_2315)
);

A2O1A1Ixp33_ASAP7_75t_L g2316 ( 
.A1(n_2016),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_2316)
);

BUFx3_ASAP7_75t_L g2317 ( 
.A(n_1909),
.Y(n_2317)
);

AND2x4_ASAP7_75t_L g2318 ( 
.A(n_1906),
.B(n_67),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2119),
.B(n_67),
.Y(n_2319)
);

OAI22xp5_ASAP7_75t_L g2320 ( 
.A1(n_2122),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_1910),
.Y(n_2321)
);

OAI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2127),
.A2(n_71),
.B1(n_68),
.B2(n_70),
.Y(n_2322)
);

AOI21xp5_ASAP7_75t_L g2323 ( 
.A1(n_2042),
.A2(n_68),
.B(n_70),
.Y(n_2323)
);

OAI22xp5_ASAP7_75t_L g2324 ( 
.A1(n_2097),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_1980),
.B(n_71),
.Y(n_2325)
);

NOR2xp67_ASAP7_75t_SL g2326 ( 
.A(n_2025),
.B(n_72),
.Y(n_2326)
);

A2O1A1Ixp33_ASAP7_75t_SL g2327 ( 
.A1(n_2072),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_2327)
);

BUFx3_ASAP7_75t_L g2328 ( 
.A(n_1992),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_1915),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1917),
.Y(n_2330)
);

INVxp67_ASAP7_75t_L g2331 ( 
.A(n_2051),
.Y(n_2331)
);

AOI21xp5_ASAP7_75t_L g2332 ( 
.A1(n_2006),
.A2(n_73),
.B(n_74),
.Y(n_2332)
);

NOR2xp33_ASAP7_75t_L g2333 ( 
.A(n_1933),
.B(n_74),
.Y(n_2333)
);

NOR3xp33_ASAP7_75t_SL g2334 ( 
.A(n_1939),
.B(n_75),
.C(n_76),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1886),
.B(n_75),
.Y(n_2335)
);

A2O1A1Ixp33_ASAP7_75t_L g2336 ( 
.A1(n_1931),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_2336)
);

AOI21xp5_ASAP7_75t_SL g2337 ( 
.A1(n_2124),
.A2(n_85),
.B(n_77),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2007),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_1998),
.Y(n_2339)
);

INVx3_ASAP7_75t_SL g2340 ( 
.A(n_1883),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2015),
.A2(n_77),
.B(n_78),
.Y(n_2341)
);

HB1xp67_ASAP7_75t_L g2342 ( 
.A(n_1981),
.Y(n_2342)
);

AOI21xp5_ASAP7_75t_L g2343 ( 
.A1(n_2019),
.A2(n_78),
.B(n_79),
.Y(n_2343)
);

INVx3_ASAP7_75t_L g2344 ( 
.A(n_2047),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_1891),
.B(n_79),
.Y(n_2345)
);

OR2x6_ASAP7_75t_L g2346 ( 
.A(n_1883),
.B(n_79),
.Y(n_2346)
);

AOI22xp33_ASAP7_75t_L g2347 ( 
.A1(n_1892),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_2347)
);

AOI221xp5_ASAP7_75t_L g2348 ( 
.A1(n_2031),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.C(n_83),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_1896),
.B(n_82),
.Y(n_2349)
);

HB1xp67_ASAP7_75t_L g2350 ( 
.A(n_2010),
.Y(n_2350)
);

AOI21xp5_ASAP7_75t_L g2351 ( 
.A1(n_2033),
.A2(n_83),
.B(n_84),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_1899),
.B(n_83),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_1901),
.B(n_84),
.Y(n_2353)
);

OAI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2036),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_2354)
);

A2O1A1Ixp33_ASAP7_75t_L g2355 ( 
.A1(n_1905),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_1927),
.B(n_86),
.Y(n_2356)
);

OA22x2_ASAP7_75t_L g2357 ( 
.A1(n_2030),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_1976),
.B(n_89),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2020),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_1929),
.B(n_88),
.Y(n_2360)
);

BUFx4_ASAP7_75t_SL g2361 ( 
.A(n_1997),
.Y(n_2361)
);

AOI21xp5_ASAP7_75t_L g2362 ( 
.A1(n_1956),
.A2(n_1962),
.B(n_2053),
.Y(n_2362)
);

AOI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_1942),
.A2(n_89),
.B(n_90),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_1976),
.B(n_90),
.Y(n_2364)
);

OR2x6_ASAP7_75t_L g2365 ( 
.A(n_1940),
.B(n_90),
.Y(n_2365)
);

HB1xp67_ASAP7_75t_L g2366 ( 
.A(n_2070),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2035),
.B(n_91),
.Y(n_2367)
);

AOI22xp5_ASAP7_75t_L g2368 ( 
.A1(n_1989),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_2368)
);

AOI22xp5_ASAP7_75t_L g2369 ( 
.A1(n_1951),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_2047),
.B(n_94),
.Y(n_2370)
);

AOI21xp5_ASAP7_75t_L g2371 ( 
.A1(n_1954),
.A2(n_93),
.B(n_94),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2069),
.B(n_95),
.Y(n_2372)
);

HB1xp67_ASAP7_75t_L g2373 ( 
.A(n_2070),
.Y(n_2373)
);

NOR2xp33_ASAP7_75t_L g2374 ( 
.A(n_1964),
.B(n_94),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2100),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_1940),
.B(n_96),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_1966),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_R g2378 ( 
.A(n_1860),
.B(n_858),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_2046),
.Y(n_2379)
);

NOR2xp67_ASAP7_75t_L g2380 ( 
.A(n_2048),
.B(n_102),
.Y(n_2380)
);

INVx2_ASAP7_75t_SL g2381 ( 
.A(n_1852),
.Y(n_2381)
);

OR2x6_ASAP7_75t_L g2382 ( 
.A(n_2079),
.B(n_104),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2059),
.B(n_105),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_1990),
.B(n_106),
.Y(n_2384)
);

AND2x2_ASAP7_75t_SL g2385 ( 
.A(n_2070),
.B(n_106),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_SL g2386 ( 
.A(n_2064),
.B(n_107),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_1984),
.B(n_107),
.Y(n_2387)
);

BUFx2_ASAP7_75t_SL g2388 ( 
.A(n_2089),
.Y(n_2388)
);

OAI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_2078),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_2389)
);

OR2x2_ASAP7_75t_L g2390 ( 
.A(n_2076),
.B(n_108),
.Y(n_2390)
);

BUFx2_ASAP7_75t_L g2391 ( 
.A(n_2089),
.Y(n_2391)
);

AOI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_2075),
.A2(n_109),
.B(n_111),
.Y(n_2392)
);

OAI22xp5_ASAP7_75t_L g2393 ( 
.A1(n_1993),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1968),
.Y(n_2394)
);

A2O1A1Ixp33_ASAP7_75t_L g2395 ( 
.A1(n_2071),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_2395)
);

OR2x6_ASAP7_75t_L g2396 ( 
.A(n_1879),
.B(n_115),
.Y(n_2396)
);

AOI22xp5_ASAP7_75t_L g2397 ( 
.A1(n_2004),
.A2(n_120),
.B1(n_116),
.B2(n_117),
.Y(n_2397)
);

AND2x4_ASAP7_75t_L g2398 ( 
.A(n_1857),
.B(n_121),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_SL g2399 ( 
.A(n_2081),
.B(n_123),
.Y(n_2399)
);

BUFx3_ASAP7_75t_L g2400 ( 
.A(n_2089),
.Y(n_2400)
);

AND2x2_ASAP7_75t_SL g2401 ( 
.A(n_2023),
.B(n_123),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2073),
.Y(n_2402)
);

AND2x4_ASAP7_75t_L g2403 ( 
.A(n_1875),
.B(n_124),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2058),
.B(n_125),
.Y(n_2404)
);

CKINVDCx20_ASAP7_75t_R g2405 ( 
.A(n_2102),
.Y(n_2405)
);

CKINVDCx8_ASAP7_75t_R g2406 ( 
.A(n_1889),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_2066),
.B(n_126),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_2065),
.B(n_862),
.Y(n_2408)
);

BUFx12f_ASAP7_75t_L g2409 ( 
.A(n_2032),
.Y(n_2409)
);

OAI22xp5_ASAP7_75t_SL g2410 ( 
.A1(n_2055),
.A2(n_131),
.B1(n_127),
.B2(n_128),
.Y(n_2410)
);

AOI21xp5_ASAP7_75t_L g2411 ( 
.A1(n_2088),
.A2(n_132),
.B(n_133),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2074),
.B(n_2077),
.Y(n_2412)
);

NAND2x1p5_ASAP7_75t_L g2413 ( 
.A(n_2105),
.B(n_133),
.Y(n_2413)
);

AOI21xp5_ASAP7_75t_L g2414 ( 
.A1(n_2098),
.A2(n_132),
.B(n_134),
.Y(n_2414)
);

AOI21xp5_ASAP7_75t_L g2415 ( 
.A1(n_2099),
.A2(n_135),
.B(n_136),
.Y(n_2415)
);

NOR2xp33_ASAP7_75t_L g2416 ( 
.A(n_2110),
.B(n_857),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2114),
.B(n_136),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2130),
.B(n_137),
.Y(n_2418)
);

NAND2x1p5_ASAP7_75t_L g2419 ( 
.A(n_2068),
.B(n_138),
.Y(n_2419)
);

BUFx2_ASAP7_75t_L g2420 ( 
.A(n_2089),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_2095),
.B(n_2085),
.Y(n_2421)
);

INVxp67_ASAP7_75t_SL g2422 ( 
.A(n_2087),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_SL g2423 ( 
.A(n_2084),
.B(n_137),
.Y(n_2423)
);

OAI21x1_ASAP7_75t_L g2424 ( 
.A1(n_2101),
.A2(n_138),
.B(n_139),
.Y(n_2424)
);

NOR2xp33_ASAP7_75t_L g2425 ( 
.A(n_2091),
.B(n_2094),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_SL g2426 ( 
.A(n_2086),
.B(n_140),
.Y(n_2426)
);

A2O1A1Ixp33_ASAP7_75t_L g2427 ( 
.A1(n_2054),
.A2(n_144),
.B(n_141),
.C(n_142),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2090),
.B(n_142),
.Y(n_2428)
);

NAND3xp33_ASAP7_75t_SL g2429 ( 
.A(n_2061),
.B(n_863),
.C(n_144),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2082),
.Y(n_2430)
);

BUFx2_ASAP7_75t_L g2431 ( 
.A(n_2082),
.Y(n_2431)
);

BUFx6f_ASAP7_75t_L g2432 ( 
.A(n_2046),
.Y(n_2432)
);

OA22x2_ASAP7_75t_L g2433 ( 
.A1(n_2096),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_2433)
);

OAI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2093),
.A2(n_151),
.B1(n_148),
.B2(n_150),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_2092),
.Y(n_2435)
);

OAI22xp5_ASAP7_75t_SL g2436 ( 
.A1(n_2092),
.A2(n_152),
.B1(n_148),
.B2(n_151),
.Y(n_2436)
);

NOR2xp33_ASAP7_75t_L g2437 ( 
.A(n_2039),
.B(n_855),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1969),
.Y(n_2438)
);

NOR2xp67_ASAP7_75t_SL g2439 ( 
.A(n_1878),
.B(n_152),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_1969),
.Y(n_2440)
);

BUFx4f_ASAP7_75t_L g2441 ( 
.A(n_1867),
.Y(n_2441)
);

NAND2x1p5_ASAP7_75t_L g2442 ( 
.A(n_1878),
.B(n_154),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_1943),
.B(n_153),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_1943),
.B(n_154),
.Y(n_2444)
);

AOI21xp5_ASAP7_75t_L g2445 ( 
.A1(n_1943),
.A2(n_155),
.B(n_156),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2014),
.B(n_156),
.Y(n_2446)
);

INVxp67_ASAP7_75t_L g2447 ( 
.A(n_2120),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_1919),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_1943),
.B(n_158),
.Y(n_2449)
);

BUFx2_ASAP7_75t_L g2450 ( 
.A(n_2120),
.Y(n_2450)
);

INVx2_ASAP7_75t_SL g2451 ( 
.A(n_1861),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_1853),
.Y(n_2452)
);

NOR3xp33_ASAP7_75t_L g2453 ( 
.A(n_2031),
.B(n_159),
.C(n_160),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_1943),
.B(n_159),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_1969),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_1943),
.B(n_162),
.Y(n_2456)
);

INVx5_ASAP7_75t_L g2457 ( 
.A(n_2120),
.Y(n_2457)
);

INVx2_ASAP7_75t_SL g2458 ( 
.A(n_1861),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_1853),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_1969),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_1943),
.B(n_163),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_SL g2462 ( 
.A(n_1878),
.B(n_164),
.Y(n_2462)
);

INVx5_ASAP7_75t_L g2463 ( 
.A(n_2120),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_1943),
.B(n_165),
.Y(n_2464)
);

AO21x1_ASAP7_75t_L g2465 ( 
.A1(n_2044),
.A2(n_166),
.B(n_167),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_1853),
.Y(n_2466)
);

BUFx6f_ASAP7_75t_L g2467 ( 
.A(n_2107),
.Y(n_2467)
);

BUFx6f_ASAP7_75t_L g2468 ( 
.A(n_2107),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_1943),
.B(n_168),
.Y(n_2469)
);

O2A1O1Ixp33_ASAP7_75t_L g2470 ( 
.A1(n_1958),
.A2(n_170),
.B(n_168),
.C(n_169),
.Y(n_2470)
);

AOI21xp5_ASAP7_75t_L g2471 ( 
.A1(n_1943),
.A2(n_169),
.B(n_170),
.Y(n_2471)
);

NOR2xp33_ASAP7_75t_R g2472 ( 
.A(n_1865),
.B(n_861),
.Y(n_2472)
);

O2A1O1Ixp5_ASAP7_75t_L g2473 ( 
.A1(n_1876),
.A2(n_174),
.B(n_172),
.C(n_173),
.Y(n_2473)
);

BUFx2_ASAP7_75t_L g2474 ( 
.A(n_2120),
.Y(n_2474)
);

BUFx6f_ASAP7_75t_L g2475 ( 
.A(n_2107),
.Y(n_2475)
);

AOI21x1_ASAP7_75t_L g2476 ( 
.A1(n_1940),
.A2(n_174),
.B(n_175),
.Y(n_2476)
);

AOI22xp33_ASAP7_75t_L g2477 ( 
.A1(n_1974),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_R g2478 ( 
.A(n_1865),
.B(n_853),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_1969),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_1943),
.B(n_178),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_1969),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_1943),
.B(n_180),
.Y(n_2482)
);

BUFx6f_ASAP7_75t_L g2483 ( 
.A(n_2107),
.Y(n_2483)
);

OAI21xp33_ASAP7_75t_SL g2484 ( 
.A1(n_1877),
.A2(n_180),
.B(n_181),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_1943),
.B(n_181),
.Y(n_2485)
);

INVx4_ASAP7_75t_L g2486 ( 
.A(n_1953),
.Y(n_2486)
);

INVx1_ASAP7_75t_SL g2487 ( 
.A(n_1867),
.Y(n_2487)
);

OAI22xp5_ASAP7_75t_L g2488 ( 
.A1(n_1877),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_2488)
);

INVx3_ASAP7_75t_L g2489 ( 
.A(n_1953),
.Y(n_2489)
);

HB1xp67_ASAP7_75t_L g2490 ( 
.A(n_2120),
.Y(n_2490)
);

BUFx6f_ASAP7_75t_L g2491 ( 
.A(n_2107),
.Y(n_2491)
);

OA22x2_ASAP7_75t_L g2492 ( 
.A1(n_1867),
.A2(n_192),
.B1(n_187),
.B2(n_189),
.Y(n_2492)
);

HB1xp67_ASAP7_75t_L g2493 ( 
.A(n_2120),
.Y(n_2493)
);

A2O1A1Ixp33_ASAP7_75t_L g2494 ( 
.A1(n_1943),
.A2(n_193),
.B(n_189),
.C(n_192),
.Y(n_2494)
);

INVx2_ASAP7_75t_SL g2495 ( 
.A(n_1861),
.Y(n_2495)
);

BUFx12f_ASAP7_75t_L g2496 ( 
.A(n_1919),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_1943),
.B(n_194),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_1943),
.B(n_194),
.Y(n_2498)
);

INVx4_ASAP7_75t_L g2499 ( 
.A(n_1953),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_1943),
.B(n_195),
.Y(n_2500)
);

BUFx3_ASAP7_75t_L g2501 ( 
.A(n_1887),
.Y(n_2501)
);

NOR2xp33_ASAP7_75t_L g2502 ( 
.A(n_2039),
.B(n_851),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_1943),
.B(n_196),
.Y(n_2503)
);

OAI22xp5_ASAP7_75t_L g2504 ( 
.A1(n_1877),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_2504)
);

OAI22xp5_ASAP7_75t_L g2505 ( 
.A1(n_1877),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_2505)
);

AOI22xp33_ASAP7_75t_L g2506 ( 
.A1(n_1974),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_SL g2507 ( 
.A(n_1878),
.B(n_201),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_1943),
.B(n_202),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_SL g2509 ( 
.A(n_1878),
.B(n_203),
.Y(n_2509)
);

BUFx3_ASAP7_75t_L g2510 ( 
.A(n_1887),
.Y(n_2510)
);

INVx5_ASAP7_75t_L g2511 ( 
.A(n_2120),
.Y(n_2511)
);

NOR2xp33_ASAP7_75t_L g2512 ( 
.A(n_2039),
.B(n_857),
.Y(n_2512)
);

INVx4_ASAP7_75t_L g2513 ( 
.A(n_1953),
.Y(n_2513)
);

CKINVDCx5p33_ASAP7_75t_R g2514 ( 
.A(n_1919),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_SL g2515 ( 
.A(n_1878),
.B(n_205),
.Y(n_2515)
);

INVx4_ASAP7_75t_L g2516 ( 
.A(n_1953),
.Y(n_2516)
);

O2A1O1Ixp33_ASAP7_75t_L g2517 ( 
.A1(n_1958),
.A2(n_209),
.B(n_207),
.C(n_208),
.Y(n_2517)
);

OAI22xp5_ASAP7_75t_L g2518 ( 
.A1(n_1877),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_2518)
);

OAI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_1877),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_1853),
.Y(n_2520)
);

OAI22xp5_ASAP7_75t_L g2521 ( 
.A1(n_1877),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_2521)
);

BUFx3_ASAP7_75t_L g2522 ( 
.A(n_1887),
.Y(n_2522)
);

AOI22xp5_ASAP7_75t_SL g2523 ( 
.A1(n_1945),
.A2(n_218),
.B1(n_215),
.B2(n_217),
.Y(n_2523)
);

OR2x2_ASAP7_75t_L g2524 ( 
.A(n_1988),
.B(n_217),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_1943),
.B(n_219),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_1878),
.B(n_221),
.Y(n_2526)
);

OAI22xp5_ASAP7_75t_L g2527 ( 
.A1(n_1877),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_1969),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_L g2529 ( 
.A(n_2039),
.B(n_850),
.Y(n_2529)
);

AOI21xp5_ASAP7_75t_L g2530 ( 
.A1(n_1943),
.A2(n_225),
.B(n_226),
.Y(n_2530)
);

INVx4_ASAP7_75t_L g2531 ( 
.A(n_1953),
.Y(n_2531)
);

OR2x6_ASAP7_75t_L g2532 ( 
.A(n_1878),
.B(n_225),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_1943),
.B(n_226),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_1943),
.B(n_227),
.Y(n_2534)
);

A2O1A1Ixp33_ASAP7_75t_L g2535 ( 
.A1(n_1943),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_2535)
);

OR2x2_ASAP7_75t_L g2536 ( 
.A(n_1988),
.B(n_230),
.Y(n_2536)
);

A2O1A1Ixp33_ASAP7_75t_L g2537 ( 
.A1(n_1943),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_2537)
);

HB1xp67_ASAP7_75t_L g2538 ( 
.A(n_2120),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_1853),
.Y(n_2539)
);

OAI22xp5_ASAP7_75t_L g2540 ( 
.A1(n_1877),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_2540)
);

AOI21xp5_ASAP7_75t_L g2541 ( 
.A1(n_1943),
.A2(n_234),
.B(n_235),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_1853),
.Y(n_2542)
);

NOR2xp33_ASAP7_75t_L g2543 ( 
.A(n_2039),
.B(n_862),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_1943),
.B(n_236),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_SL g2545 ( 
.A(n_1878),
.B(n_238),
.Y(n_2545)
);

A2O1A1Ixp33_ASAP7_75t_L g2546 ( 
.A1(n_1943),
.A2(n_241),
.B(n_239),
.C(n_240),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_1943),
.B(n_242),
.Y(n_2547)
);

AOI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_1943),
.A2(n_243),
.B(n_244),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_1853),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_1953),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_SL g2551 ( 
.A(n_1878),
.B(n_243),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_1853),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_1969),
.Y(n_2553)
);

NOR2xp33_ASAP7_75t_L g2554 ( 
.A(n_2039),
.B(n_851),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_1943),
.B(n_244),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_SL g2556 ( 
.A(n_1878),
.B(n_245),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_1943),
.B(n_245),
.Y(n_2557)
);

OAI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_1877),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_2558)
);

AOI22xp5_ASAP7_75t_L g2559 ( 
.A1(n_2126),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_2559)
);

AND2x4_ASAP7_75t_L g2560 ( 
.A(n_2057),
.B(n_250),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_SL g2561 ( 
.A(n_1878),
.B(n_251),
.Y(n_2561)
);

INVx3_ASAP7_75t_L g2562 ( 
.A(n_1953),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_SL g2563 ( 
.A(n_1878),
.B(n_251),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_1969),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_1853),
.Y(n_2565)
);

AND2x4_ASAP7_75t_L g2566 ( 
.A(n_2057),
.B(n_252),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_SL g2567 ( 
.A(n_1878),
.B(n_252),
.Y(n_2567)
);

OAI22xp5_ASAP7_75t_L g2568 ( 
.A1(n_1877),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_2568)
);

A2O1A1Ixp33_ASAP7_75t_L g2569 ( 
.A1(n_1943),
.A2(n_256),
.B(n_254),
.C(n_255),
.Y(n_2569)
);

AOI21xp5_ASAP7_75t_L g2570 ( 
.A1(n_1943),
.A2(n_256),
.B(n_257),
.Y(n_2570)
);

NOR2xp33_ASAP7_75t_L g2571 ( 
.A(n_2039),
.B(n_850),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_1919),
.Y(n_2572)
);

OAI22xp5_ASAP7_75t_L g2573 ( 
.A1(n_1877),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_2573)
);

OR2x6_ASAP7_75t_L g2574 ( 
.A(n_1878),
.B(n_259),
.Y(n_2574)
);

O2A1O1Ixp33_ASAP7_75t_SL g2575 ( 
.A1(n_1876),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_2575)
);

AOI21xp5_ASAP7_75t_L g2576 ( 
.A1(n_1943),
.A2(n_261),
.B(n_262),
.Y(n_2576)
);

NOR3xp33_ASAP7_75t_SL g2577 ( 
.A(n_1925),
.B(n_264),
.C(n_267),
.Y(n_2577)
);

AOI21xp5_ASAP7_75t_L g2578 ( 
.A1(n_1943),
.A2(n_264),
.B(n_268),
.Y(n_2578)
);

AOI21xp5_ASAP7_75t_L g2579 ( 
.A1(n_1943),
.A2(n_268),
.B(n_269),
.Y(n_2579)
);

OAI21xp33_ASAP7_75t_L g2580 ( 
.A1(n_1943),
.A2(n_269),
.B(n_270),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_1969),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_1853),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_1943),
.B(n_270),
.Y(n_2583)
);

O2A1O1Ixp33_ASAP7_75t_L g2584 ( 
.A1(n_1958),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_1943),
.B(n_271),
.Y(n_2585)
);

CKINVDCx20_ASAP7_75t_R g2586 ( 
.A(n_1919),
.Y(n_2586)
);

AOI221xp5_ASAP7_75t_L g2587 ( 
.A1(n_1916),
.A2(n_275),
.B1(n_272),
.B2(n_274),
.C(n_276),
.Y(n_2587)
);

AOI21x1_ASAP7_75t_L g2588 ( 
.A1(n_1940),
.A2(n_274),
.B(n_276),
.Y(n_2588)
);

NOR3xp33_ASAP7_75t_SL g2589 ( 
.A(n_1925),
.B(n_277),
.C(n_278),
.Y(n_2589)
);

A2O1A1Ixp33_ASAP7_75t_L g2590 ( 
.A1(n_1943),
.A2(n_281),
.B(n_277),
.C(n_280),
.Y(n_2590)
);

BUFx4f_ASAP7_75t_L g2591 ( 
.A(n_1867),
.Y(n_2591)
);

NOR2xp33_ASAP7_75t_L g2592 ( 
.A(n_2039),
.B(n_860),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_SL g2593 ( 
.A(n_1878),
.B(n_282),
.Y(n_2593)
);

INVx3_ASAP7_75t_SL g2594 ( 
.A(n_1945),
.Y(n_2594)
);

A2O1A1Ixp33_ASAP7_75t_L g2595 ( 
.A1(n_1943),
.A2(n_286),
.B(n_284),
.C(n_285),
.Y(n_2595)
);

AND2x2_ASAP7_75t_L g2596 ( 
.A(n_2014),
.B(n_286),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_1943),
.B(n_287),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_1853),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_1853),
.Y(n_2599)
);

AND2x6_ASAP7_75t_L g2600 ( 
.A(n_1926),
.B(n_289),
.Y(n_2600)
);

OAI21xp33_ASAP7_75t_SL g2601 ( 
.A1(n_1877),
.A2(n_291),
.B(n_292),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_1943),
.B(n_291),
.Y(n_2602)
);

NOR2xp33_ASAP7_75t_L g2603 ( 
.A(n_2039),
.B(n_849),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_1943),
.B(n_294),
.Y(n_2604)
);

INVx2_ASAP7_75t_SL g2605 ( 
.A(n_1861),
.Y(n_2605)
);

O2A1O1Ixp33_ASAP7_75t_L g2606 ( 
.A1(n_1958),
.A2(n_299),
.B(n_296),
.C(n_297),
.Y(n_2606)
);

NOR2xp67_ASAP7_75t_SL g2607 ( 
.A(n_1878),
.B(n_299),
.Y(n_2607)
);

INVx1_ASAP7_75t_SL g2608 ( 
.A(n_1867),
.Y(n_2608)
);

BUFx6f_ASAP7_75t_L g2609 ( 
.A(n_2107),
.Y(n_2609)
);

BUFx12f_ASAP7_75t_L g2610 ( 
.A(n_1919),
.Y(n_2610)
);

NOR2xp67_ASAP7_75t_L g2611 ( 
.A(n_2108),
.B(n_300),
.Y(n_2611)
);

NOR2xp33_ASAP7_75t_SL g2612 ( 
.A(n_1878),
.B(n_301),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_1853),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_1853),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_1943),
.B(n_301),
.Y(n_2615)
);

A2O1A1Ixp33_ASAP7_75t_L g2616 ( 
.A1(n_1943),
.A2(n_304),
.B(n_302),
.C(n_303),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_1853),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_1943),
.B(n_302),
.Y(n_2618)
);

OAI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_1877),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_2619)
);

AOI21xp5_ASAP7_75t_L g2620 ( 
.A1(n_1943),
.A2(n_306),
.B(n_307),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_R g2621 ( 
.A(n_1865),
.B(n_848),
.Y(n_2621)
);

NOR3xp33_ASAP7_75t_SL g2622 ( 
.A(n_1925),
.B(n_308),
.C(n_311),
.Y(n_2622)
);

BUFx2_ASAP7_75t_L g2623 ( 
.A(n_2120),
.Y(n_2623)
);

INVx3_ASAP7_75t_SL g2624 ( 
.A(n_1945),
.Y(n_2624)
);

AOI21xp5_ASAP7_75t_L g2625 ( 
.A1(n_1943),
.A2(n_311),
.B(n_312),
.Y(n_2625)
);

INVx1_ASAP7_75t_SL g2626 ( 
.A(n_1867),
.Y(n_2626)
);

NOR3xp33_ASAP7_75t_SL g2627 ( 
.A(n_1925),
.B(n_312),
.C(n_314),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_1853),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_1853),
.Y(n_2629)
);

OAI22xp5_ASAP7_75t_L g2630 ( 
.A1(n_1877),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_2630)
);

INVx2_ASAP7_75t_SL g2631 ( 
.A(n_1861),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_1969),
.Y(n_2632)
);

BUFx2_ASAP7_75t_L g2633 ( 
.A(n_2120),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_L g2634 ( 
.A(n_2039),
.B(n_852),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_L g2635 ( 
.A(n_2039),
.B(n_852),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2144),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2151),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2157),
.Y(n_2638)
);

BUFx12f_ASAP7_75t_L g2639 ( 
.A(n_2263),
.Y(n_2639)
);

BUFx6f_ASAP7_75t_L g2640 ( 
.A(n_2203),
.Y(n_2640)
);

INVx1_ASAP7_75t_SL g2641 ( 
.A(n_2290),
.Y(n_2641)
);

AO21x2_ASAP7_75t_L g2642 ( 
.A1(n_2465),
.A2(n_317),
.B(n_318),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2148),
.Y(n_2643)
);

INVx1_ASAP7_75t_SL g2644 ( 
.A(n_2167),
.Y(n_2644)
);

BUFx12f_ASAP7_75t_L g2645 ( 
.A(n_2496),
.Y(n_2645)
);

BUFx6f_ASAP7_75t_L g2646 ( 
.A(n_2203),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2173),
.B(n_2446),
.Y(n_2647)
);

OR2x2_ASAP7_75t_L g2648 ( 
.A(n_2138),
.B(n_317),
.Y(n_2648)
);

OA21x2_ASAP7_75t_L g2649 ( 
.A1(n_2424),
.A2(n_319),
.B(n_320),
.Y(n_2649)
);

INVx3_ASAP7_75t_L g2650 ( 
.A(n_2168),
.Y(n_2650)
);

OAI21xp5_ASAP7_75t_L g2651 ( 
.A1(n_2362),
.A2(n_320),
.B(n_321),
.Y(n_2651)
);

INVxp67_ASAP7_75t_SL g2652 ( 
.A(n_2254),
.Y(n_2652)
);

NAND2x1p5_ASAP7_75t_L g2653 ( 
.A(n_2168),
.B(n_321),
.Y(n_2653)
);

HB1xp67_ASAP7_75t_L g2654 ( 
.A(n_2254),
.Y(n_2654)
);

BUFx4f_ASAP7_75t_L g2655 ( 
.A(n_2624),
.Y(n_2655)
);

CKINVDCx14_ASAP7_75t_R g2656 ( 
.A(n_2441),
.Y(n_2656)
);

AOI22xp33_ASAP7_75t_L g2657 ( 
.A1(n_2594),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_2657)
);

INVx2_ASAP7_75t_SL g2658 ( 
.A(n_2441),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2150),
.Y(n_2659)
);

INVx2_ASAP7_75t_SL g2660 ( 
.A(n_2591),
.Y(n_2660)
);

BUFx6f_ASAP7_75t_L g2661 ( 
.A(n_2203),
.Y(n_2661)
);

BUFx6f_ASAP7_75t_L g2662 ( 
.A(n_2218),
.Y(n_2662)
);

AO21x2_ASAP7_75t_L g2663 ( 
.A1(n_2380),
.A2(n_323),
.B(n_325),
.Y(n_2663)
);

INVx3_ASAP7_75t_L g2664 ( 
.A(n_2486),
.Y(n_2664)
);

AOI22x1_ASAP7_75t_L g2665 ( 
.A1(n_2332),
.A2(n_329),
.B1(n_326),
.B2(n_327),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2153),
.Y(n_2666)
);

INVx1_ASAP7_75t_SL g2667 ( 
.A(n_2560),
.Y(n_2667)
);

BUFx3_ASAP7_75t_L g2668 ( 
.A(n_2187),
.Y(n_2668)
);

AO21x2_ASAP7_75t_L g2669 ( 
.A1(n_2380),
.A2(n_330),
.B(n_331),
.Y(n_2669)
);

BUFx2_ASAP7_75t_R g2670 ( 
.A(n_2145),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2174),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2156),
.Y(n_2672)
);

BUFx6f_ASAP7_75t_L g2673 ( 
.A(n_2218),
.Y(n_2673)
);

INVx1_ASAP7_75t_SL g2674 ( 
.A(n_2560),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2185),
.Y(n_2675)
);

INVx3_ASAP7_75t_L g2676 ( 
.A(n_2486),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2452),
.Y(n_2677)
);

AOI22x1_ASAP7_75t_L g2678 ( 
.A1(n_2341),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_2678)
);

HB1xp67_ASAP7_75t_L g2679 ( 
.A(n_2318),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2459),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2438),
.Y(n_2681)
);

INVx2_ASAP7_75t_SL g2682 ( 
.A(n_2591),
.Y(n_2682)
);

AND2x4_ASAP7_75t_L g2683 ( 
.A(n_2195),
.B(n_333),
.Y(n_2683)
);

OA21x2_ASAP7_75t_L g2684 ( 
.A1(n_2580),
.A2(n_335),
.B(n_336),
.Y(n_2684)
);

OAI21x1_ASAP7_75t_L g2685 ( 
.A1(n_2221),
.A2(n_2233),
.B(n_2225),
.Y(n_2685)
);

BUFx12f_ASAP7_75t_L g2686 ( 
.A(n_2610),
.Y(n_2686)
);

BUFx2_ASAP7_75t_L g2687 ( 
.A(n_2227),
.Y(n_2687)
);

OAI21x1_ASAP7_75t_L g2688 ( 
.A1(n_2171),
.A2(n_337),
.B(n_338),
.Y(n_2688)
);

OAI21x1_ASAP7_75t_L g2689 ( 
.A1(n_2344),
.A2(n_337),
.B(n_339),
.Y(n_2689)
);

BUFx12f_ASAP7_75t_L g2690 ( 
.A(n_2514),
.Y(n_2690)
);

INVx8_ASAP7_75t_L g2691 ( 
.A(n_2457),
.Y(n_2691)
);

INVx2_ASAP7_75t_SL g2692 ( 
.A(n_2227),
.Y(n_2692)
);

OA21x2_ASAP7_75t_L g2693 ( 
.A1(n_2473),
.A2(n_340),
.B(n_342),
.Y(n_2693)
);

INVx4_ASAP7_75t_L g2694 ( 
.A(n_2457),
.Y(n_2694)
);

BUFx3_ASAP7_75t_L g2695 ( 
.A(n_2204),
.Y(n_2695)
);

NAND2x1p5_ASAP7_75t_L g2696 ( 
.A(n_2499),
.B(n_342),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2440),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2466),
.Y(n_2698)
);

BUFx12f_ASAP7_75t_L g2699 ( 
.A(n_2448),
.Y(n_2699)
);

BUFx3_ASAP7_75t_L g2700 ( 
.A(n_2155),
.Y(n_2700)
);

OAI21x1_ASAP7_75t_SL g2701 ( 
.A1(n_2312),
.A2(n_343),
.B(n_344),
.Y(n_2701)
);

OR2x6_ASAP7_75t_L g2702 ( 
.A(n_2184),
.B(n_343),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2159),
.B(n_344),
.Y(n_2703)
);

BUFx3_ASAP7_75t_L g2704 ( 
.A(n_2501),
.Y(n_2704)
);

AO21x2_ASAP7_75t_L g2705 ( 
.A1(n_2327),
.A2(n_345),
.B(n_347),
.Y(n_2705)
);

AO21x2_ASAP7_75t_L g2706 ( 
.A1(n_2281),
.A2(n_347),
.B(n_348),
.Y(n_2706)
);

BUFx2_ASAP7_75t_SL g2707 ( 
.A(n_2510),
.Y(n_2707)
);

OAI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2343),
.A2(n_350),
.B(n_352),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2596),
.B(n_352),
.Y(n_2709)
);

INVx3_ASAP7_75t_L g2710 ( 
.A(n_2499),
.Y(n_2710)
);

INVx2_ASAP7_75t_SL g2711 ( 
.A(n_2457),
.Y(n_2711)
);

AND2x4_ASAP7_75t_L g2712 ( 
.A(n_2195),
.B(n_2463),
.Y(n_2712)
);

AOI22xp5_ASAP7_75t_L g2713 ( 
.A1(n_2365),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2291),
.B(n_353),
.Y(n_2714)
);

OAI21xp5_ASAP7_75t_L g2715 ( 
.A1(n_2351),
.A2(n_354),
.B(n_355),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2455),
.Y(n_2716)
);

INVx3_ASAP7_75t_L g2717 ( 
.A(n_2513),
.Y(n_2717)
);

NAND2x1p5_ASAP7_75t_L g2718 ( 
.A(n_2513),
.B(n_357),
.Y(n_2718)
);

BUFx3_ASAP7_75t_L g2719 ( 
.A(n_2522),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2460),
.Y(n_2720)
);

AO21x2_ASAP7_75t_L g2721 ( 
.A1(n_2248),
.A2(n_358),
.B(n_359),
.Y(n_2721)
);

OAI21xp5_ASAP7_75t_L g2722 ( 
.A1(n_2309),
.A2(n_358),
.B(n_359),
.Y(n_2722)
);

OAI21x1_ASAP7_75t_L g2723 ( 
.A1(n_2226),
.A2(n_361),
.B(n_362),
.Y(n_2723)
);

AO21x2_ASAP7_75t_L g2724 ( 
.A1(n_2286),
.A2(n_362),
.B(n_363),
.Y(n_2724)
);

OAI21x1_ASAP7_75t_L g2725 ( 
.A1(n_2226),
.A2(n_365),
.B(n_366),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2520),
.Y(n_2726)
);

NAND2x1p5_ASAP7_75t_L g2727 ( 
.A(n_2516),
.B(n_368),
.Y(n_2727)
);

CKINVDCx11_ASAP7_75t_R g2728 ( 
.A(n_2586),
.Y(n_2728)
);

INVx3_ASAP7_75t_L g2729 ( 
.A(n_2516),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2479),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2160),
.B(n_368),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_SL g2732 ( 
.A(n_2385),
.B(n_369),
.Y(n_2732)
);

INVx4_ASAP7_75t_L g2733 ( 
.A(n_2463),
.Y(n_2733)
);

INVx1_ASAP7_75t_SL g2734 ( 
.A(n_2566),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2481),
.Y(n_2735)
);

BUFx6f_ASAP7_75t_L g2736 ( 
.A(n_2218),
.Y(n_2736)
);

BUFx3_ASAP7_75t_L g2737 ( 
.A(n_2208),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2528),
.Y(n_2738)
);

BUFx12f_ASAP7_75t_L g2739 ( 
.A(n_2572),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2161),
.B(n_371),
.Y(n_2740)
);

CKINVDCx20_ASAP7_75t_R g2741 ( 
.A(n_2252),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2222),
.B(n_372),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2539),
.Y(n_2743)
);

NAND2x1p5_ASAP7_75t_L g2744 ( 
.A(n_2531),
.B(n_374),
.Y(n_2744)
);

AOI22x1_ASAP7_75t_L g2745 ( 
.A1(n_2323),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_2745)
);

AND2x4_ASAP7_75t_L g2746 ( 
.A(n_2463),
.B(n_377),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2553),
.Y(n_2747)
);

NAND2x1p5_ASAP7_75t_L g2748 ( 
.A(n_2531),
.B(n_377),
.Y(n_2748)
);

INVx3_ASAP7_75t_SL g2749 ( 
.A(n_2511),
.Y(n_2749)
);

BUFx2_ASAP7_75t_L g2750 ( 
.A(n_2170),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2564),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2511),
.B(n_378),
.Y(n_2752)
);

INVxp67_ASAP7_75t_SL g2753 ( 
.A(n_2318),
.Y(n_2753)
);

BUFx12f_ASAP7_75t_L g2754 ( 
.A(n_2346),
.Y(n_2754)
);

AO21x2_ASAP7_75t_L g2755 ( 
.A1(n_2286),
.A2(n_2588),
.B(n_2476),
.Y(n_2755)
);

AO21x2_ASAP7_75t_L g2756 ( 
.A1(n_2429),
.A2(n_2238),
.B(n_2313),
.Y(n_2756)
);

BUFx4_ASAP7_75t_SL g2757 ( 
.A(n_2532),
.Y(n_2757)
);

AO21x2_ASAP7_75t_L g2758 ( 
.A1(n_2306),
.A2(n_2370),
.B(n_2376),
.Y(n_2758)
);

BUFx2_ASAP7_75t_L g2759 ( 
.A(n_2170),
.Y(n_2759)
);

HB1xp67_ASAP7_75t_L g2760 ( 
.A(n_2244),
.Y(n_2760)
);

NAND2x1p5_ASAP7_75t_L g2761 ( 
.A(n_2234),
.B(n_380),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2581),
.Y(n_2762)
);

OAI21xp5_ASAP7_75t_L g2763 ( 
.A1(n_2285),
.A2(n_380),
.B(n_381),
.Y(n_2763)
);

BUFx3_ASAP7_75t_L g2764 ( 
.A(n_2192),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2632),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2542),
.Y(n_2766)
);

CKINVDCx8_ASAP7_75t_R g2767 ( 
.A(n_2511),
.Y(n_2767)
);

AO21x2_ASAP7_75t_L g2768 ( 
.A1(n_2611),
.A2(n_382),
.B(n_383),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2549),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2552),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2565),
.Y(n_2771)
);

BUFx3_ASAP7_75t_L g2772 ( 
.A(n_2310),
.Y(n_2772)
);

CKINVDCx5p33_ASAP7_75t_R g2773 ( 
.A(n_2361),
.Y(n_2773)
);

OAI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_2274),
.A2(n_384),
.B(n_385),
.Y(n_2774)
);

AO21x2_ASAP7_75t_L g2775 ( 
.A1(n_2307),
.A2(n_386),
.B(n_387),
.Y(n_2775)
);

BUFx6f_ASAP7_75t_L g2776 ( 
.A(n_2250),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2582),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2598),
.Y(n_2778)
);

BUFx3_ASAP7_75t_L g2779 ( 
.A(n_2209),
.Y(n_2779)
);

NAND3xp33_ASAP7_75t_L g2780 ( 
.A(n_2289),
.B(n_386),
.C(n_387),
.Y(n_2780)
);

OA21x2_ASAP7_75t_L g2781 ( 
.A1(n_2392),
.A2(n_388),
.B(n_389),
.Y(n_2781)
);

BUFx3_ASAP7_75t_L g2782 ( 
.A(n_2267),
.Y(n_2782)
);

AND2x4_ASAP7_75t_L g2783 ( 
.A(n_2350),
.B(n_388),
.Y(n_2783)
);

BUFx3_ASAP7_75t_L g2784 ( 
.A(n_2249),
.Y(n_2784)
);

BUFx3_ASAP7_75t_L g2785 ( 
.A(n_2271),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2599),
.Y(n_2786)
);

INVx5_ASAP7_75t_SL g2787 ( 
.A(n_2532),
.Y(n_2787)
);

AO21x2_ASAP7_75t_L g2788 ( 
.A1(n_2319),
.A2(n_389),
.B(n_391),
.Y(n_2788)
);

BUFx5_ASAP7_75t_L g2789 ( 
.A(n_2600),
.Y(n_2789)
);

OR2x2_ASAP7_75t_L g2790 ( 
.A(n_2162),
.B(n_392),
.Y(n_2790)
);

BUFx6f_ASAP7_75t_L g2791 ( 
.A(n_2250),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2613),
.Y(n_2792)
);

AO21x2_ASAP7_75t_L g2793 ( 
.A1(n_2335),
.A2(n_393),
.B(n_394),
.Y(n_2793)
);

INVxp67_ASAP7_75t_L g2794 ( 
.A(n_2566),
.Y(n_2794)
);

INVx2_ASAP7_75t_SL g2795 ( 
.A(n_2176),
.Y(n_2795)
);

NAND2x1p5_ASAP7_75t_L g2796 ( 
.A(n_2234),
.B(n_395),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2614),
.Y(n_2797)
);

HB1xp67_ASAP7_75t_L g2798 ( 
.A(n_2244),
.Y(n_2798)
);

BUFx3_ASAP7_75t_L g2799 ( 
.A(n_2450),
.Y(n_2799)
);

BUFx3_ASAP7_75t_L g2800 ( 
.A(n_2474),
.Y(n_2800)
);

INVx4_ASAP7_75t_L g2801 ( 
.A(n_2600),
.Y(n_2801)
);

OAI21xp5_ASAP7_75t_L g2802 ( 
.A1(n_2183),
.A2(n_397),
.B(n_398),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2617),
.Y(n_2803)
);

OAI21x1_ASAP7_75t_L g2804 ( 
.A1(n_2412),
.A2(n_400),
.B(n_401),
.Y(n_2804)
);

INVx6_ASAP7_75t_SL g2805 ( 
.A(n_2574),
.Y(n_2805)
);

INVx3_ASAP7_75t_L g2806 ( 
.A(n_2175),
.Y(n_2806)
);

OAI21xp5_ASAP7_75t_L g2807 ( 
.A1(n_2247),
.A2(n_2256),
.B(n_2255),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2628),
.Y(n_2808)
);

OAI21x1_ASAP7_75t_L g2809 ( 
.A1(n_2411),
.A2(n_403),
.B(n_404),
.Y(n_2809)
);

AOI22x1_ASAP7_75t_L g2810 ( 
.A1(n_2363),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_2810)
);

INVx3_ASAP7_75t_L g2811 ( 
.A(n_2175),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2629),
.Y(n_2812)
);

BUFx3_ASAP7_75t_L g2813 ( 
.A(n_2623),
.Y(n_2813)
);

OAI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_2147),
.A2(n_407),
.B(n_408),
.Y(n_2814)
);

BUFx6f_ASAP7_75t_L g2815 ( 
.A(n_2250),
.Y(n_2815)
);

OAI21x1_ASAP7_75t_L g2816 ( 
.A1(n_2489),
.A2(n_409),
.B(n_410),
.Y(n_2816)
);

OAI21x1_ASAP7_75t_L g2817 ( 
.A1(n_2489),
.A2(n_411),
.B(n_412),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2182),
.Y(n_2818)
);

OAI21x1_ASAP7_75t_L g2819 ( 
.A1(n_2550),
.A2(n_411),
.B(n_413),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2188),
.Y(n_2820)
);

INVx2_ASAP7_75t_SL g2821 ( 
.A(n_2328),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2202),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2216),
.Y(n_2823)
);

OA21x2_ASAP7_75t_L g2824 ( 
.A1(n_2445),
.A2(n_413),
.B(n_414),
.Y(n_2824)
);

INVx3_ASAP7_75t_SL g2825 ( 
.A(n_2574),
.Y(n_2825)
);

AND2x2_ASAP7_75t_SL g2826 ( 
.A(n_2401),
.B(n_414),
.Y(n_2826)
);

OAI21x1_ASAP7_75t_L g2827 ( 
.A1(n_2550),
.A2(n_415),
.B(n_416),
.Y(n_2827)
);

AND2x4_ASAP7_75t_L g2828 ( 
.A(n_2375),
.B(n_416),
.Y(n_2828)
);

CKINVDCx5p33_ASAP7_75t_R g2829 ( 
.A(n_2164),
.Y(n_2829)
);

HB1xp67_ASAP7_75t_L g2830 ( 
.A(n_2244),
.Y(n_2830)
);

OAI21x1_ASAP7_75t_SL g2831 ( 
.A1(n_2443),
.A2(n_417),
.B(n_418),
.Y(n_2831)
);

INVx3_ASAP7_75t_SL g2832 ( 
.A(n_2487),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2321),
.Y(n_2833)
);

CKINVDCx20_ASAP7_75t_R g2834 ( 
.A(n_2199),
.Y(n_2834)
);

OAI21x1_ASAP7_75t_L g2835 ( 
.A1(n_2562),
.A2(n_418),
.B(n_419),
.Y(n_2835)
);

NOR2xp67_ASAP7_75t_L g2836 ( 
.A(n_2288),
.B(n_419),
.Y(n_2836)
);

BUFx2_ASAP7_75t_L g2837 ( 
.A(n_2633),
.Y(n_2837)
);

OAI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2355),
.A2(n_420),
.B(n_421),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2329),
.Y(n_2839)
);

AO21x2_ASAP7_75t_L g2840 ( 
.A1(n_2345),
.A2(n_2352),
.B(n_2349),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2229),
.Y(n_2841)
);

CKINVDCx5p33_ASAP7_75t_R g2842 ( 
.A(n_2258),
.Y(n_2842)
);

INVx8_ASAP7_75t_L g2843 ( 
.A(n_2600),
.Y(n_2843)
);

OAI21x1_ASAP7_75t_SL g2844 ( 
.A1(n_2444),
.A2(n_421),
.B(n_422),
.Y(n_2844)
);

BUFx2_ASAP7_75t_SL g2845 ( 
.A(n_2600),
.Y(n_2845)
);

HB1xp67_ASAP7_75t_L g2846 ( 
.A(n_2288),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2196),
.B(n_422),
.Y(n_2847)
);

AO21x2_ASAP7_75t_L g2848 ( 
.A1(n_2353),
.A2(n_423),
.B(n_424),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2292),
.Y(n_2849)
);

BUFx2_ASAP7_75t_L g2850 ( 
.A(n_2215),
.Y(n_2850)
);

OAI21x1_ASAP7_75t_L g2851 ( 
.A1(n_2262),
.A2(n_423),
.B(n_424),
.Y(n_2851)
);

OAI21xp5_ASAP7_75t_L g2852 ( 
.A1(n_2149),
.A2(n_425),
.B(n_426),
.Y(n_2852)
);

OAI21x1_ASAP7_75t_L g2853 ( 
.A1(n_2264),
.A2(n_425),
.B(n_426),
.Y(n_2853)
);

CKINVDCx11_ASAP7_75t_R g2854 ( 
.A(n_2340),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2297),
.Y(n_2855)
);

HB1xp67_ASAP7_75t_L g2856 ( 
.A(n_2288),
.Y(n_2856)
);

AO21x2_ASAP7_75t_L g2857 ( 
.A1(n_2356),
.A2(n_427),
.B(n_428),
.Y(n_2857)
);

BUFx2_ASAP7_75t_R g2858 ( 
.A(n_2406),
.Y(n_2858)
);

AOI22x1_ASAP7_75t_L g2859 ( 
.A1(n_2371),
.A2(n_429),
.B1(n_427),
.B2(n_428),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2338),
.Y(n_2860)
);

BUFx12f_ASAP7_75t_L g2861 ( 
.A(n_2346),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2298),
.Y(n_2862)
);

INVx4_ASAP7_75t_L g2863 ( 
.A(n_2365),
.Y(n_2863)
);

BUFx12f_ASAP7_75t_L g2864 ( 
.A(n_2251),
.Y(n_2864)
);

INVx3_ASAP7_75t_SL g2865 ( 
.A(n_2608),
.Y(n_2865)
);

INVx4_ASAP7_75t_L g2866 ( 
.A(n_2382),
.Y(n_2866)
);

OAI21x1_ASAP7_75t_L g2867 ( 
.A1(n_2402),
.A2(n_429),
.B(n_430),
.Y(n_2867)
);

INVx4_ASAP7_75t_L g2868 ( 
.A(n_2382),
.Y(n_2868)
);

OR2x6_ASAP7_75t_L g2869 ( 
.A(n_2191),
.B(n_430),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2330),
.Y(n_2870)
);

NAND2x1p5_ASAP7_75t_L g2871 ( 
.A(n_2300),
.B(n_431),
.Y(n_2871)
);

NAND2x1p5_ASAP7_75t_L g2872 ( 
.A(n_2400),
.B(n_433),
.Y(n_2872)
);

BUFx2_ASAP7_75t_L g2873 ( 
.A(n_2472),
.Y(n_2873)
);

BUFx2_ASAP7_75t_SL g2874 ( 
.A(n_2451),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2359),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2240),
.B(n_434),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2304),
.Y(n_2877)
);

BUFx12f_ASAP7_75t_L g2878 ( 
.A(n_2458),
.Y(n_2878)
);

INVx3_ASAP7_75t_L g2879 ( 
.A(n_2293),
.Y(n_2879)
);

AOI22x1_ASAP7_75t_L g2880 ( 
.A1(n_2471),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2339),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2172),
.B(n_436),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2243),
.B(n_2314),
.Y(n_2883)
);

INVx2_ASAP7_75t_SL g2884 ( 
.A(n_2268),
.Y(n_2884)
);

OAI21xp5_ASAP7_75t_L g2885 ( 
.A1(n_2449),
.A2(n_438),
.B(n_439),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2433),
.Y(n_2886)
);

OAI21x1_ASAP7_75t_SL g2887 ( 
.A1(n_2454),
.A2(n_439),
.B(n_440),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2357),
.Y(n_2888)
);

BUFx3_ASAP7_75t_L g2889 ( 
.A(n_2317),
.Y(n_2889)
);

OAI21x1_ASAP7_75t_L g2890 ( 
.A1(n_2270),
.A2(n_440),
.B(n_442),
.Y(n_2890)
);

BUFx3_ASAP7_75t_L g2891 ( 
.A(n_2495),
.Y(n_2891)
);

OAI21x1_ASAP7_75t_L g2892 ( 
.A1(n_2270),
.A2(n_443),
.B(n_444),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2524),
.Y(n_2893)
);

NAND2x1_ASAP7_75t_L g2894 ( 
.A(n_2315),
.B(n_445),
.Y(n_2894)
);

OAI21x1_ASAP7_75t_SL g2895 ( 
.A1(n_2456),
.A2(n_445),
.B(n_446),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2536),
.Y(n_2896)
);

BUFx2_ASAP7_75t_R g2897 ( 
.A(n_2287),
.Y(n_2897)
);

BUFx12f_ASAP7_75t_L g2898 ( 
.A(n_2605),
.Y(n_2898)
);

BUFx2_ASAP7_75t_L g2899 ( 
.A(n_2478),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2419),
.Y(n_2900)
);

INVx1_ASAP7_75t_SL g2901 ( 
.A(n_2268),
.Y(n_2901)
);

OAI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2461),
.A2(n_449),
.B(n_450),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2442),
.Y(n_2903)
);

AND2x6_ASAP7_75t_L g2904 ( 
.A(n_2467),
.B(n_449),
.Y(n_2904)
);

INVx4_ASAP7_75t_L g2905 ( 
.A(n_2467),
.Y(n_2905)
);

BUFx3_ASAP7_75t_L g2906 ( 
.A(n_2631),
.Y(n_2906)
);

OR2x6_ASAP7_75t_L g2907 ( 
.A(n_2388),
.B(n_450),
.Y(n_2907)
);

INVxp67_ASAP7_75t_SL g2908 ( 
.A(n_2468),
.Y(n_2908)
);

AO21x2_ASAP7_75t_L g2909 ( 
.A1(n_2360),
.A2(n_451),
.B(n_452),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2213),
.Y(n_2910)
);

BUFx3_ASAP7_75t_L g2911 ( 
.A(n_2409),
.Y(n_2911)
);

INVxp67_ASAP7_75t_SL g2912 ( 
.A(n_2468),
.Y(n_2912)
);

INVx1_ASAP7_75t_SL g2913 ( 
.A(n_2391),
.Y(n_2913)
);

INVx1_ASAP7_75t_SL g2914 ( 
.A(n_2420),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2259),
.Y(n_2915)
);

INVx6_ASAP7_75t_L g2916 ( 
.A(n_2379),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2367),
.Y(n_2917)
);

OAI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2464),
.A2(n_456),
.B(n_457),
.Y(n_2918)
);

INVx2_ASAP7_75t_SL g2919 ( 
.A(n_2272),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2213),
.Y(n_2920)
);

AO21x2_ASAP7_75t_L g2921 ( 
.A1(n_2242),
.A2(n_2428),
.B(n_2386),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2236),
.Y(n_2922)
);

HB1xp67_ASAP7_75t_L g2923 ( 
.A(n_2206),
.Y(n_2923)
);

NAND2x1p5_ASAP7_75t_L g2924 ( 
.A(n_2439),
.B(n_457),
.Y(n_2924)
);

INVx1_ASAP7_75t_SL g2925 ( 
.A(n_2431),
.Y(n_2925)
);

AOI21xp5_ASAP7_75t_L g2926 ( 
.A1(n_2294),
.A2(n_2480),
.B(n_2469),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2280),
.Y(n_2927)
);

INVx5_ASAP7_75t_SL g2928 ( 
.A(n_2396),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2279),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2301),
.Y(n_2930)
);

BUFx3_ASAP7_75t_L g2931 ( 
.A(n_2295),
.Y(n_2931)
);

NAND2x1p5_ASAP7_75t_L g2932 ( 
.A(n_2607),
.B(n_458),
.Y(n_2932)
);

AO21x2_ASAP7_75t_L g2933 ( 
.A1(n_2494),
.A2(n_458),
.B(n_459),
.Y(n_2933)
);

AO21x2_ASAP7_75t_L g2934 ( 
.A1(n_2535),
.A2(n_459),
.B(n_460),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2235),
.B(n_460),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2166),
.B(n_461),
.Y(n_2936)
);

AOI21xp5_ASAP7_75t_L g2937 ( 
.A1(n_2482),
.A2(n_461),
.B(n_462),
.Y(n_2937)
);

INVx2_ASAP7_75t_SL g2938 ( 
.A(n_2158),
.Y(n_2938)
);

BUFx5_ASAP7_75t_L g2939 ( 
.A(n_2377),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2302),
.Y(n_2940)
);

AOI22x1_ASAP7_75t_L g2941 ( 
.A1(n_2530),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_2941)
);

BUFx3_ASAP7_75t_L g2942 ( 
.A(n_2626),
.Y(n_2942)
);

BUFx3_ASAP7_75t_L g2943 ( 
.A(n_2198),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2305),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2166),
.B(n_463),
.Y(n_2945)
);

BUFx4_ASAP7_75t_SL g2946 ( 
.A(n_2396),
.Y(n_2946)
);

INVx8_ASAP7_75t_L g2947 ( 
.A(n_2198),
.Y(n_2947)
);

OAI21xp5_ASAP7_75t_L g2948 ( 
.A1(n_2485),
.A2(n_2498),
.B(n_2497),
.Y(n_2948)
);

OR2x6_ASAP7_75t_L g2949 ( 
.A(n_2296),
.B(n_465),
.Y(n_2949)
);

CKINVDCx20_ASAP7_75t_R g2950 ( 
.A(n_2277),
.Y(n_2950)
);

NAND2x1p5_ASAP7_75t_L g2951 ( 
.A(n_2475),
.B(n_466),
.Y(n_2951)
);

AO21x2_ASAP7_75t_L g2952 ( 
.A1(n_2537),
.A2(n_466),
.B(n_467),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2432),
.Y(n_2953)
);

BUFx3_ASAP7_75t_L g2954 ( 
.A(n_2278),
.Y(n_2954)
);

INVx4_ASAP7_75t_L g2955 ( 
.A(n_2483),
.Y(n_2955)
);

CKINVDCx14_ASAP7_75t_R g2956 ( 
.A(n_2621),
.Y(n_2956)
);

AND2x4_ASAP7_75t_L g2957 ( 
.A(n_2394),
.B(n_469),
.Y(n_2957)
);

AO21x2_ASAP7_75t_L g2958 ( 
.A1(n_2546),
.A2(n_469),
.B(n_470),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2500),
.B(n_470),
.Y(n_2959)
);

INVx5_ASAP7_75t_L g2960 ( 
.A(n_2483),
.Y(n_2960)
);

OA21x2_ASAP7_75t_L g2961 ( 
.A1(n_2541),
.A2(n_2570),
.B(n_2548),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2503),
.B(n_472),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2246),
.Y(n_2963)
);

OR2x6_ASAP7_75t_L g2964 ( 
.A(n_2241),
.B(n_473),
.Y(n_2964)
);

OA21x2_ASAP7_75t_L g2965 ( 
.A1(n_2576),
.A2(n_2579),
.B(n_2578),
.Y(n_2965)
);

INVx5_ASAP7_75t_L g2966 ( 
.A(n_2483),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2273),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2282),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2508),
.B(n_474),
.Y(n_2969)
);

BUFx3_ASAP7_75t_L g2970 ( 
.A(n_2405),
.Y(n_2970)
);

AO21x2_ASAP7_75t_L g2971 ( 
.A1(n_2569),
.A2(n_474),
.B(n_475),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2342),
.Y(n_2972)
);

BUFx4f_ASAP7_75t_L g2973 ( 
.A(n_2398),
.Y(n_2973)
);

AND2x4_ASAP7_75t_SL g2974 ( 
.A(n_2490),
.B(n_477),
.Y(n_2974)
);

OAI21xp5_ASAP7_75t_L g2975 ( 
.A1(n_2525),
.A2(n_479),
.B(n_480),
.Y(n_2975)
);

INVx2_ASAP7_75t_SL g2976 ( 
.A(n_2493),
.Y(n_2976)
);

AO21x2_ASAP7_75t_L g2977 ( 
.A1(n_2590),
.A2(n_481),
.B(n_483),
.Y(n_2977)
);

NOR2x1_ASAP7_75t_R g2978 ( 
.A(n_2398),
.B(n_481),
.Y(n_2978)
);

OAI21xp5_ASAP7_75t_L g2979 ( 
.A1(n_2533),
.A2(n_483),
.B(n_484),
.Y(n_2979)
);

AOI21x1_ASAP7_75t_L g2980 ( 
.A1(n_2366),
.A2(n_486),
.B(n_487),
.Y(n_2980)
);

AND2x4_ASAP7_75t_L g2981 ( 
.A(n_2422),
.B(n_487),
.Y(n_2981)
);

BUFx4_ASAP7_75t_SL g2982 ( 
.A(n_2430),
.Y(n_2982)
);

BUFx12f_ASAP7_75t_L g2983 ( 
.A(n_2381),
.Y(n_2983)
);

AO21x2_ASAP7_75t_L g2984 ( 
.A1(n_2595),
.A2(n_488),
.B(n_491),
.Y(n_2984)
);

AO21x2_ASAP7_75t_L g2985 ( 
.A1(n_2616),
.A2(n_2625),
.B(n_2620),
.Y(n_2985)
);

BUFx3_ASAP7_75t_L g2986 ( 
.A(n_2538),
.Y(n_2986)
);

INVx1_ASAP7_75t_SL g2987 ( 
.A(n_2491),
.Y(n_2987)
);

AO21x2_ASAP7_75t_L g2988 ( 
.A1(n_2534),
.A2(n_494),
.B(n_496),
.Y(n_2988)
);

OAI21xp5_ASAP7_75t_L g2989 ( 
.A1(n_2544),
.A2(n_494),
.B(n_496),
.Y(n_2989)
);

OA21x2_ASAP7_75t_L g2990 ( 
.A1(n_2265),
.A2(n_497),
.B(n_499),
.Y(n_2990)
);

INVx2_ASAP7_75t_SL g2991 ( 
.A(n_2303),
.Y(n_2991)
);

BUFx6f_ASAP7_75t_L g2992 ( 
.A(n_2491),
.Y(n_2992)
);

AO21x2_ASAP7_75t_L g2993 ( 
.A1(n_2547),
.A2(n_497),
.B(n_499),
.Y(n_2993)
);

INVxp67_ASAP7_75t_SL g2994 ( 
.A(n_2609),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2320),
.Y(n_2995)
);

BUFx3_ASAP7_75t_L g2996 ( 
.A(n_2303),
.Y(n_2996)
);

AO21x2_ASAP7_75t_L g2997 ( 
.A1(n_2555),
.A2(n_500),
.B(n_501),
.Y(n_2997)
);

OAI21x1_ASAP7_75t_L g2998 ( 
.A1(n_2414),
.A2(n_500),
.B(n_501),
.Y(n_2998)
);

NAND2x1p5_ASAP7_75t_L g2999 ( 
.A(n_2609),
.B(n_502),
.Y(n_2999)
);

OR2x2_ASAP7_75t_L g3000 ( 
.A(n_2245),
.B(n_502),
.Y(n_3000)
);

INVxp67_ASAP7_75t_L g3001 ( 
.A(n_2612),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2322),
.Y(n_3002)
);

AO21x2_ASAP7_75t_L g3003 ( 
.A1(n_2557),
.A2(n_503),
.B(n_504),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2368),
.Y(n_3004)
);

AO21x2_ASAP7_75t_L g3005 ( 
.A1(n_2583),
.A2(n_503),
.B(n_505),
.Y(n_3005)
);

OAI21x1_ASAP7_75t_L g3006 ( 
.A1(n_2415),
.A2(n_505),
.B(n_508),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2137),
.B(n_508),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2585),
.B(n_510),
.Y(n_3008)
);

NAND2x1p5_ASAP7_75t_L g3009 ( 
.A(n_2326),
.B(n_510),
.Y(n_3009)
);

INVx5_ASAP7_75t_L g3010 ( 
.A(n_2435),
.Y(n_3010)
);

BUFx12f_ASAP7_75t_L g3011 ( 
.A(n_2403),
.Y(n_3011)
);

BUFx2_ASAP7_75t_L g3012 ( 
.A(n_2447),
.Y(n_3012)
);

NOR2x1_ASAP7_75t_L g3013 ( 
.A(n_2146),
.B(n_511),
.Y(n_3013)
);

BUFx2_ASAP7_75t_L g3014 ( 
.A(n_2378),
.Y(n_3014)
);

INVx4_ASAP7_75t_L g3015 ( 
.A(n_2311),
.Y(n_3015)
);

CKINVDCx5p33_ASAP7_75t_R g3016 ( 
.A(n_2207),
.Y(n_3016)
);

OR2x6_ASAP7_75t_L g3017 ( 
.A(n_2200),
.B(n_514),
.Y(n_3017)
);

BUFx12f_ASAP7_75t_L g3018 ( 
.A(n_2403),
.Y(n_3018)
);

BUFx3_ASAP7_75t_L g3019 ( 
.A(n_2311),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2324),
.Y(n_3020)
);

BUFx12f_ASAP7_75t_L g3021 ( 
.A(n_2413),
.Y(n_3021)
);

OAI21x1_ASAP7_75t_L g3022 ( 
.A1(n_2404),
.A2(n_515),
.B(n_516),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2154),
.Y(n_3023)
);

AO21x2_ASAP7_75t_L g3024 ( 
.A1(n_2597),
.A2(n_516),
.B(n_517),
.Y(n_3024)
);

AO21x2_ASAP7_75t_L g3025 ( 
.A1(n_2602),
.A2(n_517),
.B(n_518),
.Y(n_3025)
);

OAI21x1_ASAP7_75t_SL g3026 ( 
.A1(n_2604),
.A2(n_519),
.B(n_520),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2615),
.B(n_520),
.Y(n_3027)
);

NAND2x1p5_ASAP7_75t_L g3028 ( 
.A(n_2435),
.B(n_521),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2354),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2369),
.Y(n_3030)
);

OAI21xp5_ASAP7_75t_L g3031 ( 
.A1(n_2618),
.A2(n_521),
.B(n_523),
.Y(n_3031)
);

BUFx2_ASAP7_75t_L g3032 ( 
.A(n_2331),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2390),
.Y(n_3033)
);

AND2x4_ASAP7_75t_L g3034 ( 
.A(n_2373),
.B(n_523),
.Y(n_3034)
);

CKINVDCx5p33_ASAP7_75t_R g3035 ( 
.A(n_2141),
.Y(n_3035)
);

NAND3xp33_ASAP7_75t_L g3036 ( 
.A(n_2260),
.B(n_524),
.C(n_525),
.Y(n_3036)
);

AND2x4_ASAP7_75t_L g3037 ( 
.A(n_2364),
.B(n_527),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2261),
.Y(n_3038)
);

AO21x2_ASAP7_75t_L g3039 ( 
.A1(n_2232),
.A2(n_2395),
.B(n_2384),
.Y(n_3039)
);

INVx1_ASAP7_75t_SL g3040 ( 
.A(n_2275),
.Y(n_3040)
);

NAND2x1p5_ASAP7_75t_L g3041 ( 
.A(n_2181),
.B(n_527),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2139),
.B(n_528),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2266),
.B(n_528),
.Y(n_3043)
);

NAND2x1p5_ASAP7_75t_L g3044 ( 
.A(n_2237),
.B(n_529),
.Y(n_3044)
);

AND2x4_ASAP7_75t_L g3045 ( 
.A(n_2269),
.B(n_529),
.Y(n_3045)
);

INVx3_ASAP7_75t_L g3046 ( 
.A(n_2407),
.Y(n_3046)
);

BUFx8_ASAP7_75t_L g3047 ( 
.A(n_2523),
.Y(n_3047)
);

HB1xp67_ASAP7_75t_L g3048 ( 
.A(n_2206),
.Y(n_3048)
);

BUFx4f_ASAP7_75t_L g3049 ( 
.A(n_2492),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2276),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2283),
.B(n_530),
.Y(n_3051)
);

INVx4_ASAP7_75t_L g3052 ( 
.A(n_2231),
.Y(n_3052)
);

BUFx12f_ASAP7_75t_L g3053 ( 
.A(n_2152),
.Y(n_3053)
);

OAI21xp5_ASAP7_75t_L g3054 ( 
.A1(n_2189),
.A2(n_532),
.B(n_533),
.Y(n_3054)
);

AOI21x1_ASAP7_75t_L g3055 ( 
.A1(n_2399),
.A2(n_533),
.B(n_534),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2284),
.Y(n_3056)
);

AOI22x1_ASAP7_75t_L g3057 ( 
.A1(n_2194),
.A2(n_537),
.B1(n_534),
.B2(n_536),
.Y(n_3057)
);

AND2x4_ASAP7_75t_L g3058 ( 
.A(n_2425),
.B(n_537),
.Y(n_3058)
);

OAI21xp5_ASAP7_75t_L g3059 ( 
.A1(n_2257),
.A2(n_540),
.B(n_541),
.Y(n_3059)
);

BUFx2_ASAP7_75t_SL g3060 ( 
.A(n_2165),
.Y(n_3060)
);

BUFx4f_ASAP7_75t_SL g3061 ( 
.A(n_2462),
.Y(n_3061)
);

AO21x2_ASAP7_75t_L g3062 ( 
.A1(n_2427),
.A2(n_540),
.B(n_542),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2142),
.Y(n_3063)
);

AO21x2_ASAP7_75t_L g3064 ( 
.A1(n_2426),
.A2(n_543),
.B(n_544),
.Y(n_3064)
);

INVx4_ASAP7_75t_L g3065 ( 
.A(n_2423),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2417),
.Y(n_3066)
);

BUFx6f_ASAP7_75t_L g3067 ( 
.A(n_2418),
.Y(n_3067)
);

BUFx2_ASAP7_75t_L g3068 ( 
.A(n_2484),
.Y(n_3068)
);

AND2x4_ASAP7_75t_L g3069 ( 
.A(n_2372),
.B(n_545),
.Y(n_3069)
);

AOI22xp33_ASAP7_75t_L g3070 ( 
.A1(n_2253),
.A2(n_2348),
.B1(n_2453),
.B2(n_2437),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_SL g3071 ( 
.A(n_2484),
.B(n_547),
.Y(n_3071)
);

OAI21x1_ASAP7_75t_SL g3072 ( 
.A1(n_2299),
.A2(n_547),
.B(n_548),
.Y(n_3072)
);

AO21x2_ASAP7_75t_L g3073 ( 
.A1(n_2316),
.A2(n_550),
.B(n_551),
.Y(n_3073)
);

OA21x2_ASAP7_75t_L g3074 ( 
.A1(n_2336),
.A2(n_550),
.B(n_551),
.Y(n_3074)
);

INVx3_ASAP7_75t_L g3075 ( 
.A(n_2387),
.Y(n_3075)
);

INVx3_ASAP7_75t_SL g3076 ( 
.A(n_2193),
.Y(n_3076)
);

OAI21xp5_ASAP7_75t_L g3077 ( 
.A1(n_2163),
.A2(n_552),
.B(n_553),
.Y(n_3077)
);

AOI22xp33_ASAP7_75t_L g3078 ( 
.A1(n_2826),
.A2(n_2512),
.B1(n_2529),
.B2(n_2502),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2636),
.Y(n_3079)
);

BUFx8_ASAP7_75t_L g3080 ( 
.A(n_2645),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2923),
.Y(n_3081)
);

BUFx3_ASAP7_75t_L g3082 ( 
.A(n_2782),
.Y(n_3082)
);

BUFx3_ASAP7_75t_L g3083 ( 
.A(n_2668),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_3023),
.B(n_2543),
.Y(n_3084)
);

AOI22xp5_ASAP7_75t_L g3085 ( 
.A1(n_2826),
.A2(n_2180),
.B1(n_2214),
.B2(n_2224),
.Y(n_3085)
);

AOI22xp33_ASAP7_75t_L g3086 ( 
.A1(n_3049),
.A2(n_2863),
.B1(n_2732),
.B2(n_2927),
.Y(n_3086)
);

AO21x1_ASAP7_75t_L g3087 ( 
.A1(n_2732),
.A2(n_2434),
.B(n_2389),
.Y(n_3087)
);

CKINVDCx11_ASAP7_75t_R g3088 ( 
.A(n_2686),
.Y(n_3088)
);

INVx1_ASAP7_75t_SL g3089 ( 
.A(n_2741),
.Y(n_3089)
);

AOI22xp33_ASAP7_75t_SL g3090 ( 
.A1(n_2863),
.A2(n_2601),
.B1(n_2410),
.B2(n_2436),
.Y(n_3090)
);

CKINVDCx20_ASAP7_75t_R g3091 ( 
.A(n_2741),
.Y(n_3091)
);

BUFx10_ASAP7_75t_L g3092 ( 
.A(n_2773),
.Y(n_3092)
);

AOI22xp33_ASAP7_75t_L g3093 ( 
.A1(n_3049),
.A2(n_2571),
.B1(n_2592),
.B2(n_2554),
.Y(n_3093)
);

OAI21xp5_ASAP7_75t_SL g3094 ( 
.A1(n_2956),
.A2(n_2559),
.B(n_2587),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2923),
.Y(n_3095)
);

AND2x2_ASAP7_75t_L g3096 ( 
.A(n_2883),
.B(n_2577),
.Y(n_3096)
);

AOI22xp33_ASAP7_75t_L g3097 ( 
.A1(n_2963),
.A2(n_2634),
.B1(n_2635),
.B2(n_2603),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_3048),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_3048),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2643),
.Y(n_3100)
);

BUFx12f_ASAP7_75t_L g3101 ( 
.A(n_2728),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_2637),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2638),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_2671),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2675),
.Y(n_3105)
);

BUFx6f_ASAP7_75t_L g3106 ( 
.A(n_2960),
.Y(n_3106)
);

NAND2x1p5_ASAP7_75t_L g3107 ( 
.A(n_2687),
.B(n_2212),
.Y(n_3107)
);

CKINVDCx11_ASAP7_75t_R g3108 ( 
.A(n_2728),
.Y(n_3108)
);

HB1xp67_ASAP7_75t_L g3109 ( 
.A(n_2644),
.Y(n_3109)
);

BUFx5_ASAP7_75t_L g3110 ( 
.A(n_2904),
.Y(n_3110)
);

AOI22xp33_ASAP7_75t_L g3111 ( 
.A1(n_3004),
.A2(n_2358),
.B1(n_2333),
.B2(n_2374),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2917),
.B(n_2239),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_2647),
.B(n_2589),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_2973),
.A2(n_2408),
.B1(n_2416),
.B2(n_2507),
.Y(n_3114)
);

BUFx6f_ASAP7_75t_L g3115 ( 
.A(n_2960),
.Y(n_3115)
);

INVx4_ASAP7_75t_L g3116 ( 
.A(n_2843),
.Y(n_3116)
);

HB1xp67_ASAP7_75t_L g3117 ( 
.A(n_2644),
.Y(n_3117)
);

OAI22xp33_ASAP7_75t_L g3118 ( 
.A1(n_3017),
.A2(n_2397),
.B1(n_2504),
.B2(n_2488),
.Y(n_3118)
);

CKINVDCx5p33_ASAP7_75t_R g3119 ( 
.A(n_2946),
.Y(n_3119)
);

OAI22xp5_ASAP7_75t_L g3120 ( 
.A1(n_2652),
.A2(n_2334),
.B1(n_2506),
.B2(n_2477),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_2936),
.B(n_2622),
.Y(n_3121)
);

AO21x2_ASAP7_75t_L g3122 ( 
.A1(n_2910),
.A2(n_2575),
.B(n_2220),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2677),
.Y(n_3123)
);

AOI22xp33_ASAP7_75t_L g3124 ( 
.A1(n_2973),
.A2(n_2509),
.B1(n_2526),
.B2(n_2515),
.Y(n_3124)
);

OAI21x1_ASAP7_75t_L g3125 ( 
.A1(n_2685),
.A2(n_2421),
.B(n_2223),
.Y(n_3125)
);

CKINVDCx11_ASAP7_75t_R g3126 ( 
.A(n_2639),
.Y(n_3126)
);

BUFx6f_ASAP7_75t_L g3127 ( 
.A(n_2960),
.Y(n_3127)
);

AOI22xp33_ASAP7_75t_L g3128 ( 
.A1(n_3047),
.A2(n_2545),
.B1(n_2556),
.B2(n_2551),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2659),
.Y(n_3129)
);

NOR2x1_ASAP7_75t_SL g3130 ( 
.A(n_2845),
.B(n_2561),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2666),
.Y(n_3131)
);

BUFx2_ASAP7_75t_L g3132 ( 
.A(n_2805),
.Y(n_3132)
);

BUFx2_ASAP7_75t_L g3133 ( 
.A(n_2805),
.Y(n_3133)
);

INVx4_ASAP7_75t_L g3134 ( 
.A(n_2843),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2680),
.Y(n_3135)
);

OAI22xp33_ASAP7_75t_L g3136 ( 
.A1(n_3017),
.A2(n_2505),
.B1(n_2519),
.B2(n_2518),
.Y(n_3136)
);

OAI22xp5_ASAP7_75t_L g3137 ( 
.A1(n_2652),
.A2(n_2347),
.B1(n_2567),
.B2(n_2563),
.Y(n_3137)
);

AOI21x1_ASAP7_75t_L g3138 ( 
.A1(n_2926),
.A2(n_2593),
.B(n_2219),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2698),
.Y(n_3139)
);

CKINVDCx11_ASAP7_75t_R g3140 ( 
.A(n_2690),
.Y(n_3140)
);

HB1xp67_ASAP7_75t_L g3141 ( 
.A(n_2679),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2672),
.Y(n_3142)
);

INVx6_ASAP7_75t_L g3143 ( 
.A(n_2691),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2681),
.Y(n_3144)
);

AOI22xp33_ASAP7_75t_SL g3145 ( 
.A1(n_2956),
.A2(n_2601),
.B1(n_2521),
.B2(n_2540),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2726),
.Y(n_3146)
);

INVx3_ASAP7_75t_L g3147 ( 
.A(n_2801),
.Y(n_3147)
);

INVx6_ASAP7_75t_L g3148 ( 
.A(n_2691),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2697),
.Y(n_3149)
);

INVx3_ASAP7_75t_L g3150 ( 
.A(n_2801),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2716),
.Y(n_3151)
);

AOI22xp33_ASAP7_75t_L g3152 ( 
.A1(n_3047),
.A2(n_2308),
.B1(n_2325),
.B2(n_2383),
.Y(n_3152)
);

INVx3_ASAP7_75t_L g3153 ( 
.A(n_2843),
.Y(n_3153)
);

OAI21x1_ASAP7_75t_L g3154 ( 
.A1(n_2926),
.A2(n_2517),
.B(n_2470),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2720),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2743),
.Y(n_3156)
);

AOI22xp33_ASAP7_75t_L g3157 ( 
.A1(n_3011),
.A2(n_2393),
.B1(n_2558),
.B2(n_2527),
.Y(n_3157)
);

BUFx6f_ASAP7_75t_L g3158 ( 
.A(n_2960),
.Y(n_3158)
);

AOI22xp33_ASAP7_75t_SL g3159 ( 
.A1(n_2787),
.A2(n_2568),
.B1(n_2619),
.B2(n_2573),
.Y(n_3159)
);

OAI22xp33_ASAP7_75t_L g3160 ( 
.A1(n_3017),
.A2(n_2630),
.B1(n_2210),
.B2(n_2211),
.Y(n_3160)
);

BUFx2_ASAP7_75t_L g3161 ( 
.A(n_2947),
.Y(n_3161)
);

OAI22xp33_ASAP7_75t_L g3162 ( 
.A1(n_2702),
.A2(n_2825),
.B1(n_2753),
.B2(n_2713),
.Y(n_3162)
);

CKINVDCx20_ASAP7_75t_R g3163 ( 
.A(n_2834),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2730),
.Y(n_3164)
);

INVx3_ASAP7_75t_L g3165 ( 
.A(n_2650),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2735),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2738),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2747),
.Y(n_3168)
);

OA21x2_ASAP7_75t_L g3169 ( 
.A1(n_2920),
.A2(n_2627),
.B(n_2179),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2751),
.Y(n_3170)
);

HB1xp67_ASAP7_75t_L g3171 ( 
.A(n_2679),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2770),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2762),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2765),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2778),
.Y(n_3175)
);

BUFx6f_ASAP7_75t_L g3176 ( 
.A(n_2966),
.Y(n_3176)
);

BUFx4f_ASAP7_75t_L g3177 ( 
.A(n_2825),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_2945),
.B(n_2205),
.Y(n_3178)
);

INVx1_ASAP7_75t_SL g3179 ( 
.A(n_2832),
.Y(n_3179)
);

BUFx2_ASAP7_75t_L g3180 ( 
.A(n_2947),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2818),
.Y(n_3181)
);

AOI22xp5_ASAP7_75t_L g3182 ( 
.A1(n_2950),
.A2(n_2177),
.B1(n_2228),
.B2(n_2217),
.Y(n_3182)
);

AOI21x1_ASAP7_75t_L g3183 ( 
.A1(n_3068),
.A2(n_2186),
.B(n_2169),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2893),
.B(n_2140),
.Y(n_3184)
);

CKINVDCx5p33_ASAP7_75t_R g3185 ( 
.A(n_2946),
.Y(n_3185)
);

INVx2_ASAP7_75t_SL g3186 ( 
.A(n_2757),
.Y(n_3186)
);

AOI22xp5_ASAP7_75t_L g3187 ( 
.A1(n_2950),
.A2(n_2230),
.B1(n_2197),
.B2(n_2143),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2820),
.Y(n_3188)
);

AOI22xp33_ASAP7_75t_L g3189 ( 
.A1(n_3018),
.A2(n_3046),
.B1(n_3020),
.B2(n_3050),
.Y(n_3189)
);

BUFx3_ASAP7_75t_L g3190 ( 
.A(n_2700),
.Y(n_3190)
);

OAI22xp33_ASAP7_75t_L g3191 ( 
.A1(n_2702),
.A2(n_2190),
.B1(n_2201),
.B2(n_2178),
.Y(n_3191)
);

BUFx2_ASAP7_75t_L g3192 ( 
.A(n_2947),
.Y(n_3192)
);

AND2x4_ASAP7_75t_L g3193 ( 
.A(n_2650),
.B(n_555),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2822),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2792),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2823),
.Y(n_3196)
);

INVx1_ASAP7_75t_SL g3197 ( 
.A(n_2832),
.Y(n_3197)
);

INVx4_ASAP7_75t_SL g3198 ( 
.A(n_2904),
.Y(n_3198)
);

OAI21xp5_ASAP7_75t_L g3199 ( 
.A1(n_3070),
.A2(n_2882),
.B(n_2876),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_2808),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2862),
.Y(n_3201)
);

AOI21x1_ASAP7_75t_L g3202 ( 
.A1(n_2684),
.A2(n_2337),
.B(n_2584),
.Y(n_3202)
);

CKINVDCx20_ASAP7_75t_R g3203 ( 
.A(n_2834),
.Y(n_3203)
);

OAI22xp5_ASAP7_75t_L g3204 ( 
.A1(n_2654),
.A2(n_2606),
.B1(n_558),
.B2(n_556),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2870),
.Y(n_3205)
);

BUFx4f_ASAP7_75t_L g3206 ( 
.A(n_2754),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2875),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_2812),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2841),
.Y(n_3209)
);

CKINVDCx5p33_ASAP7_75t_R g3210 ( 
.A(n_2757),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2833),
.Y(n_3211)
);

BUFx2_ASAP7_75t_R g3212 ( 
.A(n_2773),
.Y(n_3212)
);

CKINVDCx20_ASAP7_75t_R g3213 ( 
.A(n_2656),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2849),
.Y(n_3214)
);

BUFx2_ASAP7_75t_L g3215 ( 
.A(n_2889),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2855),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2860),
.Y(n_3217)
);

CKINVDCx11_ASAP7_75t_R g3218 ( 
.A(n_2699),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2766),
.Y(n_3219)
);

NAND2x1p5_ASAP7_75t_L g3220 ( 
.A(n_2704),
.B(n_863),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_2839),
.Y(n_3221)
);

INVxp67_ASAP7_75t_SL g3222 ( 
.A(n_2654),
.Y(n_3222)
);

OAI21x1_ASAP7_75t_L g3223 ( 
.A1(n_2879),
.A2(n_559),
.B(n_560),
.Y(n_3223)
);

BUFx2_ASAP7_75t_L g3224 ( 
.A(n_2691),
.Y(n_3224)
);

NAND2x1p5_ASAP7_75t_L g3225 ( 
.A(n_2719),
.B(n_562),
.Y(n_3225)
);

INVx4_ASAP7_75t_L g3226 ( 
.A(n_2749),
.Y(n_3226)
);

OAI22xp33_ASAP7_75t_L g3227 ( 
.A1(n_2702),
.A2(n_564),
.B1(n_562),
.B2(n_563),
.Y(n_3227)
);

BUFx6f_ASAP7_75t_L g3228 ( 
.A(n_2966),
.Y(n_3228)
);

AO21x1_ASAP7_75t_L g3229 ( 
.A1(n_3071),
.A2(n_563),
.B(n_565),
.Y(n_3229)
);

AOI22xp5_ASAP7_75t_L g3230 ( 
.A1(n_2828),
.A2(n_567),
.B1(n_565),
.B2(n_566),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2769),
.Y(n_3231)
);

OAI22xp5_ASAP7_75t_L g3232 ( 
.A1(n_2787),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.Y(n_3232)
);

INVx3_ASAP7_75t_L g3233 ( 
.A(n_2664),
.Y(n_3233)
);

HB1xp67_ASAP7_75t_L g3234 ( 
.A(n_2641),
.Y(n_3234)
);

AND2x4_ASAP7_75t_L g3235 ( 
.A(n_2664),
.B(n_569),
.Y(n_3235)
);

AND2x2_ASAP7_75t_L g3236 ( 
.A(n_2742),
.B(n_571),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2649),
.Y(n_3237)
);

HB1xp67_ASAP7_75t_L g3238 ( 
.A(n_2641),
.Y(n_3238)
);

BUFx2_ASAP7_75t_L g3239 ( 
.A(n_2943),
.Y(n_3239)
);

AND2x2_ASAP7_75t_L g3240 ( 
.A(n_2683),
.B(n_571),
.Y(n_3240)
);

BUFx6f_ASAP7_75t_L g3241 ( 
.A(n_2966),
.Y(n_3241)
);

OAI21x1_ASAP7_75t_L g3242 ( 
.A1(n_2879),
.A2(n_572),
.B(n_573),
.Y(n_3242)
);

BUFx3_ASAP7_75t_L g3243 ( 
.A(n_2784),
.Y(n_3243)
);

BUFx3_ASAP7_75t_L g3244 ( 
.A(n_2785),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2649),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2896),
.B(n_574),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2867),
.Y(n_3247)
);

NAND2x1p5_ASAP7_75t_L g3248 ( 
.A(n_2692),
.B(n_574),
.Y(n_3248)
);

HB1xp67_ASAP7_75t_L g3249 ( 
.A(n_3040),
.Y(n_3249)
);

OR2x2_ASAP7_75t_L g3250 ( 
.A(n_2790),
.B(n_575),
.Y(n_3250)
);

AO21x1_ASAP7_75t_L g3251 ( 
.A1(n_3071),
.A2(n_576),
.B(n_577),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_2771),
.Y(n_3252)
);

BUFx8_ASAP7_75t_L g3253 ( 
.A(n_2864),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2777),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_2683),
.B(n_576),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_2786),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_2797),
.Y(n_3257)
);

INVx2_ASAP7_75t_L g3258 ( 
.A(n_2803),
.Y(n_3258)
);

OAI22xp33_ASAP7_75t_L g3259 ( 
.A1(n_2713),
.A2(n_579),
.B1(n_577),
.B2(n_578),
.Y(n_3259)
);

BUFx4f_ASAP7_75t_L g3260 ( 
.A(n_2861),
.Y(n_3260)
);

HB1xp67_ASAP7_75t_L g3261 ( 
.A(n_3040),
.Y(n_3261)
);

AND2x4_ASAP7_75t_L g3262 ( 
.A(n_2676),
.B(n_579),
.Y(n_3262)
);

INVx6_ASAP7_75t_L g3263 ( 
.A(n_2878),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2930),
.Y(n_3264)
);

INVx2_ASAP7_75t_SL g3265 ( 
.A(n_2737),
.Y(n_3265)
);

OAI22xp5_ASAP7_75t_SL g3266 ( 
.A1(n_2656),
.A2(n_582),
.B1(n_580),
.B2(n_581),
.Y(n_3266)
);

OR2x6_ASAP7_75t_L g3267 ( 
.A(n_2707),
.B(n_580),
.Y(n_3267)
);

INVx2_ASAP7_75t_SL g3268 ( 
.A(n_2772),
.Y(n_3268)
);

INVx3_ASAP7_75t_L g3269 ( 
.A(n_2676),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_2968),
.B(n_581),
.Y(n_3270)
);

AOI22xp33_ASAP7_75t_L g3271 ( 
.A1(n_3046),
.A2(n_585),
.B1(n_583),
.B2(n_584),
.Y(n_3271)
);

OAI22xp5_ASAP7_75t_L g3272 ( 
.A1(n_2787),
.A2(n_587),
.B1(n_585),
.B2(n_586),
.Y(n_3272)
);

BUFx2_ASAP7_75t_L g3273 ( 
.A(n_2749),
.Y(n_3273)
);

AOI22xp33_ASAP7_75t_L g3274 ( 
.A1(n_3056),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_3274)
);

AOI22xp33_ASAP7_75t_SL g3275 ( 
.A1(n_2928),
.A2(n_593),
.B1(n_591),
.B2(n_592),
.Y(n_3275)
);

AOI22xp33_ASAP7_75t_SL g3276 ( 
.A1(n_2928),
.A2(n_593),
.B1(n_591),
.B2(n_592),
.Y(n_3276)
);

CKINVDCx11_ASAP7_75t_R g3277 ( 
.A(n_2739),
.Y(n_3277)
);

INVx3_ASAP7_75t_L g3278 ( 
.A(n_2710),
.Y(n_3278)
);

OR2x6_ASAP7_75t_L g3279 ( 
.A(n_2907),
.B(n_594),
.Y(n_3279)
);

INVx4_ASAP7_75t_L g3280 ( 
.A(n_2854),
.Y(n_3280)
);

AOI22xp33_ASAP7_75t_L g3281 ( 
.A1(n_2949),
.A2(n_2944),
.B1(n_2967),
.B2(n_2940),
.Y(n_3281)
);

BUFx6f_ASAP7_75t_L g3282 ( 
.A(n_2966),
.Y(n_3282)
);

OA21x2_ASAP7_75t_L g3283 ( 
.A1(n_2688),
.A2(n_594),
.B(n_595),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2723),
.Y(n_3284)
);

BUFx3_ASAP7_75t_L g3285 ( 
.A(n_2764),
.Y(n_3285)
);

OAI22xp5_ASAP7_75t_SL g3286 ( 
.A1(n_3035),
.A2(n_2829),
.B1(n_2868),
.B2(n_2866),
.Y(n_3286)
);

AOI22xp5_ASAP7_75t_L g3287 ( 
.A1(n_2828),
.A2(n_597),
.B1(n_595),
.B2(n_596),
.Y(n_3287)
);

AND2x4_ASAP7_75t_L g3288 ( 
.A(n_2710),
.B(n_2717),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_2881),
.Y(n_3289)
);

AND2x2_ASAP7_75t_L g3290 ( 
.A(n_3037),
.B(n_596),
.Y(n_3290)
);

INVx4_ASAP7_75t_L g3291 ( 
.A(n_2854),
.Y(n_3291)
);

AOI22xp33_ASAP7_75t_L g3292 ( 
.A1(n_2949),
.A2(n_600),
.B1(n_597),
.B2(n_598),
.Y(n_3292)
);

AOI22xp33_ASAP7_75t_L g3293 ( 
.A1(n_2949),
.A2(n_604),
.B1(n_601),
.B2(n_603),
.Y(n_3293)
);

BUFx12f_ASAP7_75t_L g3294 ( 
.A(n_2695),
.Y(n_3294)
);

OA21x2_ASAP7_75t_L g3295 ( 
.A1(n_2651),
.A2(n_605),
.B(n_606),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2725),
.Y(n_3296)
);

INVx6_ASAP7_75t_L g3297 ( 
.A(n_2898),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2804),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_2890),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_2892),
.Y(n_3300)
);

INVx3_ASAP7_75t_L g3301 ( 
.A(n_2717),
.Y(n_3301)
);

BUFx4f_ASAP7_75t_SL g3302 ( 
.A(n_2911),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2689),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2703),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2703),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3063),
.B(n_605),
.Y(n_3306)
);

BUFx3_ASAP7_75t_L g3307 ( 
.A(n_2779),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_3037),
.B(n_606),
.Y(n_3308)
);

AND2x2_ASAP7_75t_L g3309 ( 
.A(n_2783),
.B(n_607),
.Y(n_3309)
);

AND2x4_ASAP7_75t_L g3310 ( 
.A(n_2729),
.B(n_607),
.Y(n_3310)
);

AOI22xp33_ASAP7_75t_L g3311 ( 
.A1(n_2866),
.A2(n_611),
.B1(n_609),
.B2(n_610),
.Y(n_3311)
);

BUFx3_ASAP7_75t_L g3312 ( 
.A(n_2821),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2731),
.Y(n_3313)
);

AO21x2_ASAP7_75t_L g3314 ( 
.A1(n_2755),
.A2(n_860),
.B(n_613),
.Y(n_3314)
);

AO21x1_ASAP7_75t_L g3315 ( 
.A1(n_3065),
.A2(n_614),
.B(n_615),
.Y(n_3315)
);

INVx1_ASAP7_75t_SL g3316 ( 
.A(n_2865),
.Y(n_3316)
);

OAI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_2667),
.A2(n_617),
.B1(n_615),
.B2(n_616),
.Y(n_3317)
);

AOI22xp33_ASAP7_75t_L g3318 ( 
.A1(n_2868),
.A2(n_620),
.B1(n_617),
.B2(n_619),
.Y(n_3318)
);

OAI22xp5_ASAP7_75t_L g3319 ( 
.A1(n_2667),
.A2(n_621),
.B1(n_619),
.B2(n_620),
.Y(n_3319)
);

AOI22xp33_ASAP7_75t_L g3320 ( 
.A1(n_2915),
.A2(n_623),
.B1(n_621),
.B2(n_622),
.Y(n_3320)
);

AOI22xp33_ASAP7_75t_L g3321 ( 
.A1(n_2886),
.A2(n_624),
.B1(n_622),
.B2(n_623),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2731),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_2740),
.Y(n_3323)
);

INVx3_ASAP7_75t_L g3324 ( 
.A(n_2729),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_2740),
.Y(n_3325)
);

AND2x2_ASAP7_75t_L g3326 ( 
.A(n_2783),
.B(n_625),
.Y(n_3326)
);

AOI22xp33_ASAP7_75t_L g3327 ( 
.A1(n_2888),
.A2(n_628),
.B1(n_626),
.B2(n_627),
.Y(n_3327)
);

BUFx3_ASAP7_75t_L g3328 ( 
.A(n_2865),
.Y(n_3328)
);

HB1xp67_ASAP7_75t_L g3329 ( 
.A(n_2981),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_2972),
.B(n_626),
.Y(n_3330)
);

INVx3_ASAP7_75t_L g3331 ( 
.A(n_2767),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_2981),
.Y(n_3332)
);

BUFx2_ASAP7_75t_L g3333 ( 
.A(n_2750),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_2957),
.Y(n_3334)
);

OAI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_3070),
.A2(n_627),
.B(n_628),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_2957),
.Y(n_3336)
);

CKINVDCx6p67_ASAP7_75t_R g3337 ( 
.A(n_2931),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_2816),
.Y(n_3338)
);

BUFx2_ASAP7_75t_SL g3339 ( 
.A(n_2658),
.Y(n_3339)
);

AOI22xp33_ASAP7_75t_SL g3340 ( 
.A1(n_2928),
.A2(n_631),
.B1(n_629),
.B2(n_630),
.Y(n_3340)
);

AOI22xp33_ASAP7_75t_L g3341 ( 
.A1(n_3043),
.A2(n_633),
.B1(n_631),
.B2(n_632),
.Y(n_3341)
);

OR2x2_ASAP7_75t_L g3342 ( 
.A(n_2759),
.B(n_633),
.Y(n_3342)
);

OAI22xp5_ASAP7_75t_SL g3343 ( 
.A1(n_3035),
.A2(n_636),
.B1(n_634),
.B2(n_635),
.Y(n_3343)
);

OAI22xp33_ASAP7_75t_L g3344 ( 
.A1(n_3014),
.A2(n_637),
.B1(n_634),
.B2(n_636),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2817),
.Y(n_3345)
);

INVxp67_ASAP7_75t_SL g3346 ( 
.A(n_2794),
.Y(n_3346)
);

BUFx8_ASAP7_75t_L g3347 ( 
.A(n_2660),
.Y(n_3347)
);

INVx3_ASAP7_75t_L g3348 ( 
.A(n_3010),
.Y(n_3348)
);

INVxp33_ASAP7_75t_L g3349 ( 
.A(n_2978),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_2653),
.Y(n_3350)
);

BUFx2_ASAP7_75t_R g3351 ( 
.A(n_3016),
.Y(n_3351)
);

HB1xp67_ASAP7_75t_L g3352 ( 
.A(n_2760),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_2653),
.Y(n_3353)
);

NAND3xp33_ASAP7_75t_L g3354 ( 
.A(n_3036),
.B(n_637),
.C(n_638),
.Y(n_3354)
);

BUFx8_ASAP7_75t_L g3355 ( 
.A(n_2682),
.Y(n_3355)
);

OA21x2_ASAP7_75t_L g3356 ( 
.A1(n_2651),
.A2(n_638),
.B(n_640),
.Y(n_3356)
);

OR2x2_ASAP7_75t_L g3357 ( 
.A(n_3000),
.B(n_640),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_2696),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_SL g3359 ( 
.A1(n_3065),
.A2(n_643),
.B1(n_641),
.B2(n_642),
.Y(n_3359)
);

BUFx2_ASAP7_75t_L g3360 ( 
.A(n_2760),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_2819),
.Y(n_3361)
);

OAI22xp5_ASAP7_75t_L g3362 ( 
.A1(n_2674),
.A2(n_645),
.B1(n_642),
.B2(n_644),
.Y(n_3362)
);

OAI22xp5_ASAP7_75t_SL g3363 ( 
.A1(n_2829),
.A2(n_646),
.B1(n_644),
.B2(n_645),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_2827),
.Y(n_3364)
);

OAI21xp5_ASAP7_75t_SL g3365 ( 
.A1(n_3001),
.A2(n_647),
.B(n_648),
.Y(n_3365)
);

BUFx2_ASAP7_75t_R g3366 ( 
.A(n_3016),
.Y(n_3366)
);

BUFx4f_ASAP7_75t_SL g3367 ( 
.A(n_3053),
.Y(n_3367)
);

OAI21xp5_ASAP7_75t_L g3368 ( 
.A1(n_2882),
.A2(n_647),
.B(n_648),
.Y(n_3368)
);

BUFx12f_ASAP7_75t_L g3369 ( 
.A(n_2842),
.Y(n_3369)
);

AOI21x1_ASAP7_75t_L g3370 ( 
.A1(n_2980),
.A2(n_649),
.B(n_650),
.Y(n_3370)
);

OAI22xp5_ASAP7_75t_L g3371 ( 
.A1(n_2674),
.A2(n_652),
.B1(n_650),
.B2(n_651),
.Y(n_3371)
);

INVx3_ASAP7_75t_L g3372 ( 
.A(n_3010),
.Y(n_3372)
);

AOI22xp33_ASAP7_75t_L g3373 ( 
.A1(n_3043),
.A2(n_655),
.B1(n_653),
.B2(n_654),
.Y(n_3373)
);

AOI22xp33_ASAP7_75t_SL g3374 ( 
.A1(n_2873),
.A2(n_656),
.B1(n_654),
.B2(n_655),
.Y(n_3374)
);

HB1xp67_ASAP7_75t_L g3375 ( 
.A(n_2798),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_2696),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_2718),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3058),
.B(n_656),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_2718),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_2727),
.Y(n_3380)
);

BUFx2_ASAP7_75t_L g3381 ( 
.A(n_2798),
.Y(n_3381)
);

AND2x4_ASAP7_75t_L g3382 ( 
.A(n_3010),
.B(n_659),
.Y(n_3382)
);

OAI22xp33_ASAP7_75t_L g3383 ( 
.A1(n_2964),
.A2(n_662),
.B1(n_660),
.B2(n_661),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_2727),
.Y(n_3384)
);

AOI22xp33_ASAP7_75t_L g3385 ( 
.A1(n_2995),
.A2(n_664),
.B1(n_661),
.B2(n_663),
.Y(n_3385)
);

AOI22xp33_ASAP7_75t_L g3386 ( 
.A1(n_3002),
.A2(n_665),
.B1(n_663),
.B2(n_664),
.Y(n_3386)
);

HB1xp67_ASAP7_75t_L g3387 ( 
.A(n_2830),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_2922),
.B(n_665),
.Y(n_3388)
);

INVx6_ASAP7_75t_L g3389 ( 
.A(n_2694),
.Y(n_3389)
);

OR2x2_ASAP7_75t_L g3390 ( 
.A(n_2925),
.B(n_666),
.Y(n_3390)
);

AOI21x1_ASAP7_75t_L g3391 ( 
.A1(n_2948),
.A2(n_668),
.B(n_669),
.Y(n_3391)
);

CKINVDCx6p67_ASAP7_75t_R g3392 ( 
.A(n_2869),
.Y(n_3392)
);

AO21x2_ASAP7_75t_L g3393 ( 
.A1(n_2755),
.A2(n_854),
.B(n_669),
.Y(n_3393)
);

BUFx6f_ASAP7_75t_L g3394 ( 
.A(n_2640),
.Y(n_3394)
);

AOI22xp33_ASAP7_75t_SL g3395 ( 
.A1(n_2899),
.A2(n_672),
.B1(n_670),
.B2(n_671),
.Y(n_3395)
);

BUFx3_ASAP7_75t_L g3396 ( 
.A(n_2799),
.Y(n_3396)
);

CKINVDCx16_ASAP7_75t_R g3397 ( 
.A(n_2970),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_2744),
.Y(n_3398)
);

HB1xp67_ASAP7_75t_L g3399 ( 
.A(n_2830),
.Y(n_3399)
);

INVx1_ASAP7_75t_SL g3400 ( 
.A(n_2874),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_2744),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_2824),
.Y(n_3402)
);

AND2x2_ASAP7_75t_L g3403 ( 
.A(n_3058),
.B(n_2648),
.Y(n_3403)
);

BUFx3_ASAP7_75t_L g3404 ( 
.A(n_2800),
.Y(n_3404)
);

CKINVDCx11_ASAP7_75t_R g3405 ( 
.A(n_2983),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_2824),
.Y(n_3406)
);

AOI22xp33_ASAP7_75t_SL g3407 ( 
.A1(n_2964),
.A2(n_675),
.B1(n_673),
.B2(n_674),
.Y(n_3407)
);

INVx8_ASAP7_75t_L g3408 ( 
.A(n_2869),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_2748),
.Y(n_3409)
);

CKINVDCx5p33_ASAP7_75t_R g3410 ( 
.A(n_2858),
.Y(n_3410)
);

BUFx2_ASAP7_75t_L g3411 ( 
.A(n_2846),
.Y(n_3411)
);

HB1xp67_ASAP7_75t_L g3412 ( 
.A(n_2846),
.Y(n_3412)
);

CKINVDCx6p67_ASAP7_75t_R g3413 ( 
.A(n_2869),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_2748),
.Y(n_3414)
);

OA21x2_ASAP7_75t_L g3415 ( 
.A1(n_2948),
.A2(n_673),
.B(n_675),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_2761),
.Y(n_3416)
);

OAI21xp5_ASAP7_75t_L g3417 ( 
.A1(n_2807),
.A2(n_676),
.B(n_677),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_2761),
.Y(n_3418)
);

AND2x4_ASAP7_75t_L g3419 ( 
.A(n_3010),
.B(n_676),
.Y(n_3419)
);

AOI22xp33_ASAP7_75t_L g3420 ( 
.A1(n_2780),
.A2(n_680),
.B1(n_678),
.B2(n_679),
.Y(n_3420)
);

INVx4_ASAP7_75t_L g3421 ( 
.A(n_2907),
.Y(n_3421)
);

INVx4_ASAP7_75t_L g3422 ( 
.A(n_2904),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_2835),
.Y(n_3423)
);

INVx6_ASAP7_75t_L g3424 ( 
.A(n_2694),
.Y(n_3424)
);

OAI22xp5_ASAP7_75t_L g3425 ( 
.A1(n_2734),
.A2(n_682),
.B1(n_679),
.B2(n_681),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_2663),
.Y(n_3426)
);

BUFx2_ASAP7_75t_L g3427 ( 
.A(n_2856),
.Y(n_3427)
);

NAND2x1p5_ASAP7_75t_L g3428 ( 
.A(n_2733),
.B(n_854),
.Y(n_3428)
);

AOI22xp33_ASAP7_75t_L g3429 ( 
.A1(n_2780),
.A2(n_685),
.B1(n_683),
.B2(n_684),
.Y(n_3429)
);

INVx4_ASAP7_75t_L g3430 ( 
.A(n_2904),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_2663),
.Y(n_3431)
);

AOI22xp33_ASAP7_75t_SL g3432 ( 
.A1(n_2964),
.A2(n_687),
.B1(n_684),
.B2(n_686),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_2781),
.Y(n_3433)
);

INVx2_ASAP7_75t_SL g3434 ( 
.A(n_2655),
.Y(n_3434)
);

OAI21x1_ASAP7_75t_SL g3435 ( 
.A1(n_2852),
.A2(n_687),
.B(n_688),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_2781),
.Y(n_3436)
);

AOI22xp33_ASAP7_75t_L g3437 ( 
.A1(n_3029),
.A2(n_690),
.B1(n_688),
.B2(n_689),
.Y(n_3437)
);

INVx3_ASAP7_75t_L g3438 ( 
.A(n_2905),
.Y(n_3438)
);

INVx3_ASAP7_75t_L g3439 ( 
.A(n_2905),
.Y(n_3439)
);

BUFx3_ASAP7_75t_L g3440 ( 
.A(n_2813),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_2669),
.Y(n_3441)
);

BUFx4f_ASAP7_75t_L g3442 ( 
.A(n_2924),
.Y(n_3442)
);

AOI22xp33_ASAP7_75t_SL g3443 ( 
.A1(n_3061),
.A2(n_691),
.B1(n_689),
.B2(n_690),
.Y(n_3443)
);

HB1xp67_ASAP7_75t_L g3444 ( 
.A(n_2856),
.Y(n_3444)
);

INVx3_ASAP7_75t_L g3445 ( 
.A(n_2955),
.Y(n_3445)
);

OR2x6_ASAP7_75t_L g3446 ( 
.A(n_3060),
.B(n_693),
.Y(n_3446)
);

BUFx6f_ASAP7_75t_L g3447 ( 
.A(n_2640),
.Y(n_3447)
);

BUFx2_ASAP7_75t_L g3448 ( 
.A(n_3021),
.Y(n_3448)
);

CKINVDCx20_ASAP7_75t_R g3449 ( 
.A(n_2842),
.Y(n_3449)
);

INVx2_ASAP7_75t_SL g3450 ( 
.A(n_2655),
.Y(n_3450)
);

AO21x1_ASAP7_75t_L g3451 ( 
.A1(n_2796),
.A2(n_694),
.B(n_695),
.Y(n_3451)
);

BUFx2_ASAP7_75t_L g3452 ( 
.A(n_2733),
.Y(n_3452)
);

INVxp67_ASAP7_75t_L g3453 ( 
.A(n_2978),
.Y(n_3453)
);

BUFx2_ASAP7_75t_L g3454 ( 
.A(n_2942),
.Y(n_3454)
);

AOI22xp5_ASAP7_75t_L g3455 ( 
.A1(n_3069),
.A2(n_698),
.B1(n_696),
.B2(n_697),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_2669),
.Y(n_3456)
);

INVx3_ASAP7_75t_L g3457 ( 
.A(n_2955),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_2724),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_2724),
.Y(n_3459)
);

INVx2_ASAP7_75t_SL g3460 ( 
.A(n_2982),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_2768),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_2768),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_2810),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_2642),
.Y(n_3464)
);

BUFx2_ASAP7_75t_L g3465 ( 
.A(n_2877),
.Y(n_3465)
);

NOR2x1_ASAP7_75t_R g3466 ( 
.A(n_2746),
.B(n_697),
.Y(n_3466)
);

INVx2_ASAP7_75t_L g3467 ( 
.A(n_2859),
.Y(n_3467)
);

CKINVDCx11_ASAP7_75t_R g3468 ( 
.A(n_3076),
.Y(n_3468)
);

BUFx3_ASAP7_75t_L g3469 ( 
.A(n_2986),
.Y(n_3469)
);

AND2x2_ASAP7_75t_L g3470 ( 
.A(n_2709),
.B(n_699),
.Y(n_3470)
);

AOI22xp5_ASAP7_75t_L g3471 ( 
.A1(n_3069),
.A2(n_701),
.B1(n_699),
.B2(n_700),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_2665),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3033),
.B(n_700),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_2642),
.Y(n_3474)
);

OAI22xp33_ASAP7_75t_L g3475 ( 
.A1(n_3061),
.A2(n_705),
.B1(n_702),
.B2(n_703),
.Y(n_3475)
);

AND2x2_ASAP7_75t_L g3476 ( 
.A(n_2901),
.B(n_702),
.Y(n_3476)
);

OAI22x1_ASAP7_75t_L g3477 ( 
.A1(n_3001),
.A2(n_706),
.B1(n_703),
.B2(n_705),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_2884),
.B(n_707),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_2714),
.B(n_708),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3074),
.Y(n_3480)
);

INVx3_ASAP7_75t_L g3481 ( 
.A(n_2789),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3074),
.Y(n_3482)
);

BUFx10_ASAP7_75t_L g3483 ( 
.A(n_2746),
.Y(n_3483)
);

INVxp67_ASAP7_75t_L g3484 ( 
.A(n_2850),
.Y(n_3484)
);

CKINVDCx11_ASAP7_75t_R g3485 ( 
.A(n_3076),
.Y(n_3485)
);

AOI22xp33_ASAP7_75t_L g3486 ( 
.A1(n_3036),
.A2(n_711),
.B1(n_709),
.B2(n_710),
.Y(n_3486)
);

AND2x2_ASAP7_75t_L g3487 ( 
.A(n_2929),
.B(n_711),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_L g3488 ( 
.A1(n_3052),
.A2(n_714),
.B1(n_712),
.B2(n_713),
.Y(n_3488)
);

HB1xp67_ASAP7_75t_L g3489 ( 
.A(n_2925),
.Y(n_3489)
);

INVx3_ASAP7_75t_L g3490 ( 
.A(n_2789),
.Y(n_3490)
);

BUFx3_ASAP7_75t_L g3491 ( 
.A(n_2891),
.Y(n_3491)
);

AOI22xp33_ASAP7_75t_SL g3492 ( 
.A1(n_2796),
.A2(n_719),
.B1(n_715),
.B2(n_718),
.Y(n_3492)
);

AND2x2_ASAP7_75t_L g3493 ( 
.A(n_3038),
.B(n_719),
.Y(n_3493)
);

AND2x2_ASAP7_75t_L g3494 ( 
.A(n_3007),
.B(n_720),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_2706),
.Y(n_3495)
);

OAI22xp5_ASAP7_75t_L g3496 ( 
.A1(n_2871),
.A2(n_723),
.B1(n_721),
.B2(n_722),
.Y(n_3496)
);

BUFx10_ASAP7_75t_L g3497 ( 
.A(n_2752),
.Y(n_3497)
);

AND2x2_ASAP7_75t_L g3498 ( 
.A(n_2752),
.B(n_722),
.Y(n_3498)
);

OAI22xp5_ASAP7_75t_L g3499 ( 
.A1(n_3034),
.A2(n_725),
.B1(n_723),
.B2(n_724),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3264),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3100),
.Y(n_3501)
);

INVx2_ASAP7_75t_SL g3502 ( 
.A(n_3302),
.Y(n_3502)
);

OR2x6_ASAP7_75t_L g3503 ( 
.A(n_3408),
.B(n_2924),
.Y(n_3503)
);

CKINVDCx5p33_ASAP7_75t_R g3504 ( 
.A(n_3080),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3100),
.Y(n_3505)
);

NOR3xp33_ASAP7_75t_SL g3506 ( 
.A(n_3119),
.B(n_3185),
.C(n_3210),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3170),
.Y(n_3507)
);

OR2x6_ASAP7_75t_L g3508 ( 
.A(n_3408),
.B(n_2932),
.Y(n_3508)
);

OR2x2_ASAP7_75t_L g3509 ( 
.A(n_3109),
.B(n_2837),
.Y(n_3509)
);

INVxp67_ASAP7_75t_L g3510 ( 
.A(n_3352),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3079),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3290),
.B(n_3045),
.Y(n_3512)
);

AND2x2_ASAP7_75t_L g3513 ( 
.A(n_3308),
.B(n_3045),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_3102),
.Y(n_3514)
);

OR2x2_ASAP7_75t_L g3515 ( 
.A(n_3117),
.B(n_2938),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_R g3516 ( 
.A(n_3213),
.B(n_2789),
.Y(n_3516)
);

NOR2xp33_ASAP7_75t_R g3517 ( 
.A(n_3091),
.B(n_2789),
.Y(n_3517)
);

OAI22xp5_ASAP7_75t_L g3518 ( 
.A1(n_3279),
.A2(n_2657),
.B1(n_2872),
.B2(n_3034),
.Y(n_3518)
);

INVx2_ASAP7_75t_L g3519 ( 
.A(n_3103),
.Y(n_3519)
);

NOR2xp33_ASAP7_75t_R g3520 ( 
.A(n_3367),
.B(n_2789),
.Y(n_3520)
);

AND2x2_ASAP7_75t_L g3521 ( 
.A(n_3470),
.B(n_2976),
.Y(n_3521)
);

CKINVDCx6p67_ASAP7_75t_R g3522 ( 
.A(n_3088),
.Y(n_3522)
);

BUFx2_ASAP7_75t_L g3523 ( 
.A(n_3224),
.Y(n_3523)
);

HB1xp67_ASAP7_75t_L g3524 ( 
.A(n_3375),
.Y(n_3524)
);

NAND2xp33_ASAP7_75t_R g3525 ( 
.A(n_3267),
.B(n_2903),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3170),
.Y(n_3526)
);

NOR2xp33_ASAP7_75t_R g3527 ( 
.A(n_3080),
.B(n_2795),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3104),
.Y(n_3528)
);

HB1xp67_ASAP7_75t_L g3529 ( 
.A(n_3387),
.Y(n_3529)
);

NAND2xp33_ASAP7_75t_R g3530 ( 
.A(n_3267),
.B(n_2900),
.Y(n_3530)
);

BUFx3_ASAP7_75t_L g3531 ( 
.A(n_3082),
.Y(n_3531)
);

NAND2xp33_ASAP7_75t_R g3532 ( 
.A(n_3279),
.B(n_3446),
.Y(n_3532)
);

AND2x4_ASAP7_75t_L g3533 ( 
.A(n_3198),
.B(n_2836),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3105),
.Y(n_3534)
);

O2A1O1Ixp33_ASAP7_75t_L g3535 ( 
.A1(n_3160),
.A2(n_2814),
.B(n_2701),
.C(n_3066),
.Y(n_3535)
);

BUFx2_ASAP7_75t_L g3536 ( 
.A(n_3360),
.Y(n_3536)
);

CKINVDCx5p33_ASAP7_75t_R g3537 ( 
.A(n_3108),
.Y(n_3537)
);

AND2x2_ASAP7_75t_L g3538 ( 
.A(n_3236),
.B(n_3052),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3403),
.B(n_2847),
.Y(n_3539)
);

NOR2xp33_ASAP7_75t_R g3540 ( 
.A(n_3206),
.B(n_2906),
.Y(n_3540)
);

HB1xp67_ASAP7_75t_L g3541 ( 
.A(n_3399),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3173),
.Y(n_3542)
);

AND2x2_ASAP7_75t_L g3543 ( 
.A(n_3178),
.B(n_2919),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3173),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3129),
.B(n_2847),
.Y(n_3545)
);

OAI22xp5_ASAP7_75t_L g3546 ( 
.A1(n_3090),
.A2(n_2657),
.B1(n_2872),
.B2(n_2932),
.Y(n_3546)
);

AND2x2_ASAP7_75t_L g3547 ( 
.A(n_3096),
.B(n_2712),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_3309),
.B(n_2712),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_3326),
.B(n_3032),
.Y(n_3549)
);

CKINVDCx5p33_ASAP7_75t_R g3550 ( 
.A(n_3253),
.Y(n_3550)
);

AND2x2_ASAP7_75t_L g3551 ( 
.A(n_3113),
.B(n_3012),
.Y(n_3551)
);

AO31x2_ASAP7_75t_L g3552 ( 
.A1(n_3480),
.A2(n_2953),
.A3(n_2937),
.B(n_2959),
.Y(n_3552)
);

CKINVDCx5p33_ASAP7_75t_R g3553 ( 
.A(n_3253),
.Y(n_3553)
);

NAND3xp33_ASAP7_75t_SL g3554 ( 
.A(n_3349),
.B(n_3009),
.C(n_2814),
.Y(n_3554)
);

BUFx3_ASAP7_75t_L g3555 ( 
.A(n_3083),
.Y(n_3555)
);

OR2x2_ASAP7_75t_L g3556 ( 
.A(n_3249),
.B(n_2913),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3174),
.Y(n_3557)
);

INVx2_ASAP7_75t_L g3558 ( 
.A(n_3123),
.Y(n_3558)
);

AOI22xp33_ASAP7_75t_L g3559 ( 
.A1(n_3145),
.A2(n_3030),
.B1(n_2802),
.B2(n_3013),
.Y(n_3559)
);

INVx5_ASAP7_75t_SL g3560 ( 
.A(n_3392),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3240),
.B(n_3051),
.Y(n_3561)
);

BUFx3_ASAP7_75t_L g3562 ( 
.A(n_3190),
.Y(n_3562)
);

BUFx2_ASAP7_75t_L g3563 ( 
.A(n_3381),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3135),
.Y(n_3564)
);

AND2x2_ASAP7_75t_L g3565 ( 
.A(n_3255),
.B(n_2974),
.Y(n_3565)
);

CKINVDCx5p33_ASAP7_75t_R g3566 ( 
.A(n_3126),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3139),
.Y(n_3567)
);

NAND2xp33_ASAP7_75t_R g3568 ( 
.A(n_3446),
.B(n_2990),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3174),
.Y(n_3569)
);

NAND2xp33_ASAP7_75t_SL g3570 ( 
.A(n_3422),
.B(n_2852),
.Y(n_3570)
);

AOI22xp33_ASAP7_75t_L g3571 ( 
.A1(n_3162),
.A2(n_2802),
.B1(n_3077),
.B2(n_3054),
.Y(n_3571)
);

INVx2_ASAP7_75t_SL g3572 ( 
.A(n_3143),
.Y(n_3572)
);

AOI22xp33_ASAP7_75t_L g3573 ( 
.A1(n_3159),
.A2(n_3191),
.B1(n_3136),
.B2(n_3421),
.Y(n_3573)
);

OAI22xp33_ASAP7_75t_L g3574 ( 
.A1(n_3413),
.A2(n_3009),
.B1(n_3054),
.B2(n_3077),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3181),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3146),
.Y(n_3576)
);

BUFx6f_ASAP7_75t_L g3577 ( 
.A(n_3106),
.Y(n_3577)
);

OAI222xp33_ASAP7_75t_L g3578 ( 
.A1(n_3421),
.A2(n_3028),
.B1(n_2951),
.B2(n_2999),
.C1(n_3041),
.C2(n_2913),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3181),
.Y(n_3579)
);

AND2x2_ASAP7_75t_L g3580 ( 
.A(n_3378),
.B(n_2806),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3131),
.B(n_2935),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3188),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3188),
.Y(n_3583)
);

AND2x4_ASAP7_75t_L g3584 ( 
.A(n_3198),
.B(n_2836),
.Y(n_3584)
);

NOR2xp33_ASAP7_75t_L g3585 ( 
.A(n_3453),
.B(n_2858),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3196),
.Y(n_3586)
);

AND2x2_ASAP7_75t_L g3587 ( 
.A(n_3498),
.B(n_3330),
.Y(n_3587)
);

AND2x4_ASAP7_75t_L g3588 ( 
.A(n_3422),
.B(n_2914),
.Y(n_3588)
);

INVx11_ASAP7_75t_L g3589 ( 
.A(n_3347),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3196),
.Y(n_3590)
);

NAND3xp33_ASAP7_75t_L g3591 ( 
.A(n_3189),
.B(n_2937),
.C(n_2678),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3142),
.Y(n_3592)
);

INVx2_ASAP7_75t_L g3593 ( 
.A(n_3156),
.Y(n_3593)
);

CKINVDCx16_ASAP7_75t_R g3594 ( 
.A(n_3163),
.Y(n_3594)
);

INVx2_ASAP7_75t_L g3595 ( 
.A(n_3172),
.Y(n_3595)
);

INVx3_ASAP7_75t_L g3596 ( 
.A(n_3143),
.Y(n_3596)
);

INVx3_ASAP7_75t_SL g3597 ( 
.A(n_3263),
.Y(n_3597)
);

NOR3xp33_ASAP7_75t_SL g3598 ( 
.A(n_3410),
.B(n_2902),
.C(n_2885),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_3494),
.B(n_2806),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3479),
.B(n_2811),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3144),
.Y(n_3601)
);

OAI21xp5_ASAP7_75t_SL g3602 ( 
.A1(n_3365),
.A2(n_3085),
.B(n_3407),
.Y(n_3602)
);

INVxp33_ASAP7_75t_SL g3603 ( 
.A(n_3466),
.Y(n_3603)
);

OR2x6_ASAP7_75t_L g3604 ( 
.A(n_3186),
.B(n_3041),
.Y(n_3604)
);

AOI22xp33_ASAP7_75t_SL g3605 ( 
.A1(n_3442),
.A2(n_3430),
.B1(n_3329),
.B2(n_3110),
.Y(n_3605)
);

NOR2x1_ASAP7_75t_SL g3606 ( 
.A(n_3430),
.B(n_3073),
.Y(n_3606)
);

OR2x6_ASAP7_75t_L g3607 ( 
.A(n_3460),
.B(n_2711),
.Y(n_3607)
);

NOR2xp33_ASAP7_75t_R g3608 ( 
.A(n_3206),
.B(n_2670),
.Y(n_3608)
);

NOR3xp33_ASAP7_75t_SL g3609 ( 
.A(n_3094),
.B(n_2902),
.C(n_2885),
.Y(n_3609)
);

AND2x2_ASAP7_75t_L g3610 ( 
.A(n_3411),
.B(n_2811),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3149),
.Y(n_3611)
);

OR2x2_ASAP7_75t_L g3612 ( 
.A(n_3261),
.B(n_3234),
.Y(n_3612)
);

INVxp67_ASAP7_75t_L g3613 ( 
.A(n_3412),
.Y(n_3613)
);

OAI22xp5_ASAP7_75t_L g3614 ( 
.A1(n_3442),
.A2(n_2838),
.B1(n_3059),
.B2(n_2951),
.Y(n_3614)
);

AO31x2_ASAP7_75t_L g3615 ( 
.A1(n_3482),
.A2(n_2962),
.A3(n_2969),
.B(n_2959),
.Y(n_3615)
);

NAND2xp33_ASAP7_75t_R g3616 ( 
.A(n_3448),
.B(n_2990),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3151),
.Y(n_3617)
);

NOR2xp33_ASAP7_75t_R g3618 ( 
.A(n_3260),
.B(n_2670),
.Y(n_3618)
);

AND2x4_ASAP7_75t_L g3619 ( 
.A(n_3116),
.B(n_2914),
.Y(n_3619)
);

INVx3_ASAP7_75t_L g3620 ( 
.A(n_3148),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3155),
.Y(n_3621)
);

CKINVDCx5p33_ASAP7_75t_R g3622 ( 
.A(n_3140),
.Y(n_3622)
);

OR2x6_ASAP7_75t_L g3623 ( 
.A(n_3148),
.B(n_3028),
.Y(n_3623)
);

HB1xp67_ASAP7_75t_L g3624 ( 
.A(n_3444),
.Y(n_3624)
);

NOR2xp33_ASAP7_75t_R g3625 ( 
.A(n_3260),
.B(n_2954),
.Y(n_3625)
);

AOI22xp33_ASAP7_75t_L g3626 ( 
.A1(n_3118),
.A2(n_3199),
.B1(n_3120),
.B2(n_3078),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3164),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3166),
.B(n_3167),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3168),
.Y(n_3629)
);

AOI22xp33_ASAP7_75t_L g3630 ( 
.A1(n_3087),
.A2(n_3075),
.B1(n_2838),
.B2(n_3072),
.Y(n_3630)
);

OAI22xp5_ASAP7_75t_L g3631 ( 
.A1(n_3086),
.A2(n_3059),
.B1(n_2918),
.B2(n_2979),
.Y(n_3631)
);

OAI22xp5_ASAP7_75t_L g3632 ( 
.A1(n_3432),
.A2(n_3230),
.B1(n_3287),
.B2(n_3292),
.Y(n_3632)
);

NOR3xp33_ASAP7_75t_SL g3633 ( 
.A(n_3286),
.B(n_2975),
.C(n_2918),
.Y(n_3633)
);

BUFx2_ASAP7_75t_L g3634 ( 
.A(n_3427),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3194),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3201),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_3465),
.B(n_2975),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3205),
.B(n_2935),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3207),
.Y(n_3639)
);

OR2x2_ASAP7_75t_L g3640 ( 
.A(n_3238),
.B(n_2775),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3209),
.Y(n_3641)
);

BUFx10_ASAP7_75t_L g3642 ( 
.A(n_3263),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3214),
.Y(n_3643)
);

CKINVDCx5p33_ASAP7_75t_R g3644 ( 
.A(n_3218),
.Y(n_3644)
);

AND2x4_ASAP7_75t_L g3645 ( 
.A(n_3116),
.B(n_2908),
.Y(n_3645)
);

INVxp67_ASAP7_75t_L g3646 ( 
.A(n_3215),
.Y(n_3646)
);

CKINVDCx16_ASAP7_75t_R g3647 ( 
.A(n_3203),
.Y(n_3647)
);

NOR2xp33_ASAP7_75t_R g3648 ( 
.A(n_3468),
.B(n_2996),
.Y(n_3648)
);

AND2x4_ASAP7_75t_L g3649 ( 
.A(n_3134),
.B(n_2908),
.Y(n_3649)
);

NAND2xp33_ASAP7_75t_R g3650 ( 
.A(n_3273),
.B(n_724),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3175),
.Y(n_3651)
);

BUFx2_ASAP7_75t_L g3652 ( 
.A(n_3285),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3216),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_3195),
.Y(n_3654)
);

CKINVDCx5p33_ASAP7_75t_R g3655 ( 
.A(n_3277),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3217),
.B(n_2775),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3252),
.B(n_2788),
.Y(n_3657)
);

AO31x2_ASAP7_75t_L g3658 ( 
.A1(n_3482),
.A2(n_2962),
.A3(n_3008),
.B(n_2969),
.Y(n_3658)
);

CKINVDCx16_ASAP7_75t_R g3659 ( 
.A(n_3449),
.Y(n_3659)
);

BUFx2_ASAP7_75t_L g3660 ( 
.A(n_3452),
.Y(n_3660)
);

CKINVDCx16_ASAP7_75t_R g3661 ( 
.A(n_3101),
.Y(n_3661)
);

AO31x2_ASAP7_75t_L g3662 ( 
.A1(n_3426),
.A2(n_3008),
.A3(n_3027),
.B(n_3042),
.Y(n_3662)
);

OR2x6_ASAP7_75t_L g3663 ( 
.A(n_3297),
.B(n_3044),
.Y(n_3663)
);

CKINVDCx5p33_ASAP7_75t_R g3664 ( 
.A(n_3405),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3200),
.Y(n_3665)
);

CKINVDCx16_ASAP7_75t_R g3666 ( 
.A(n_3092),
.Y(n_3666)
);

AND2x2_ASAP7_75t_L g3667 ( 
.A(n_3473),
.B(n_2979),
.Y(n_3667)
);

O2A1O1Ixp33_ASAP7_75t_L g3668 ( 
.A1(n_3084),
.A2(n_3042),
.B(n_2844),
.C(n_2887),
.Y(n_3668)
);

AOI22xp33_ASAP7_75t_L g3669 ( 
.A1(n_3121),
.A2(n_3075),
.B1(n_3057),
.B2(n_3067),
.Y(n_3669)
);

OAI22xp5_ASAP7_75t_L g3670 ( 
.A1(n_3293),
.A2(n_2989),
.B1(n_3031),
.B2(n_3044),
.Y(n_3670)
);

AND2x4_ASAP7_75t_L g3671 ( 
.A(n_3134),
.B(n_2912),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3250),
.B(n_3031),
.Y(n_3672)
);

CKINVDCx20_ASAP7_75t_R g3673 ( 
.A(n_3485),
.Y(n_3673)
);

AND2x2_ASAP7_75t_L g3674 ( 
.A(n_3231),
.B(n_2991),
.Y(n_3674)
);

BUFx3_ASAP7_75t_L g3675 ( 
.A(n_3243),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3219),
.Y(n_3676)
);

OR2x6_ASAP7_75t_L g3677 ( 
.A(n_3297),
.B(n_3015),
.Y(n_3677)
);

AND2x2_ASAP7_75t_L g3678 ( 
.A(n_3256),
.B(n_726),
.Y(n_3678)
);

BUFx3_ASAP7_75t_L g3679 ( 
.A(n_3244),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3252),
.Y(n_3680)
);

NAND2xp33_ASAP7_75t_R g3681 ( 
.A(n_3161),
.B(n_727),
.Y(n_3681)
);

OR2x2_ASAP7_75t_L g3682 ( 
.A(n_3489),
.B(n_2788),
.Y(n_3682)
);

OAI22xp5_ASAP7_75t_L g3683 ( 
.A1(n_3455),
.A2(n_2722),
.B1(n_2708),
.B2(n_2715),
.Y(n_3683)
);

NAND2xp33_ASAP7_75t_R g3684 ( 
.A(n_3180),
.B(n_728),
.Y(n_3684)
);

CKINVDCx5p33_ASAP7_75t_R g3685 ( 
.A(n_3369),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3254),
.B(n_2793),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3254),
.B(n_2793),
.Y(n_3687)
);

AND2x2_ASAP7_75t_L g3688 ( 
.A(n_3257),
.B(n_728),
.Y(n_3688)
);

NOR2xp33_ASAP7_75t_R g3689 ( 
.A(n_3177),
.B(n_3347),
.Y(n_3689)
);

NAND2xp33_ASAP7_75t_R g3690 ( 
.A(n_3192),
.B(n_729),
.Y(n_3690)
);

CKINVDCx5p33_ASAP7_75t_R g3691 ( 
.A(n_3294),
.Y(n_3691)
);

NOR3xp33_ASAP7_75t_SL g3692 ( 
.A(n_3343),
.B(n_2715),
.C(n_2708),
.Y(n_3692)
);

OR2x2_ASAP7_75t_L g3693 ( 
.A(n_3258),
.B(n_3222),
.Y(n_3693)
);

OR2x6_ASAP7_75t_L g3694 ( 
.A(n_3280),
.B(n_3015),
.Y(n_3694)
);

BUFx10_ASAP7_75t_L g3695 ( 
.A(n_3434),
.Y(n_3695)
);

AND2x2_ASAP7_75t_L g3696 ( 
.A(n_3487),
.B(n_729),
.Y(n_3696)
);

AOI22xp33_ASAP7_75t_L g3697 ( 
.A1(n_3335),
.A2(n_3067),
.B1(n_2745),
.B2(n_2941),
.Y(n_3697)
);

OAI22xp5_ASAP7_75t_L g3698 ( 
.A1(n_3471),
.A2(n_2722),
.B1(n_2763),
.B2(n_3027),
.Y(n_3698)
);

AOI22xp33_ASAP7_75t_SL g3699 ( 
.A1(n_3110),
.A2(n_2880),
.B1(n_2895),
.B2(n_2831),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3281),
.B(n_2848),
.Y(n_3700)
);

OR2x6_ASAP7_75t_L g3701 ( 
.A(n_3280),
.B(n_3291),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3304),
.B(n_2848),
.Y(n_3702)
);

OAI21xp5_ASAP7_75t_L g3703 ( 
.A1(n_3097),
.A2(n_2763),
.B(n_2774),
.Y(n_3703)
);

OAI22xp5_ASAP7_75t_L g3704 ( 
.A1(n_3157),
.A2(n_2774),
.B1(n_2807),
.B2(n_3067),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3208),
.Y(n_3705)
);

AND2x4_ASAP7_75t_L g3706 ( 
.A(n_3288),
.B(n_2912),
.Y(n_3706)
);

CKINVDCx5p33_ASAP7_75t_R g3707 ( 
.A(n_3212),
.Y(n_3707)
);

A2O1A1Ixp33_ASAP7_75t_L g3708 ( 
.A1(n_3417),
.A2(n_3006),
.B(n_2998),
.C(n_2853),
.Y(n_3708)
);

NAND2xp33_ASAP7_75t_SL g3709 ( 
.A(n_3226),
.B(n_2857),
.Y(n_3709)
);

OR2x6_ASAP7_75t_L g3710 ( 
.A(n_3291),
.B(n_3019),
.Y(n_3710)
);

INVx2_ASAP7_75t_L g3711 ( 
.A(n_3211),
.Y(n_3711)
);

NAND2xp33_ASAP7_75t_R g3712 ( 
.A(n_3132),
.B(n_730),
.Y(n_3712)
);

OR2x2_ASAP7_75t_L g3713 ( 
.A(n_3141),
.B(n_2857),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3493),
.B(n_730),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3305),
.B(n_2909),
.Y(n_3715)
);

NOR2xp33_ASAP7_75t_R g3716 ( 
.A(n_3177),
.B(n_2897),
.Y(n_3716)
);

AND2x2_ASAP7_75t_L g3717 ( 
.A(n_3469),
.B(n_731),
.Y(n_3717)
);

INVx2_ASAP7_75t_L g3718 ( 
.A(n_3221),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3313),
.B(n_2909),
.Y(n_3719)
);

OR2x2_ASAP7_75t_L g3720 ( 
.A(n_3171),
.B(n_2988),
.Y(n_3720)
);

CKINVDCx16_ASAP7_75t_R g3721 ( 
.A(n_3092),
.Y(n_3721)
);

NAND2xp33_ASAP7_75t_R g3722 ( 
.A(n_3133),
.B(n_3331),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3322),
.B(n_2840),
.Y(n_3723)
);

OR2x6_ASAP7_75t_L g3724 ( 
.A(n_3339),
.B(n_3226),
.Y(n_3724)
);

AND2x2_ASAP7_75t_L g3725 ( 
.A(n_3476),
.B(n_731),
.Y(n_3725)
);

NOR2x1p5_ASAP7_75t_L g3726 ( 
.A(n_3328),
.B(n_2894),
.Y(n_3726)
);

AND2x2_ASAP7_75t_SL g3727 ( 
.A(n_3382),
.B(n_2897),
.Y(n_3727)
);

NAND2xp33_ASAP7_75t_R g3728 ( 
.A(n_3331),
.B(n_732),
.Y(n_3728)
);

OAI21xp33_ASAP7_75t_L g3729 ( 
.A1(n_3093),
.A2(n_3055),
.B(n_3022),
.Y(n_3729)
);

NOR2xp33_ASAP7_75t_R g3730 ( 
.A(n_3355),
.B(n_2646),
.Y(n_3730)
);

NOR3xp33_ASAP7_75t_SL g3731 ( 
.A(n_3266),
.B(n_2982),
.C(n_2994),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3193),
.B(n_732),
.Y(n_3732)
);

AND2x2_ASAP7_75t_L g3733 ( 
.A(n_3193),
.B(n_733),
.Y(n_3733)
);

OAI22xp5_ASAP7_75t_L g3734 ( 
.A1(n_3492),
.A2(n_2994),
.B1(n_2916),
.B2(n_2987),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3323),
.B(n_2840),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3325),
.B(n_2988),
.Y(n_3736)
);

AO31x2_ASAP7_75t_L g3737 ( 
.A1(n_3431),
.A2(n_2705),
.A3(n_2721),
.B(n_2985),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3289),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3246),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3235),
.Y(n_3740)
);

CKINVDCx5p33_ASAP7_75t_R g3741 ( 
.A(n_3337),
.Y(n_3741)
);

CKINVDCx5p33_ASAP7_75t_R g3742 ( 
.A(n_3351),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3235),
.Y(n_3743)
);

AOI22xp33_ASAP7_75t_L g3744 ( 
.A1(n_3137),
.A2(n_2758),
.B1(n_3026),
.B2(n_2756),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_3184),
.B(n_2993),
.Y(n_3745)
);

CKINVDCx5p33_ASAP7_75t_R g3746 ( 
.A(n_3366),
.Y(n_3746)
);

AO31x2_ASAP7_75t_L g3747 ( 
.A1(n_3441),
.A2(n_2705),
.A3(n_2721),
.B(n_2985),
.Y(n_3747)
);

OAI21xp5_ASAP7_75t_L g3748 ( 
.A1(n_3354),
.A2(n_2851),
.B(n_2809),
.Y(n_3748)
);

AND2x4_ASAP7_75t_L g3749 ( 
.A(n_3288),
.B(n_2987),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3262),
.Y(n_3750)
);

HB1xp67_ASAP7_75t_L g3751 ( 
.A(n_3484),
.Y(n_3751)
);

CKINVDCx5p33_ASAP7_75t_R g3752 ( 
.A(n_3355),
.Y(n_3752)
);

BUFx3_ASAP7_75t_L g3753 ( 
.A(n_3307),
.Y(n_3753)
);

HB1xp67_ASAP7_75t_L g3754 ( 
.A(n_3333),
.Y(n_3754)
);

BUFx2_ASAP7_75t_L g3755 ( 
.A(n_3396),
.Y(n_3755)
);

NAND2xp33_ASAP7_75t_SL g3756 ( 
.A(n_3147),
.B(n_2993),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3270),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3262),
.B(n_3310),
.Y(n_3758)
);

BUFx3_ASAP7_75t_L g3759 ( 
.A(n_3491),
.Y(n_3759)
);

NOR3xp33_ASAP7_75t_SL g3760 ( 
.A(n_3363),
.B(n_3003),
.C(n_2997),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3310),
.Y(n_3761)
);

AOI22xp33_ASAP7_75t_L g3762 ( 
.A1(n_3111),
.A2(n_3259),
.B1(n_3227),
.B2(n_3383),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_3478),
.B(n_733),
.Y(n_3763)
);

HB1xp67_ASAP7_75t_L g3764 ( 
.A(n_3454),
.Y(n_3764)
);

A2O1A1Ixp33_ASAP7_75t_L g3765 ( 
.A1(n_3368),
.A2(n_3353),
.B(n_3358),
.C(n_3350),
.Y(n_3765)
);

OR2x2_ASAP7_75t_L g3766 ( 
.A(n_3390),
.B(n_2997),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3223),
.Y(n_3767)
);

NAND2xp33_ASAP7_75t_R g3768 ( 
.A(n_3382),
.B(n_734),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3334),
.B(n_3003),
.Y(n_3769)
);

CKINVDCx5p33_ASAP7_75t_R g3770 ( 
.A(n_3397),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3336),
.B(n_3332),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_3357),
.B(n_734),
.Y(n_3772)
);

O2A1O1Ixp33_ASAP7_75t_SL g3773 ( 
.A1(n_3475),
.A2(n_2939),
.B(n_3073),
.C(n_3024),
.Y(n_3773)
);

AND2x2_ASAP7_75t_L g3774 ( 
.A(n_3404),
.B(n_735),
.Y(n_3774)
);

OR2x4_ASAP7_75t_L g3775 ( 
.A(n_3342),
.B(n_736),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3112),
.B(n_3005),
.Y(n_3776)
);

OAI22xp33_ASAP7_75t_L g3777 ( 
.A1(n_3428),
.A2(n_2693),
.B1(n_2916),
.B2(n_2961),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3440),
.B(n_738),
.Y(n_3778)
);

AND2x4_ASAP7_75t_L g3779 ( 
.A(n_3348),
.B(n_3372),
.Y(n_3779)
);

INVx2_ASAP7_75t_L g3780 ( 
.A(n_3242),
.Y(n_3780)
);

AND2x2_ASAP7_75t_L g3781 ( 
.A(n_3400),
.B(n_739),
.Y(n_3781)
);

CKINVDCx5p33_ASAP7_75t_R g3782 ( 
.A(n_3089),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_3346),
.B(n_3005),
.Y(n_3783)
);

NOR2xp33_ASAP7_75t_R g3784 ( 
.A(n_3450),
.B(n_2646),
.Y(n_3784)
);

OAI22xp5_ASAP7_75t_L g3785 ( 
.A1(n_3376),
.A2(n_2916),
.B1(n_2693),
.B2(n_2961),
.Y(n_3785)
);

AND2x2_ASAP7_75t_L g3786 ( 
.A(n_3312),
.B(n_740),
.Y(n_3786)
);

HB1xp67_ASAP7_75t_L g3787 ( 
.A(n_3377),
.Y(n_3787)
);

CKINVDCx14_ASAP7_75t_R g3788 ( 
.A(n_3239),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3081),
.Y(n_3789)
);

O2A1O1Ixp33_ASAP7_75t_L g3790 ( 
.A1(n_3232),
.A2(n_2934),
.B(n_2952),
.C(n_2933),
.Y(n_3790)
);

INVx2_ASAP7_75t_SL g3791 ( 
.A(n_3268),
.Y(n_3791)
);

CKINVDCx5p33_ASAP7_75t_R g3792 ( 
.A(n_3179),
.Y(n_3792)
);

NOR2x1p5_ASAP7_75t_L g3793 ( 
.A(n_3153),
.B(n_2646),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_3197),
.B(n_740),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_3379),
.B(n_3024),
.Y(n_3795)
);

INVxp67_ASAP7_75t_SL g3796 ( 
.A(n_3110),
.Y(n_3796)
);

CKINVDCx14_ASAP7_75t_R g3797 ( 
.A(n_3483),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3081),
.Y(n_3798)
);

CKINVDCx16_ASAP7_75t_R g3799 ( 
.A(n_3265),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3316),
.B(n_741),
.Y(n_3800)
);

HB1xp67_ASAP7_75t_L g3801 ( 
.A(n_3380),
.Y(n_3801)
);

NOR2xp33_ASAP7_75t_L g3802 ( 
.A(n_3107),
.B(n_741),
.Y(n_3802)
);

AND2x2_ASAP7_75t_L g3803 ( 
.A(n_3419),
.B(n_742),
.Y(n_3803)
);

AOI21xp33_ASAP7_75t_L g3804 ( 
.A1(n_3169),
.A2(n_2921),
.B(n_2756),
.Y(n_3804)
);

BUFx6f_ASAP7_75t_L g3805 ( 
.A(n_3106),
.Y(n_3805)
);

NAND3xp33_ASAP7_75t_SL g3806 ( 
.A(n_3220),
.B(n_742),
.C(n_743),
.Y(n_3806)
);

AND2x2_ASAP7_75t_L g3807 ( 
.A(n_3419),
.B(n_743),
.Y(n_3807)
);

NOR2xp33_ASAP7_75t_R g3808 ( 
.A(n_3153),
.B(n_2661),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3306),
.B(n_744),
.Y(n_3809)
);

NOR3xp33_ASAP7_75t_SL g3810 ( 
.A(n_3272),
.B(n_3025),
.C(n_2706),
.Y(n_3810)
);

HB1xp67_ASAP7_75t_L g3811 ( 
.A(n_3384),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3398),
.B(n_3025),
.Y(n_3812)
);

BUFx3_ASAP7_75t_L g3813 ( 
.A(n_3389),
.Y(n_3813)
);

AOI22xp33_ASAP7_75t_SL g3814 ( 
.A1(n_3110),
.A2(n_2933),
.B1(n_2952),
.B2(n_2934),
.Y(n_3814)
);

AND2x2_ASAP7_75t_L g3815 ( 
.A(n_3483),
.B(n_746),
.Y(n_3815)
);

NOR2xp33_ASAP7_75t_R g3816 ( 
.A(n_3110),
.B(n_2661),
.Y(n_3816)
);

INVx3_ASAP7_75t_L g3817 ( 
.A(n_3389),
.Y(n_3817)
);

BUFx6f_ASAP7_75t_L g3818 ( 
.A(n_3106),
.Y(n_3818)
);

NOR3xp33_ASAP7_75t_SL g3819 ( 
.A(n_3344),
.B(n_2971),
.C(n_2958),
.Y(n_3819)
);

CKINVDCx20_ASAP7_75t_R g3820 ( 
.A(n_3424),
.Y(n_3820)
);

BUFx3_ASAP7_75t_L g3821 ( 
.A(n_3424),
.Y(n_3821)
);

OR2x2_ASAP7_75t_SL g3822 ( 
.A(n_3295),
.B(n_2965),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3095),
.Y(n_3823)
);

BUFx6f_ASAP7_75t_L g3824 ( 
.A(n_3115),
.Y(n_3824)
);

AOI22xp33_ASAP7_75t_L g3825 ( 
.A1(n_3401),
.A2(n_2758),
.B1(n_2921),
.B2(n_2958),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3409),
.B(n_2971),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3095),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3098),
.Y(n_3828)
);

CKINVDCx5p33_ASAP7_75t_R g3829 ( 
.A(n_3497),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3098),
.Y(n_3830)
);

NAND3xp33_ASAP7_75t_SL g3831 ( 
.A(n_3225),
.B(n_3248),
.C(n_3275),
.Y(n_3831)
);

CKINVDCx16_ASAP7_75t_R g3832 ( 
.A(n_3497),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3099),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3099),
.Y(n_3834)
);

NAND2xp33_ASAP7_75t_R g3835 ( 
.A(n_3348),
.B(n_746),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3477),
.B(n_747),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3414),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3416),
.Y(n_3838)
);

CKINVDCx5p33_ASAP7_75t_R g3839 ( 
.A(n_3276),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3418),
.Y(n_3840)
);

NAND2xp33_ASAP7_75t_SL g3841 ( 
.A(n_3147),
.B(n_2977),
.Y(n_3841)
);

INVx1_ASAP7_75t_L g3842 ( 
.A(n_3388),
.Y(n_3842)
);

CKINVDCx5p33_ASAP7_75t_R g3843 ( 
.A(n_3340),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3372),
.B(n_747),
.Y(n_3844)
);

HB1xp67_ASAP7_75t_L g3845 ( 
.A(n_3165),
.Y(n_3845)
);

CKINVDCx16_ASAP7_75t_R g3846 ( 
.A(n_3115),
.Y(n_3846)
);

AND2x2_ASAP7_75t_SL g3847 ( 
.A(n_3150),
.B(n_2661),
.Y(n_3847)
);

BUFx6f_ASAP7_75t_L g3848 ( 
.A(n_3127),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3229),
.Y(n_3849)
);

BUFx6f_ASAP7_75t_SL g3850 ( 
.A(n_3127),
.Y(n_3850)
);

OR2x6_ASAP7_75t_L g3851 ( 
.A(n_3127),
.B(n_2662),
.Y(n_3851)
);

AOI22xp33_ASAP7_75t_L g3852 ( 
.A1(n_3496),
.A2(n_2984),
.B1(n_3062),
.B2(n_3039),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3251),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3152),
.B(n_748),
.Y(n_3854)
);

AOI22xp33_ASAP7_75t_L g3855 ( 
.A1(n_3435),
.A2(n_3064),
.B1(n_2939),
.B2(n_2673),
.Y(n_3855)
);

CKINVDCx5p33_ASAP7_75t_R g3856 ( 
.A(n_3158),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3341),
.B(n_2939),
.Y(n_3857)
);

CKINVDCx20_ASAP7_75t_R g3858 ( 
.A(n_3158),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3373),
.B(n_2939),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3182),
.B(n_2939),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3165),
.B(n_749),
.Y(n_3861)
);

HB1xp67_ASAP7_75t_L g3862 ( 
.A(n_3233),
.Y(n_3862)
);

CKINVDCx11_ASAP7_75t_R g3863 ( 
.A(n_3158),
.Y(n_3863)
);

OR2x6_ASAP7_75t_L g3864 ( 
.A(n_3176),
.B(n_2673),
.Y(n_3864)
);

INVx2_ASAP7_75t_SL g3865 ( 
.A(n_3176),
.Y(n_3865)
);

CKINVDCx5p33_ASAP7_75t_R g3866 ( 
.A(n_3176),
.Y(n_3866)
);

OR2x2_ASAP7_75t_L g3867 ( 
.A(n_3233),
.B(n_2736),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3451),
.Y(n_3868)
);

NOR2xp33_ASAP7_75t_R g3869 ( 
.A(n_3150),
.B(n_2736),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3269),
.B(n_3278),
.Y(n_3870)
);

CKINVDCx11_ASAP7_75t_R g3871 ( 
.A(n_3228),
.Y(n_3871)
);

AOI22xp5_ASAP7_75t_L g3872 ( 
.A1(n_3187),
.A2(n_2776),
.B1(n_2791),
.B2(n_2736),
.Y(n_3872)
);

NOR2xp33_ASAP7_75t_L g3873 ( 
.A(n_3128),
.B(n_749),
.Y(n_3873)
);

NOR2xp33_ASAP7_75t_R g3874 ( 
.A(n_3228),
.B(n_2776),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3269),
.B(n_2776),
.Y(n_3875)
);

NAND2xp33_ASAP7_75t_SL g3876 ( 
.A(n_3228),
.B(n_2992),
.Y(n_3876)
);

AND2x2_ASAP7_75t_L g3877 ( 
.A(n_3278),
.B(n_750),
.Y(n_3877)
);

NAND3xp33_ASAP7_75t_SL g3878 ( 
.A(n_3443),
.B(n_750),
.C(n_751),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3314),
.Y(n_3879)
);

NOR2xp33_ASAP7_75t_R g3880 ( 
.A(n_3241),
.B(n_2791),
.Y(n_3880)
);

AND2x2_ASAP7_75t_L g3881 ( 
.A(n_3587),
.B(n_3393),
.Y(n_3881)
);

OR2x2_ASAP7_75t_L g3882 ( 
.A(n_3693),
.B(n_3495),
.Y(n_3882)
);

HB1xp67_ASAP7_75t_L g3883 ( 
.A(n_3524),
.Y(n_3883)
);

AOI221xp5_ASAP7_75t_L g3884 ( 
.A1(n_3626),
.A2(n_3499),
.B1(n_3317),
.B2(n_3371),
.C(n_3362),
.Y(n_3884)
);

INVx2_ASAP7_75t_L g3885 ( 
.A(n_3511),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_3543),
.B(n_3393),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3501),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3505),
.Y(n_3888)
);

INVx2_ASAP7_75t_L g3889 ( 
.A(n_3514),
.Y(n_3889)
);

BUFx6f_ASAP7_75t_L g3890 ( 
.A(n_3863),
.Y(n_3890)
);

INVxp67_ASAP7_75t_L g3891 ( 
.A(n_3660),
.Y(n_3891)
);

AND2x2_ASAP7_75t_L g3892 ( 
.A(n_3551),
.B(n_3301),
.Y(n_3892)
);

AND2x2_ASAP7_75t_L g3893 ( 
.A(n_3561),
.B(n_3301),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3507),
.Y(n_3894)
);

BUFx3_ASAP7_75t_L g3895 ( 
.A(n_3531),
.Y(n_3895)
);

AND2x2_ASAP7_75t_SL g3896 ( 
.A(n_3727),
.B(n_3295),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3526),
.Y(n_3897)
);

HB1xp67_ASAP7_75t_L g3898 ( 
.A(n_3529),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3519),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3542),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3544),
.Y(n_3901)
);

AND2x2_ASAP7_75t_L g3902 ( 
.A(n_3512),
.B(n_3324),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3557),
.Y(n_3903)
);

BUFx3_ASAP7_75t_L g3904 ( 
.A(n_3752),
.Y(n_3904)
);

BUFx2_ASAP7_75t_L g3905 ( 
.A(n_3724),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3528),
.Y(n_3906)
);

INVx2_ASAP7_75t_L g3907 ( 
.A(n_3534),
.Y(n_3907)
);

NOR2xp33_ASAP7_75t_L g3908 ( 
.A(n_3603),
.B(n_3324),
.Y(n_3908)
);

INVx2_ASAP7_75t_L g3909 ( 
.A(n_3558),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3500),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3676),
.B(n_3464),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3592),
.Y(n_3912)
);

AND2x2_ASAP7_75t_L g3913 ( 
.A(n_3513),
.B(n_3438),
.Y(n_3913)
);

HB1xp67_ASAP7_75t_L g3914 ( 
.A(n_3541),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3601),
.Y(n_3915)
);

INVx3_ASAP7_75t_L g3916 ( 
.A(n_3588),
.Y(n_3916)
);

CKINVDCx6p67_ASAP7_75t_R g3917 ( 
.A(n_3597),
.Y(n_3917)
);

AO21x2_ASAP7_75t_L g3918 ( 
.A1(n_3804),
.A2(n_3462),
.B(n_3461),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3611),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3547),
.B(n_3438),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3617),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3621),
.Y(n_3922)
);

AND2x2_ASAP7_75t_L g3923 ( 
.A(n_3521),
.B(n_3439),
.Y(n_3923)
);

INVx8_ASAP7_75t_L g3924 ( 
.A(n_3724),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3627),
.Y(n_3925)
);

BUFx3_ASAP7_75t_L g3926 ( 
.A(n_3555),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3629),
.Y(n_3927)
);

BUFx3_ASAP7_75t_L g3928 ( 
.A(n_3562),
.Y(n_3928)
);

INVx2_ASAP7_75t_SL g3929 ( 
.A(n_3589),
.Y(n_3929)
);

AND2x2_ASAP7_75t_L g3930 ( 
.A(n_3549),
.B(n_3439),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3569),
.Y(n_3931)
);

AOI22xp33_ASAP7_75t_L g3932 ( 
.A1(n_3573),
.A2(n_3359),
.B1(n_3169),
.B2(n_3315),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3564),
.Y(n_3933)
);

BUFx3_ASAP7_75t_L g3934 ( 
.A(n_3675),
.Y(n_3934)
);

INVx3_ASAP7_75t_L g3935 ( 
.A(n_3588),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3536),
.B(n_3445),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3567),
.Y(n_3937)
);

INVx5_ASAP7_75t_L g3938 ( 
.A(n_3677),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3635),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_3576),
.Y(n_3940)
);

AND2x4_ASAP7_75t_L g3941 ( 
.A(n_3706),
.B(n_3458),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3636),
.B(n_3464),
.Y(n_3942)
);

AOI211xp5_ASAP7_75t_L g3943 ( 
.A1(n_3831),
.A2(n_3319),
.B(n_3425),
.C(n_3204),
.Y(n_3943)
);

AND2x2_ASAP7_75t_L g3944 ( 
.A(n_3563),
.B(n_3445),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3639),
.Y(n_3945)
);

AOI22xp33_ASAP7_75t_L g3946 ( 
.A1(n_3546),
.A2(n_3374),
.B1(n_3395),
.B2(n_3114),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3575),
.Y(n_3947)
);

HB1xp67_ASAP7_75t_L g3948 ( 
.A(n_3624),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_3593),
.Y(n_3949)
);

BUFx3_ASAP7_75t_L g3950 ( 
.A(n_3679),
.Y(n_3950)
);

INVx3_ASAP7_75t_L g3951 ( 
.A(n_3847),
.Y(n_3951)
);

OR2x2_ASAP7_75t_L g3952 ( 
.A(n_3612),
.B(n_3474),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3579),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3582),
.Y(n_3954)
);

OAI211xp5_ASAP7_75t_L g3955 ( 
.A1(n_3602),
.A2(n_3311),
.B(n_3318),
.C(n_3488),
.Y(n_3955)
);

AND2x2_ASAP7_75t_L g3956 ( 
.A(n_3634),
.B(n_3457),
.Y(n_3956)
);

INVx2_ASAP7_75t_L g3957 ( 
.A(n_3595),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3651),
.Y(n_3958)
);

AND2x2_ASAP7_75t_L g3959 ( 
.A(n_3758),
.B(n_3457),
.Y(n_3959)
);

AND2x4_ASAP7_75t_L g3960 ( 
.A(n_3706),
.B(n_3458),
.Y(n_3960)
);

AND2x4_ASAP7_75t_L g3961 ( 
.A(n_3789),
.B(n_3459),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3654),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3665),
.Y(n_3963)
);

NOR2xp33_ASAP7_75t_L g3964 ( 
.A(n_3799),
.B(n_3124),
.Y(n_3964)
);

INVxp67_ASAP7_75t_L g3965 ( 
.A(n_3523),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3641),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3705),
.Y(n_3967)
);

INVx2_ASAP7_75t_L g3968 ( 
.A(n_3711),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_3548),
.B(n_3674),
.Y(n_3969)
);

HB1xp67_ASAP7_75t_L g3970 ( 
.A(n_3510),
.Y(n_3970)
);

INVx2_ASAP7_75t_SL g3971 ( 
.A(n_3527),
.Y(n_3971)
);

AND2x2_ASAP7_75t_L g3972 ( 
.A(n_3538),
.B(n_3441),
.Y(n_3972)
);

INVx2_ASAP7_75t_L g3973 ( 
.A(n_3718),
.Y(n_3973)
);

AND2x2_ASAP7_75t_L g3974 ( 
.A(n_3764),
.B(n_3456),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3583),
.Y(n_3975)
);

INVx3_ASAP7_75t_L g3976 ( 
.A(n_3779),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3599),
.B(n_3600),
.Y(n_3977)
);

AND2x2_ASAP7_75t_L g3978 ( 
.A(n_3580),
.B(n_3456),
.Y(n_3978)
);

INVx3_ASAP7_75t_L g3979 ( 
.A(n_3779),
.Y(n_3979)
);

NOR2xp33_ASAP7_75t_L g3980 ( 
.A(n_3788),
.B(n_752),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3586),
.Y(n_3981)
);

AND2x2_ASAP7_75t_L g3982 ( 
.A(n_3610),
.B(n_3459),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3643),
.B(n_3474),
.Y(n_3983)
);

INVx4_ASAP7_75t_L g3984 ( 
.A(n_3503),
.Y(n_3984)
);

NOR2xp33_ASAP7_75t_L g3985 ( 
.A(n_3594),
.B(n_753),
.Y(n_3985)
);

BUFx3_ASAP7_75t_L g3986 ( 
.A(n_3820),
.Y(n_3986)
);

AND2x2_ASAP7_75t_L g3987 ( 
.A(n_3787),
.B(n_3461),
.Y(n_3987)
);

AND2x2_ASAP7_75t_L g3988 ( 
.A(n_3801),
.B(n_3462),
.Y(n_3988)
);

INVx4_ASAP7_75t_L g3989 ( 
.A(n_3503),
.Y(n_3989)
);

AND2x2_ASAP7_75t_L g3990 ( 
.A(n_3811),
.B(n_3754),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3590),
.Y(n_3991)
);

AND2x2_ASAP7_75t_L g3992 ( 
.A(n_3613),
.B(n_3284),
.Y(n_3992)
);

OR2x2_ASAP7_75t_L g3993 ( 
.A(n_3556),
.B(n_3237),
.Y(n_3993)
);

BUFx2_ASAP7_75t_L g3994 ( 
.A(n_3869),
.Y(n_3994)
);

INVx2_ASAP7_75t_L g3995 ( 
.A(n_3738),
.Y(n_3995)
);

INVx2_ASAP7_75t_L g3996 ( 
.A(n_3680),
.Y(n_3996)
);

AND2x2_ASAP7_75t_L g3997 ( 
.A(n_3751),
.B(n_3284),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3653),
.B(n_3296),
.Y(n_3998)
);

AND2x2_ASAP7_75t_L g3999 ( 
.A(n_3837),
.B(n_3296),
.Y(n_3999)
);

INVx2_ASAP7_75t_L g4000 ( 
.A(n_3798),
.Y(n_4000)
);

INVx2_ASAP7_75t_L g4001 ( 
.A(n_3823),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3827),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3828),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3838),
.B(n_3241),
.Y(n_4004)
);

OR2x6_ASAP7_75t_L g4005 ( 
.A(n_3508),
.B(n_3241),
.Y(n_4005)
);

BUFx2_ASAP7_75t_L g4006 ( 
.A(n_3858),
.Y(n_4006)
);

BUFx3_ASAP7_75t_L g4007 ( 
.A(n_3753),
.Y(n_4007)
);

AND2x2_ASAP7_75t_L g4008 ( 
.A(n_3840),
.B(n_3509),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3830),
.Y(n_4009)
);

OR2x2_ASAP7_75t_L g4010 ( 
.A(n_3515),
.B(n_3237),
.Y(n_4010)
);

BUFx3_ASAP7_75t_L g4011 ( 
.A(n_3759),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3628),
.Y(n_4012)
);

AOI211xp5_ASAP7_75t_L g4013 ( 
.A1(n_3518),
.A2(n_3554),
.B(n_3574),
.C(n_3632),
.Y(n_4013)
);

INVx3_ASAP7_75t_L g4014 ( 
.A(n_3645),
.Y(n_4014)
);

HB1xp67_ASAP7_75t_L g4015 ( 
.A(n_3646),
.Y(n_4015)
);

AND2x2_ASAP7_75t_L g4016 ( 
.A(n_3652),
.B(n_3282),
.Y(n_4016)
);

OAI221xp5_ASAP7_75t_L g4017 ( 
.A1(n_3532),
.A2(n_3486),
.B1(n_3420),
.B2(n_3429),
.C(n_3321),
.Y(n_4017)
);

INVx2_ASAP7_75t_L g4018 ( 
.A(n_3833),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3755),
.B(n_3282),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3846),
.B(n_3282),
.Y(n_4020)
);

AND2x2_ASAP7_75t_L g4021 ( 
.A(n_3637),
.B(n_3717),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3834),
.Y(n_4022)
);

AOI22xp5_ASAP7_75t_L g4023 ( 
.A1(n_3768),
.A2(n_3327),
.B1(n_3274),
.B2(n_3271),
.Y(n_4023)
);

AND2x2_ASAP7_75t_L g4024 ( 
.A(n_3725),
.B(n_3183),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_3539),
.B(n_3672),
.Y(n_4025)
);

INVx2_ASAP7_75t_L g4026 ( 
.A(n_3771),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3723),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3735),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3657),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_3842),
.B(n_3739),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_3732),
.B(n_3356),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3686),
.Y(n_4032)
);

BUFx3_ASAP7_75t_L g4033 ( 
.A(n_3642),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3757),
.B(n_3320),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3640),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3733),
.B(n_3356),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3667),
.B(n_3385),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_L g4038 ( 
.A(n_3545),
.B(n_3386),
.Y(n_4038)
);

INVx2_ASAP7_75t_L g4039 ( 
.A(n_3867),
.Y(n_4039)
);

INVx2_ASAP7_75t_L g4040 ( 
.A(n_3870),
.Y(n_4040)
);

AND2x2_ASAP7_75t_L g4041 ( 
.A(n_3774),
.B(n_3415),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_3581),
.B(n_3437),
.Y(n_4042)
);

BUFx2_ASAP7_75t_SL g4043 ( 
.A(n_3502),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3682),
.Y(n_4044)
);

HB1xp67_ASAP7_75t_L g4045 ( 
.A(n_3845),
.Y(n_4045)
);

INVx2_ASAP7_75t_L g4046 ( 
.A(n_3577),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3720),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3713),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_3778),
.B(n_3415),
.Y(n_4049)
);

NOR2xp33_ASAP7_75t_L g4050 ( 
.A(n_3647),
.B(n_755),
.Y(n_4050)
);

INVxp67_ASAP7_75t_SL g4051 ( 
.A(n_3862),
.Y(n_4051)
);

AOI22xp5_ASAP7_75t_L g4052 ( 
.A1(n_3839),
.A2(n_3472),
.B1(n_3345),
.B2(n_3361),
.Y(n_4052)
);

AND2x4_ASAP7_75t_L g4053 ( 
.A(n_3796),
.B(n_3481),
.Y(n_4053)
);

AND2x2_ASAP7_75t_L g4054 ( 
.A(n_3803),
.B(n_3338),
.Y(n_4054)
);

OR2x2_ASAP7_75t_L g4055 ( 
.A(n_3766),
.B(n_3656),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3687),
.Y(n_4056)
);

AND2x2_ASAP7_75t_L g4057 ( 
.A(n_3807),
.B(n_3338),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_3740),
.B(n_3345),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_3743),
.B(n_3361),
.Y(n_4059)
);

INVx2_ASAP7_75t_L g4060 ( 
.A(n_3577),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3577),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3638),
.B(n_3298),
.Y(n_4062)
);

HB1xp67_ASAP7_75t_L g4063 ( 
.A(n_3750),
.Y(n_4063)
);

AND2x4_ASAP7_75t_L g4064 ( 
.A(n_3645),
.B(n_3481),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3805),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_3761),
.B(n_3364),
.Y(n_4066)
);

AND2x2_ASAP7_75t_L g4067 ( 
.A(n_3786),
.B(n_3364),
.Y(n_4067)
);

AND2x4_ASAP7_75t_SL g4068 ( 
.A(n_3508),
.B(n_3394),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3736),
.Y(n_4069)
);

OR2x2_ASAP7_75t_L g4070 ( 
.A(n_3791),
.B(n_3245),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3702),
.Y(n_4071)
);

INVxp67_ASAP7_75t_L g4072 ( 
.A(n_3530),
.Y(n_4072)
);

BUFx3_ASAP7_75t_L g4073 ( 
.A(n_3504),
.Y(n_4073)
);

INVxp67_ASAP7_75t_L g4074 ( 
.A(n_3525),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3609),
.B(n_3678),
.Y(n_4075)
);

AND2x2_ASAP7_75t_L g4076 ( 
.A(n_3749),
.B(n_3423),
.Y(n_4076)
);

BUFx2_ASAP7_75t_L g4077 ( 
.A(n_3730),
.Y(n_4077)
);

AND2x2_ASAP7_75t_L g4078 ( 
.A(n_3749),
.B(n_3423),
.Y(n_4078)
);

INVx2_ASAP7_75t_L g4079 ( 
.A(n_3805),
.Y(n_4079)
);

OR2x2_ASAP7_75t_L g4080 ( 
.A(n_3715),
.B(n_3245),
.Y(n_4080)
);

BUFx2_ASAP7_75t_L g4081 ( 
.A(n_3856),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_3719),
.Y(n_4082)
);

AND2x4_ASAP7_75t_L g4083 ( 
.A(n_3649),
.B(n_3490),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_3763),
.B(n_3298),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_3805),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3795),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_3688),
.B(n_3247),
.Y(n_4087)
);

OR2x2_ASAP7_75t_L g4088 ( 
.A(n_3769),
.B(n_3433),
.Y(n_4088)
);

BUFx6f_ASAP7_75t_L g4089 ( 
.A(n_3871),
.Y(n_4089)
);

AND2x2_ASAP7_75t_L g4090 ( 
.A(n_3794),
.B(n_3303),
.Y(n_4090)
);

HB1xp67_ASAP7_75t_L g4091 ( 
.A(n_3649),
.Y(n_4091)
);

NOR2x1_ASAP7_75t_L g4092 ( 
.A(n_3701),
.B(n_3490),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_3818),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3615),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_3800),
.B(n_3299),
.Y(n_4095)
);

NOR2xp33_ASAP7_75t_L g4096 ( 
.A(n_3792),
.B(n_755),
.Y(n_4096)
);

INVx2_ASAP7_75t_L g4097 ( 
.A(n_3818),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_3615),
.Y(n_4098)
);

INVx2_ASAP7_75t_L g4099 ( 
.A(n_3818),
.Y(n_4099)
);

HB1xp67_ASAP7_75t_L g4100 ( 
.A(n_3671),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3615),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3658),
.Y(n_4102)
);

HB1xp67_ASAP7_75t_L g4103 ( 
.A(n_3671),
.Y(n_4103)
);

AND2x4_ASAP7_75t_L g4104 ( 
.A(n_3533),
.B(n_3247),
.Y(n_4104)
);

INVx2_ASAP7_75t_L g4105 ( 
.A(n_3824),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_3658),
.Y(n_4106)
);

NOR2x1_ASAP7_75t_L g4107 ( 
.A(n_3701),
.B(n_3300),
.Y(n_4107)
);

INVx1_ASAP7_75t_SL g4108 ( 
.A(n_3689),
.Y(n_4108)
);

BUFx2_ASAP7_75t_L g4109 ( 
.A(n_3866),
.Y(n_4109)
);

NOR2xp33_ASAP7_75t_L g4110 ( 
.A(n_3782),
.B(n_756),
.Y(n_4110)
);

OR2x2_ASAP7_75t_L g4111 ( 
.A(n_3812),
.B(n_3436),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_3824),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_3658),
.Y(n_4113)
);

AOI22xp33_ASAP7_75t_L g4114 ( 
.A1(n_3878),
.A2(n_3463),
.B1(n_3467),
.B2(n_3122),
.Y(n_4114)
);

OR2x2_ASAP7_75t_L g4115 ( 
.A(n_3783),
.B(n_3402),
.Y(n_4115)
);

BUFx2_ASAP7_75t_L g4116 ( 
.A(n_3874),
.Y(n_4116)
);

INVx4_ASAP7_75t_L g4117 ( 
.A(n_3694),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3662),
.Y(n_4118)
);

BUFx2_ASAP7_75t_L g4119 ( 
.A(n_3880),
.Y(n_4119)
);

AND2x2_ASAP7_75t_L g4120 ( 
.A(n_3696),
.B(n_3138),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_3703),
.B(n_3130),
.Y(n_4121)
);

AND2x2_ASAP7_75t_L g4122 ( 
.A(n_3714),
.B(n_3122),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_3772),
.B(n_3394),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_3781),
.B(n_3394),
.Y(n_4124)
);

INVx2_ASAP7_75t_L g4125 ( 
.A(n_3824),
.Y(n_4125)
);

BUFx2_ASAP7_75t_L g4126 ( 
.A(n_3784),
.Y(n_4126)
);

OR2x2_ASAP7_75t_L g4127 ( 
.A(n_3745),
.B(n_3406),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3848),
.Y(n_4128)
);

INVx1_ASAP7_75t_SL g4129 ( 
.A(n_3648),
.Y(n_4129)
);

HB1xp67_ASAP7_75t_L g4130 ( 
.A(n_3619),
.Y(n_4130)
);

INVxp67_ASAP7_75t_L g4131 ( 
.A(n_3895),
.Y(n_4131)
);

AND2x2_ASAP7_75t_SL g4132 ( 
.A(n_4117),
.B(n_3666),
.Y(n_4132)
);

AND2x2_ASAP7_75t_L g4133 ( 
.A(n_3977),
.B(n_3860),
.Y(n_4133)
);

BUFx2_ASAP7_75t_L g4134 ( 
.A(n_3994),
.Y(n_4134)
);

INVx3_ASAP7_75t_L g4135 ( 
.A(n_4117),
.Y(n_4135)
);

AND2x2_ASAP7_75t_L g4136 ( 
.A(n_4021),
.B(n_3826),
.Y(n_4136)
);

OR2x2_ASAP7_75t_L g4137 ( 
.A(n_3883),
.B(n_3898),
.Y(n_4137)
);

OR2x2_ASAP7_75t_L g4138 ( 
.A(n_3914),
.B(n_3776),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_3910),
.Y(n_4139)
);

AND2x2_ASAP7_75t_L g4140 ( 
.A(n_3990),
.B(n_3700),
.Y(n_4140)
);

INVx2_ASAP7_75t_L g4141 ( 
.A(n_3885),
.Y(n_4141)
);

AND2x2_ASAP7_75t_L g4142 ( 
.A(n_3972),
.B(n_3565),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_3881),
.B(n_3704),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_3912),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_4012),
.B(n_3868),
.Y(n_4145)
);

AND2x4_ASAP7_75t_L g4146 ( 
.A(n_4014),
.B(n_3879),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_4025),
.B(n_3662),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_4026),
.B(n_3662),
.Y(n_4148)
);

HB1xp67_ASAP7_75t_L g4149 ( 
.A(n_3948),
.Y(n_4149)
);

AND2x4_ASAP7_75t_L g4150 ( 
.A(n_4014),
.B(n_3533),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_3886),
.B(n_3571),
.Y(n_4151)
);

INVx2_ASAP7_75t_L g4152 ( 
.A(n_3889),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_3899),
.Y(n_4153)
);

AND2x2_ASAP7_75t_L g4154 ( 
.A(n_4040),
.B(n_3619),
.Y(n_4154)
);

AND2x2_ASAP7_75t_L g4155 ( 
.A(n_3893),
.B(n_3552),
.Y(n_4155)
);

AND2x2_ASAP7_75t_L g4156 ( 
.A(n_4091),
.B(n_3552),
.Y(n_4156)
);

HB1xp67_ASAP7_75t_L g4157 ( 
.A(n_4045),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_3906),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_4047),
.B(n_3631),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_4048),
.B(n_3683),
.Y(n_4160)
);

AND2x2_ASAP7_75t_L g4161 ( 
.A(n_4100),
.B(n_4103),
.Y(n_4161)
);

HB1xp67_ASAP7_75t_L g4162 ( 
.A(n_4130),
.Y(n_4162)
);

NAND2x1_ASAP7_75t_SL g4163 ( 
.A(n_3984),
.B(n_3585),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_4035),
.B(n_3836),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_3915),
.Y(n_4165)
);

AND2x2_ASAP7_75t_L g4166 ( 
.A(n_3969),
.B(n_3552),
.Y(n_4166)
);

AND2x2_ASAP7_75t_L g4167 ( 
.A(n_4008),
.B(n_3872),
.Y(n_4167)
);

AND2x2_ASAP7_75t_L g4168 ( 
.A(n_3892),
.B(n_3606),
.Y(n_4168)
);

NOR2xp33_ASAP7_75t_L g4169 ( 
.A(n_3926),
.B(n_3661),
.Y(n_4169)
);

OR2x2_ASAP7_75t_L g4170 ( 
.A(n_4055),
.B(n_3721),
.Y(n_4170)
);

INVxp67_ASAP7_75t_R g4171 ( 
.A(n_3917),
.Y(n_4171)
);

HB1xp67_ASAP7_75t_L g4172 ( 
.A(n_3970),
.Y(n_4172)
);

AND2x4_ASAP7_75t_L g4173 ( 
.A(n_4104),
.B(n_3584),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_3887),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_4044),
.B(n_3997),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_3919),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_L g4177 ( 
.A(n_3995),
.B(n_3978),
.Y(n_4177)
);

AND2x4_ASAP7_75t_L g4178 ( 
.A(n_4104),
.B(n_3584),
.Y(n_4178)
);

OR2x2_ASAP7_75t_L g4179 ( 
.A(n_3952),
.B(n_3560),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_3921),
.Y(n_4180)
);

OR2x2_ASAP7_75t_L g4181 ( 
.A(n_3882),
.B(n_3560),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_3922),
.Y(n_4182)
);

AOI22xp33_ASAP7_75t_L g4183 ( 
.A1(n_3946),
.A2(n_3570),
.B1(n_3614),
.B2(n_3762),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_3925),
.Y(n_4184)
);

OR2x2_ASAP7_75t_L g4185 ( 
.A(n_3993),
.B(n_3822),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3927),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_3930),
.B(n_3607),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_3939),
.Y(n_4188)
);

INVx2_ASAP7_75t_L g4189 ( 
.A(n_3907),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_3945),
.Y(n_4190)
);

INVx2_ASAP7_75t_L g4191 ( 
.A(n_3909),
.Y(n_4191)
);

AOI221xp5_ASAP7_75t_L g4192 ( 
.A1(n_4013),
.A2(n_3802),
.B1(n_3535),
.B2(n_3873),
.C(n_3806),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_3974),
.B(n_3692),
.Y(n_4193)
);

AND2x2_ASAP7_75t_L g4194 ( 
.A(n_4090),
.B(n_3607),
.Y(n_4194)
);

AOI211xp5_ASAP7_75t_L g4195 ( 
.A1(n_3980),
.A2(n_3608),
.B(n_3618),
.C(n_3716),
.Y(n_4195)
);

HB1xp67_ASAP7_75t_L g4196 ( 
.A(n_3891),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_4095),
.B(n_3854),
.Y(n_4197)
);

AOI22xp33_ASAP7_75t_L g4198 ( 
.A1(n_3896),
.A2(n_3559),
.B1(n_3670),
.B2(n_3698),
.Y(n_4198)
);

AND2x4_ASAP7_75t_L g4199 ( 
.A(n_3916),
.B(n_3813),
.Y(n_4199)
);

NOR2xp33_ASAP7_75t_L g4200 ( 
.A(n_3928),
.B(n_3659),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_3992),
.B(n_3849),
.Y(n_4201)
);

AND2x2_ASAP7_75t_L g4202 ( 
.A(n_4054),
.B(n_3821),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_3966),
.Y(n_4203)
);

AND2x2_ASAP7_75t_L g4204 ( 
.A(n_4057),
.B(n_3815),
.Y(n_4204)
);

AND2x2_ASAP7_75t_L g4205 ( 
.A(n_3902),
.B(n_3832),
.Y(n_4205)
);

INVx2_ASAP7_75t_L g4206 ( 
.A(n_3933),
.Y(n_4206)
);

INVx3_ASAP7_75t_L g4207 ( 
.A(n_3924),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_4084),
.B(n_3853),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_3887),
.Y(n_4209)
);

AND2x2_ASAP7_75t_L g4210 ( 
.A(n_3923),
.B(n_3797),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_L g4211 ( 
.A(n_4000),
.B(n_3765),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_3888),
.Y(n_4212)
);

INVx2_ASAP7_75t_L g4213 ( 
.A(n_3937),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_3888),
.Y(n_4214)
);

OR2x2_ASAP7_75t_L g4215 ( 
.A(n_4010),
.B(n_3737),
.Y(n_4215)
);

INVx2_ASAP7_75t_L g4216 ( 
.A(n_3940),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_4001),
.B(n_3630),
.Y(n_4217)
);

AND2x2_ASAP7_75t_L g4218 ( 
.A(n_3959),
.B(n_3865),
.Y(n_4218)
);

AND2x4_ASAP7_75t_SL g4219 ( 
.A(n_3890),
.B(n_3677),
.Y(n_4219)
);

INVxp67_ASAP7_75t_SL g4220 ( 
.A(n_4051),
.Y(n_4220)
);

INVxp67_ASAP7_75t_SL g4221 ( 
.A(n_4107),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_4018),
.B(n_3598),
.Y(n_4222)
);

NAND4xp25_ASAP7_75t_L g4223 ( 
.A(n_3943),
.B(n_3650),
.C(n_3684),
.D(n_3681),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_L g4224 ( 
.A(n_4002),
.B(n_4003),
.Y(n_4224)
);

AND2x2_ASAP7_75t_L g4225 ( 
.A(n_3936),
.B(n_3710),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_4002),
.B(n_3633),
.Y(n_4226)
);

AND2x4_ASAP7_75t_L g4227 ( 
.A(n_3916),
.B(n_3694),
.Y(n_4227)
);

NAND2x1_ASAP7_75t_SL g4228 ( 
.A(n_3984),
.B(n_3989),
.Y(n_4228)
);

NOR2xp33_ASAP7_75t_L g4229 ( 
.A(n_3934),
.B(n_3537),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_3949),
.Y(n_4230)
);

OR2x2_ASAP7_75t_L g4231 ( 
.A(n_4070),
.B(n_3737),
.Y(n_4231)
);

AND2x2_ASAP7_75t_L g4232 ( 
.A(n_3944),
.B(n_3710),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_3956),
.B(n_3844),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_3894),
.Y(n_4234)
);

OR2x2_ASAP7_75t_L g4235 ( 
.A(n_4039),
.B(n_3747),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_3897),
.Y(n_4236)
);

OR2x2_ASAP7_75t_L g4237 ( 
.A(n_4086),
.B(n_3747),
.Y(n_4237)
);

HB1xp67_ASAP7_75t_L g4238 ( 
.A(n_3965),
.Y(n_4238)
);

NAND3xp33_ASAP7_75t_L g4239 ( 
.A(n_4075),
.B(n_3760),
.C(n_3810),
.Y(n_4239)
);

INVx4_ASAP7_75t_L g4240 ( 
.A(n_3924),
.Y(n_4240)
);

INVx2_ASAP7_75t_L g4241 ( 
.A(n_3957),
.Y(n_4241)
);

OR2x2_ASAP7_75t_L g4242 ( 
.A(n_3982),
.B(n_3747),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_3897),
.Y(n_4243)
);

AND2x2_ASAP7_75t_L g4244 ( 
.A(n_3913),
.B(n_3817),
.Y(n_4244)
);

INVx2_ASAP7_75t_L g4245 ( 
.A(n_3958),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_3962),
.Y(n_4246)
);

AND2x4_ASAP7_75t_L g4247 ( 
.A(n_3935),
.B(n_3726),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_4003),
.B(n_3744),
.Y(n_4248)
);

HB1xp67_ASAP7_75t_L g4249 ( 
.A(n_4015),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_4139),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4144),
.Y(n_4251)
);

INVxp67_ASAP7_75t_SL g4252 ( 
.A(n_4220),
.Y(n_4252)
);

INVx2_ASAP7_75t_L g4253 ( 
.A(n_4137),
.Y(n_4253)
);

HB1xp67_ASAP7_75t_L g4254 ( 
.A(n_4162),
.Y(n_4254)
);

BUFx2_ASAP7_75t_L g4255 ( 
.A(n_4134),
.Y(n_4255)
);

OR2x2_ASAP7_75t_L g4256 ( 
.A(n_4138),
.B(n_4115),
.Y(n_4256)
);

INVx3_ASAP7_75t_L g4257 ( 
.A(n_4135),
.Y(n_4257)
);

INVx3_ASAP7_75t_L g4258 ( 
.A(n_4135),
.Y(n_4258)
);

AND2x2_ASAP7_75t_L g4259 ( 
.A(n_4161),
.B(n_4133),
.Y(n_4259)
);

OR2x2_ASAP7_75t_L g4260 ( 
.A(n_4175),
.B(n_4027),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4165),
.Y(n_4261)
);

INVx2_ASAP7_75t_L g4262 ( 
.A(n_4157),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4176),
.Y(n_4263)
);

OR2x2_ASAP7_75t_L g4264 ( 
.A(n_4177),
.B(n_4027),
.Y(n_4264)
);

INVx5_ASAP7_75t_L g4265 ( 
.A(n_4240),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_4235),
.Y(n_4266)
);

OR2x2_ASAP7_75t_L g4267 ( 
.A(n_4166),
.B(n_4028),
.Y(n_4267)
);

BUFx2_ASAP7_75t_L g4268 ( 
.A(n_4132),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_4147),
.B(n_4029),
.Y(n_4269)
);

HB1xp67_ASAP7_75t_L g4270 ( 
.A(n_4149),
.Y(n_4270)
);

BUFx2_ASAP7_75t_L g4271 ( 
.A(n_4228),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4180),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4182),
.Y(n_4273)
);

INVx2_ASAP7_75t_L g4274 ( 
.A(n_4141),
.Y(n_4274)
);

HB1xp67_ASAP7_75t_L g4275 ( 
.A(n_4172),
.Y(n_4275)
);

AND2x2_ASAP7_75t_L g4276 ( 
.A(n_4194),
.B(n_3935),
.Y(n_4276)
);

NOR2xp67_ASAP7_75t_L g4277 ( 
.A(n_4240),
.B(n_3989),
.Y(n_4277)
);

BUFx2_ASAP7_75t_L g4278 ( 
.A(n_4131),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4184),
.Y(n_4279)
);

OR2x2_ASAP7_75t_L g4280 ( 
.A(n_4140),
.B(n_4028),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4186),
.Y(n_4281)
);

INVx2_ASAP7_75t_SL g4282 ( 
.A(n_4219),
.Y(n_4282)
);

INVx2_ASAP7_75t_L g4283 ( 
.A(n_4152),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4188),
.Y(n_4284)
);

OR2x2_ASAP7_75t_L g4285 ( 
.A(n_4160),
.B(n_4029),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4136),
.B(n_4067),
.Y(n_4286)
);

AND2x4_ASAP7_75t_SL g4287 ( 
.A(n_4207),
.B(n_3890),
.Y(n_4287)
);

INVx2_ASAP7_75t_L g4288 ( 
.A(n_4153),
.Y(n_4288)
);

AND2x2_ASAP7_75t_L g4289 ( 
.A(n_4249),
.B(n_4076),
.Y(n_4289)
);

AND2x2_ASAP7_75t_L g4290 ( 
.A(n_4202),
.B(n_4078),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_4154),
.B(n_4142),
.Y(n_4291)
);

AND2x2_ASAP7_75t_L g4292 ( 
.A(n_4168),
.B(n_3941),
.Y(n_4292)
);

AND2x4_ASAP7_75t_L g4293 ( 
.A(n_4221),
.B(n_3941),
.Y(n_4293)
);

INVx3_ASAP7_75t_L g4294 ( 
.A(n_4227),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4190),
.Y(n_4295)
);

AND2x2_ASAP7_75t_L g4296 ( 
.A(n_4196),
.B(n_3960),
.Y(n_4296)
);

AND2x2_ASAP7_75t_L g4297 ( 
.A(n_4238),
.B(n_3960),
.Y(n_4297)
);

AND2x2_ASAP7_75t_L g4298 ( 
.A(n_4167),
.B(n_4233),
.Y(n_4298)
);

OR2x2_ASAP7_75t_L g4299 ( 
.A(n_4208),
.B(n_4032),
.Y(n_4299)
);

AND2x4_ASAP7_75t_L g4300 ( 
.A(n_4173),
.B(n_3987),
.Y(n_4300)
);

INVxp33_ASAP7_75t_L g4301 ( 
.A(n_4163),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_4159),
.B(n_4032),
.Y(n_4302)
);

INVx1_ASAP7_75t_SL g4303 ( 
.A(n_4210),
.Y(n_4303)
);

INVx3_ASAP7_75t_L g4304 ( 
.A(n_4227),
.Y(n_4304)
);

AND2x2_ASAP7_75t_L g4305 ( 
.A(n_4204),
.B(n_3976),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4203),
.Y(n_4306)
);

AND2x2_ASAP7_75t_L g4307 ( 
.A(n_4155),
.B(n_3976),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_4174),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_4158),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4224),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_4173),
.B(n_3979),
.Y(n_4311)
);

INVx1_ASAP7_75t_SL g4312 ( 
.A(n_4187),
.Y(n_4312)
);

AND2x2_ASAP7_75t_L g4313 ( 
.A(n_4178),
.B(n_3979),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_4148),
.B(n_4145),
.Y(n_4314)
);

AND2x2_ASAP7_75t_L g4315 ( 
.A(n_4178),
.B(n_3920),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4174),
.Y(n_4316)
);

AND2x4_ASAP7_75t_SL g4317 ( 
.A(n_4207),
.B(n_3890),
.Y(n_4317)
);

OR2x2_ASAP7_75t_L g4318 ( 
.A(n_4201),
.B(n_4056),
.Y(n_4318)
);

NAND4xp75_ASAP7_75t_L g4319 ( 
.A(n_4192),
.B(n_3971),
.C(n_4092),
.D(n_3731),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_4189),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4212),
.Y(n_4321)
);

INVx2_ASAP7_75t_L g4322 ( 
.A(n_4191),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_4244),
.B(n_4225),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4232),
.B(n_4122),
.Y(n_4324)
);

INVx2_ASAP7_75t_SL g4325 ( 
.A(n_4169),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4212),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4214),
.Y(n_4327)
);

HB1xp67_ASAP7_75t_L g4328 ( 
.A(n_4156),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4214),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_4218),
.B(n_4124),
.Y(n_4330)
);

AND2x4_ASAP7_75t_L g4331 ( 
.A(n_4146),
.B(n_3988),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_4170),
.B(n_4123),
.Y(n_4332)
);

CKINVDCx16_ASAP7_75t_R g4333 ( 
.A(n_4200),
.Y(n_4333)
);

NAND2x1_ASAP7_75t_L g4334 ( 
.A(n_4247),
.B(n_3905),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_4151),
.B(n_4069),
.Y(n_4335)
);

AND2x2_ASAP7_75t_L g4336 ( 
.A(n_4197),
.B(n_4016),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4205),
.B(n_4019),
.Y(n_4337)
);

AND2x2_ASAP7_75t_L g4338 ( 
.A(n_4150),
.B(n_4024),
.Y(n_4338)
);

AND2x2_ASAP7_75t_L g4339 ( 
.A(n_4150),
.B(n_4063),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_4269),
.B(n_4226),
.Y(n_4340)
);

INVxp67_ASAP7_75t_L g4341 ( 
.A(n_4255),
.Y(n_4341)
);

AND2x2_ASAP7_75t_L g4342 ( 
.A(n_4338),
.B(n_4324),
.Y(n_4342)
);

AOI22xp5_ASAP7_75t_L g4343 ( 
.A1(n_4319),
.A2(n_4223),
.B1(n_4183),
.B2(n_4198),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4252),
.Y(n_4344)
);

OAI322xp33_ASAP7_75t_L g4345 ( 
.A1(n_4285),
.A2(n_4193),
.A3(n_4164),
.B1(n_4222),
.B2(n_4074),
.C1(n_4072),
.C2(n_3985),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4252),
.Y(n_4346)
);

AND2x2_ASAP7_75t_L g4347 ( 
.A(n_4339),
.B(n_4185),
.Y(n_4347)
);

INVx2_ASAP7_75t_SL g4348 ( 
.A(n_4287),
.Y(n_4348)
);

NOR2xp33_ASAP7_75t_L g4349 ( 
.A(n_4333),
.B(n_4129),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4270),
.Y(n_4350)
);

OAI21xp5_ASAP7_75t_L g4351 ( 
.A1(n_4277),
.A2(n_4239),
.B(n_4108),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_4270),
.Y(n_4352)
);

NAND4xp25_ASAP7_75t_L g4353 ( 
.A(n_4268),
.B(n_4195),
.C(n_3712),
.D(n_3690),
.Y(n_4353)
);

INVx5_ASAP7_75t_L g4354 ( 
.A(n_4265),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_4296),
.B(n_4199),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4275),
.Y(n_4356)
);

AOI22xp5_ASAP7_75t_L g4357 ( 
.A1(n_4277),
.A2(n_3835),
.B1(n_3728),
.B2(n_3568),
.Y(n_4357)
);

NOR2xp33_ASAP7_75t_L g4358 ( 
.A(n_4287),
.B(n_4317),
.Y(n_4358)
);

A2O1A1Ixp33_ASAP7_75t_L g4359 ( 
.A1(n_4334),
.A2(n_4077),
.B(n_4007),
.C(n_4011),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_SL g4360 ( 
.A(n_4265),
.B(n_4271),
.Y(n_4360)
);

INVx1_ASAP7_75t_SL g4361 ( 
.A(n_4303),
.Y(n_4361)
);

AND2x2_ASAP7_75t_L g4362 ( 
.A(n_4297),
.B(n_4199),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_4300),
.B(n_4146),
.Y(n_4363)
);

HB1xp67_ASAP7_75t_L g4364 ( 
.A(n_4254),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4275),
.Y(n_4365)
);

XOR2x2_ASAP7_75t_L g4366 ( 
.A(n_4303),
.B(n_3929),
.Y(n_4366)
);

INVxp67_ASAP7_75t_SL g4367 ( 
.A(n_4254),
.Y(n_4367)
);

AOI32xp33_ASAP7_75t_L g4368 ( 
.A1(n_4301),
.A2(n_4126),
.A3(n_4050),
.B1(n_3950),
.B2(n_4006),
.Y(n_4368)
);

INVx2_ASAP7_75t_L g4369 ( 
.A(n_4266),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4256),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4250),
.Y(n_4371)
);

OAI211xp5_ASAP7_75t_SL g4372 ( 
.A1(n_4335),
.A2(n_4181),
.B(n_4179),
.C(n_4052),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4251),
.Y(n_4373)
);

AOI22xp5_ASAP7_75t_L g4374 ( 
.A1(n_4265),
.A2(n_4143),
.B1(n_3964),
.B2(n_3843),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4261),
.Y(n_4375)
);

INVx2_ASAP7_75t_L g4376 ( 
.A(n_4266),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_4308),
.Y(n_4377)
);

NAND2xp33_ASAP7_75t_SL g4378 ( 
.A(n_4301),
.B(n_4089),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4263),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_4269),
.B(n_4248),
.Y(n_4380)
);

OR2x2_ASAP7_75t_L g4381 ( 
.A(n_4267),
.B(n_4242),
.Y(n_4381)
);

INVxp67_ASAP7_75t_L g4382 ( 
.A(n_4278),
.Y(n_4382)
);

INVxp67_ASAP7_75t_SL g4383 ( 
.A(n_4328),
.Y(n_4383)
);

AND2x4_ASAP7_75t_SL g4384 ( 
.A(n_4282),
.B(n_4089),
.Y(n_4384)
);

INVxp67_ASAP7_75t_SL g4385 ( 
.A(n_4328),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4272),
.Y(n_4386)
);

AND2x2_ASAP7_75t_L g4387 ( 
.A(n_4300),
.B(n_4247),
.Y(n_4387)
);

AND2x2_ASAP7_75t_L g4388 ( 
.A(n_4312),
.B(n_4215),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4273),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_SL g4390 ( 
.A(n_4265),
.B(n_4089),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4279),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4308),
.Y(n_4392)
);

OAI322xp33_ASAP7_75t_L g4393 ( 
.A1(n_4335),
.A2(n_4110),
.A3(n_4217),
.B1(n_4096),
.B2(n_4030),
.C1(n_4231),
.C2(n_4211),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_SL g4394 ( 
.A(n_4257),
.B(n_3938),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4281),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_L g4396 ( 
.A(n_4314),
.B(n_4071),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4284),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4295),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_4306),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4316),
.Y(n_4400)
);

AND2x2_ASAP7_75t_L g4401 ( 
.A(n_4312),
.B(n_4206),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_SL g4402 ( 
.A(n_4257),
.B(n_3938),
.Y(n_4402)
);

AND2x2_ASAP7_75t_L g4403 ( 
.A(n_4331),
.B(n_4213),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4321),
.Y(n_4404)
);

INVx2_ASAP7_75t_L g4405 ( 
.A(n_4274),
.Y(n_4405)
);

INVx2_ASAP7_75t_L g4406 ( 
.A(n_4283),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4326),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4327),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4329),
.Y(n_4409)
);

NOR4xp25_ASAP7_75t_L g4410 ( 
.A(n_4325),
.B(n_4229),
.C(n_3955),
.D(n_3790),
.Y(n_4410)
);

NOR3xp33_ASAP7_75t_L g4411 ( 
.A(n_4302),
.B(n_4017),
.C(n_3578),
.Y(n_4411)
);

INVx3_ASAP7_75t_L g4412 ( 
.A(n_4258),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4310),
.Y(n_4413)
);

AND2x4_ASAP7_75t_L g4414 ( 
.A(n_4293),
.B(n_4236),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_4411),
.B(n_4302),
.Y(n_4415)
);

O2A1O1Ixp33_ASAP7_75t_L g4416 ( 
.A1(n_4410),
.A2(n_4262),
.B(n_4121),
.C(n_3986),
.Y(n_4416)
);

AOI22xp33_ASAP7_75t_L g4417 ( 
.A1(n_4343),
.A2(n_4331),
.B1(n_4304),
.B2(n_4294),
.Y(n_4417)
);

OAI21xp5_ASAP7_75t_L g4418 ( 
.A1(n_4359),
.A2(n_3932),
.B(n_4258),
.Y(n_4418)
);

XNOR2xp5_ASAP7_75t_L g4419 ( 
.A(n_4366),
.B(n_3550),
.Y(n_4419)
);

AOI22xp5_ASAP7_75t_L g4420 ( 
.A1(n_4353),
.A2(n_4289),
.B1(n_4253),
.B2(n_4305),
.Y(n_4420)
);

NOR3xp33_ASAP7_75t_L g4421 ( 
.A(n_4351),
.B(n_3591),
.C(n_3908),
.Y(n_4421)
);

NOR3xp33_ASAP7_75t_L g4422 ( 
.A(n_4393),
.B(n_3734),
.C(n_3729),
.Y(n_4422)
);

INVxp67_ASAP7_75t_L g4423 ( 
.A(n_4349),
.Y(n_4423)
);

OAI21xp5_ASAP7_75t_L g4424 ( 
.A1(n_4383),
.A2(n_4293),
.B(n_4119),
.Y(n_4424)
);

A2O1A1Ixp33_ASAP7_75t_L g4425 ( 
.A1(n_4368),
.A2(n_4317),
.B(n_4081),
.C(n_4109),
.Y(n_4425)
);

INVx1_ASAP7_75t_L g4426 ( 
.A(n_4364),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4350),
.Y(n_4427)
);

OAI21xp5_ASAP7_75t_L g4428 ( 
.A1(n_4385),
.A2(n_4116),
.B(n_3938),
.Y(n_4428)
);

NOR3xp33_ASAP7_75t_L g4429 ( 
.A(n_4372),
.B(n_3668),
.C(n_3709),
.Y(n_4429)
);

AOI21xp5_ASAP7_75t_L g4430 ( 
.A1(n_4390),
.A2(n_4171),
.B(n_4294),
.Y(n_4430)
);

NAND3xp33_ASAP7_75t_L g4431 ( 
.A(n_4344),
.B(n_3616),
.C(n_3819),
.Y(n_4431)
);

INVxp67_ASAP7_75t_L g4432 ( 
.A(n_4367),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_SL g4433 ( 
.A(n_4354),
.B(n_4304),
.Y(n_4433)
);

AOI22xp5_ASAP7_75t_L g4434 ( 
.A1(n_4382),
.A2(n_4332),
.B1(n_4276),
.B2(n_4307),
.Y(n_4434)
);

INVx2_ASAP7_75t_L g4435 ( 
.A(n_4361),
.Y(n_4435)
);

INVxp33_ASAP7_75t_SL g4436 ( 
.A(n_4357),
.Y(n_4436)
);

OAI21xp33_ASAP7_75t_L g4437 ( 
.A1(n_4340),
.A2(n_4318),
.B(n_4299),
.Y(n_4437)
);

OAI22xp5_ASAP7_75t_L g4438 ( 
.A1(n_4348),
.A2(n_4280),
.B1(n_4292),
.B2(n_4315),
.Y(n_4438)
);

AO22x1_ASAP7_75t_L g4439 ( 
.A1(n_4354),
.A2(n_3707),
.B1(n_3553),
.B2(n_3742),
.Y(n_4439)
);

NAND4xp75_ASAP7_75t_L g4440 ( 
.A(n_4360),
.B(n_3506),
.C(n_4120),
.D(n_4023),
.Y(n_4440)
);

OAI21xp5_ASAP7_75t_L g4441 ( 
.A1(n_4341),
.A2(n_3604),
.B(n_4114),
.Y(n_4441)
);

OAI21xp33_ASAP7_75t_L g4442 ( 
.A1(n_4380),
.A2(n_4264),
.B(n_4260),
.Y(n_4442)
);

AOI21xp33_ASAP7_75t_L g4443 ( 
.A1(n_4374),
.A2(n_3722),
.B(n_3572),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_4352),
.Y(n_4444)
);

INVxp67_ASAP7_75t_L g4445 ( 
.A(n_4356),
.Y(n_4445)
);

OAI211xp5_ASAP7_75t_SL g4446 ( 
.A1(n_4346),
.A2(n_3884),
.B(n_3605),
.C(n_4034),
.Y(n_4446)
);

INVxp67_ASAP7_75t_L g4447 ( 
.A(n_4365),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_4369),
.Y(n_4448)
);

AOI22xp5_ASAP7_75t_L g4449 ( 
.A1(n_4378),
.A2(n_4330),
.B1(n_4298),
.B2(n_4336),
.Y(n_4449)
);

AOI221xp5_ASAP7_75t_L g4450 ( 
.A1(n_4345),
.A2(n_4286),
.B1(n_4259),
.B2(n_4337),
.C(n_4290),
.Y(n_4450)
);

OAI22xp33_ASAP7_75t_L g4451 ( 
.A1(n_4354),
.A2(n_4412),
.B1(n_4381),
.B2(n_4402),
.Y(n_4451)
);

OAI21xp5_ASAP7_75t_L g4452 ( 
.A1(n_4412),
.A2(n_3604),
.B(n_3673),
.Y(n_4452)
);

INVxp67_ASAP7_75t_SL g4453 ( 
.A(n_4405),
.Y(n_4453)
);

NAND3xp33_ASAP7_75t_L g4454 ( 
.A(n_4413),
.B(n_3814),
.C(n_4237),
.Y(n_4454)
);

AOI211xp5_ASAP7_75t_SL g4455 ( 
.A1(n_4358),
.A2(n_3596),
.B(n_3620),
.C(n_3951),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_L g4456 ( 
.A(n_4370),
.B(n_4396),
.Y(n_4456)
);

NAND3xp33_ASAP7_75t_L g4457 ( 
.A(n_4371),
.B(n_3756),
.C(n_4118),
.Y(n_4457)
);

AOI22xp33_ASAP7_75t_L g4458 ( 
.A1(n_4414),
.A2(n_4036),
.B1(n_4031),
.B2(n_4041),
.Y(n_4458)
);

OAI21xp5_ASAP7_75t_L g4459 ( 
.A1(n_4414),
.A2(n_4291),
.B(n_3699),
.Y(n_4459)
);

OAI221xp5_ASAP7_75t_L g4460 ( 
.A1(n_4373),
.A2(n_4043),
.B1(n_4033),
.B2(n_3852),
.C(n_3663),
.Y(n_4460)
);

AND2x2_ASAP7_75t_SL g4461 ( 
.A(n_4384),
.B(n_3951),
.Y(n_4461)
);

NAND2xp33_ASAP7_75t_SL g4462 ( 
.A(n_4387),
.B(n_3625),
.Y(n_4462)
);

AOI22xp5_ASAP7_75t_L g4463 ( 
.A1(n_4388),
.A2(n_4313),
.B1(n_4311),
.B2(n_4323),
.Y(n_4463)
);

AND2x2_ASAP7_75t_L g4464 ( 
.A(n_4363),
.B(n_4288),
.Y(n_4464)
);

OAI21xp5_ASAP7_75t_L g4465 ( 
.A1(n_4394),
.A2(n_3663),
.B(n_4005),
.Y(n_4465)
);

AOI21xp5_ASAP7_75t_L g4466 ( 
.A1(n_4403),
.A2(n_4005),
.B(n_4309),
.Y(n_4466)
);

NOR2xp33_ASAP7_75t_L g4467 ( 
.A(n_4436),
.B(n_3522),
.Y(n_4467)
);

OAI22xp5_ASAP7_75t_L g4468 ( 
.A1(n_4417),
.A2(n_4355),
.B1(n_4362),
.B2(n_4347),
.Y(n_4468)
);

OAI221xp5_ASAP7_75t_SL g4469 ( 
.A1(n_4420),
.A2(n_4401),
.B1(n_4037),
.B2(n_3669),
.C(n_4379),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4435),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4426),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4415),
.B(n_4375),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4432),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4456),
.Y(n_4474)
);

AOI22xp5_ASAP7_75t_L g4475 ( 
.A1(n_4440),
.A2(n_4389),
.B1(n_4391),
.B2(n_4386),
.Y(n_4475)
);

AOI221xp5_ASAP7_75t_L g4476 ( 
.A1(n_4416),
.A2(n_4397),
.B1(n_4399),
.B2(n_4398),
.C(n_4395),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_L g4477 ( 
.A(n_4437),
.B(n_4400),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_4442),
.B(n_4404),
.Y(n_4478)
);

OAI21xp5_ASAP7_75t_L g4479 ( 
.A1(n_4425),
.A2(n_4408),
.B(n_4407),
.Y(n_4479)
);

AND2x2_ASAP7_75t_L g4480 ( 
.A(n_4461),
.B(n_4342),
.Y(n_4480)
);

A2O1A1Ixp33_ASAP7_75t_L g4481 ( 
.A1(n_4462),
.A2(n_3904),
.B(n_4073),
.C(n_3746),
.Y(n_4481)
);

OAI22xp5_ASAP7_75t_L g4482 ( 
.A1(n_4449),
.A2(n_4376),
.B1(n_4409),
.B2(n_4406),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_4445),
.B(n_4392),
.Y(n_4483)
);

AND2x4_ASAP7_75t_L g4484 ( 
.A(n_4452),
.B(n_4392),
.Y(n_4484)
);

OAI211xp5_ASAP7_75t_L g4485 ( 
.A1(n_4418),
.A2(n_4441),
.B(n_4443),
.C(n_4455),
.Y(n_4485)
);

NOR2xp33_ASAP7_75t_L g4486 ( 
.A(n_4419),
.B(n_4423),
.Y(n_4486)
);

NAND2x1p5_ASAP7_75t_L g4487 ( 
.A(n_4430),
.B(n_4433),
.Y(n_4487)
);

AOI21xp33_ASAP7_75t_L g4488 ( 
.A1(n_4460),
.A2(n_3770),
.B(n_3829),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4427),
.Y(n_4489)
);

AOI211xp5_ASAP7_75t_L g4490 ( 
.A1(n_4451),
.A2(n_3540),
.B(n_3741),
.C(n_3664),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4444),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_4447),
.B(n_4377),
.Y(n_4492)
);

AOI211xp5_ASAP7_75t_L g4493 ( 
.A1(n_4439),
.A2(n_3566),
.B(n_3644),
.C(n_3622),
.Y(n_4493)
);

OAI21xp5_ASAP7_75t_SL g4494 ( 
.A1(n_4455),
.A2(n_4068),
.B(n_4049),
.Y(n_4494)
);

OAI22xp33_ASAP7_75t_L g4495 ( 
.A1(n_4424),
.A2(n_3775),
.B1(n_4322),
.B2(n_4320),
.Y(n_4495)
);

AOI21xp5_ASAP7_75t_L g4496 ( 
.A1(n_4466),
.A2(n_3655),
.B(n_3773),
.Y(n_4496)
);

AOI21xp33_ASAP7_75t_L g4497 ( 
.A1(n_4454),
.A2(n_4042),
.B(n_4038),
.Y(n_4497)
);

HB1xp67_ASAP7_75t_L g4498 ( 
.A(n_4453),
.Y(n_4498)
);

AOI21xp33_ASAP7_75t_L g4499 ( 
.A1(n_4446),
.A2(n_3809),
.B(n_4118),
.Y(n_4499)
);

INVxp67_ASAP7_75t_SL g4500 ( 
.A(n_4429),
.Y(n_4500)
);

OR2x2_ASAP7_75t_L g4501 ( 
.A(n_4448),
.B(n_4246),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4438),
.Y(n_4502)
);

OAI21xp5_ASAP7_75t_L g4503 ( 
.A1(n_4459),
.A2(n_3841),
.B(n_3708),
.Y(n_4503)
);

O2A1O1Ixp33_ASAP7_75t_L g4504 ( 
.A1(n_4422),
.A2(n_3777),
.B(n_3748),
.C(n_3623),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4464),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4434),
.Y(n_4506)
);

HB1xp67_ASAP7_75t_L g4507 ( 
.A(n_4428),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_4450),
.B(n_4236),
.Y(n_4508)
);

O2A1O1Ixp33_ASAP7_75t_L g4509 ( 
.A1(n_4421),
.A2(n_3623),
.B(n_3877),
.C(n_3861),
.Y(n_4509)
);

AND2x2_ASAP7_75t_L g4510 ( 
.A(n_4463),
.B(n_4020),
.Y(n_4510)
);

OR2x2_ASAP7_75t_L g4511 ( 
.A(n_4458),
.B(n_4245),
.Y(n_4511)
);

INVx2_ASAP7_75t_L g4512 ( 
.A(n_4431),
.Y(n_4512)
);

OAI22xp33_ASAP7_75t_L g4513 ( 
.A1(n_4465),
.A2(n_4216),
.B1(n_4241),
.B2(n_4230),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4457),
.Y(n_4514)
);

OAI22xp5_ASAP7_75t_SL g4515 ( 
.A1(n_4419),
.A2(n_3691),
.B1(n_3685),
.B2(n_4064),
.Y(n_4515)
);

INVx3_ASAP7_75t_L g4516 ( 
.A(n_4461),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_4415),
.B(n_4243),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_4461),
.B(n_4064),
.Y(n_4518)
);

OAI21xp33_ASAP7_75t_L g4519 ( 
.A1(n_4436),
.A2(n_4082),
.B(n_4243),
.Y(n_4519)
);

NOR3xp33_ASAP7_75t_L g4520 ( 
.A(n_4440),
.B(n_3391),
.C(n_3370),
.Y(n_4520)
);

OA211x2_ASAP7_75t_L g4521 ( 
.A1(n_4418),
.A2(n_3697),
.B(n_3855),
.C(n_3825),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_4502),
.B(n_4209),
.Y(n_4522)
);

INVxp67_ASAP7_75t_L g4523 ( 
.A(n_4467),
.Y(n_4523)
);

OA22x2_ASAP7_75t_L g4524 ( 
.A1(n_4485),
.A2(n_4083),
.B1(n_4234),
.B2(n_4022),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_SL g4525 ( 
.A(n_4498),
.B(n_3520),
.Y(n_4525)
);

AND2x2_ASAP7_75t_L g4526 ( 
.A(n_4487),
.B(n_4083),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_SL g4527 ( 
.A(n_4476),
.B(n_3516),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_L g4528 ( 
.A(n_4500),
.B(n_4009),
.Y(n_4528)
);

NOR2xp33_ASAP7_75t_L g4529 ( 
.A(n_4486),
.B(n_3695),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_SL g4530 ( 
.A(n_4516),
.B(n_4495),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_4501),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_4470),
.Y(n_4532)
);

OAI21xp5_ASAP7_75t_L g4533 ( 
.A1(n_4504),
.A2(n_4004),
.B(n_3154),
.Y(n_4533)
);

AOI21xp5_ASAP7_75t_L g4534 ( 
.A1(n_4515),
.A2(n_3876),
.B(n_4062),
.Y(n_4534)
);

OAI221xp5_ASAP7_75t_SL g4535 ( 
.A1(n_4494),
.A2(n_4087),
.B1(n_4009),
.B2(n_3903),
.C(n_3931),
.Y(n_4535)
);

NOR3x1_ASAP7_75t_L g4536 ( 
.A(n_4506),
.B(n_3859),
.C(n_3857),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4473),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_4474),
.B(n_3900),
.Y(n_4538)
);

NAND3xp33_ASAP7_75t_SL g4539 ( 
.A(n_4512),
.B(n_3808),
.C(n_3517),
.Y(n_4539)
);

NOR2xp67_ASAP7_75t_L g4540 ( 
.A(n_4516),
.B(n_756),
.Y(n_4540)
);

INVx2_ASAP7_75t_L g4541 ( 
.A(n_4505),
.Y(n_4541)
);

NOR3xp33_ASAP7_75t_L g4542 ( 
.A(n_4520),
.B(n_3202),
.C(n_4128),
.Y(n_4542)
);

OR2x2_ASAP7_75t_L g4543 ( 
.A(n_4517),
.B(n_4127),
.Y(n_4543)
);

AOI221xp5_ASAP7_75t_L g4544 ( 
.A1(n_4514),
.A2(n_3900),
.B1(n_3931),
.B2(n_3903),
.C(n_3901),
.Y(n_4544)
);

AOI21xp5_ASAP7_75t_L g4545 ( 
.A1(n_4490),
.A2(n_3942),
.B(n_3911),
.Y(n_4545)
);

INVx2_ASAP7_75t_SL g4546 ( 
.A(n_4518),
.Y(n_4546)
);

INVx1_ASAP7_75t_SL g4547 ( 
.A(n_4488),
.Y(n_4547)
);

NOR2x1_ASAP7_75t_L g4548 ( 
.A(n_4481),
.B(n_3793),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4471),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4489),
.Y(n_4550)
);

OAI21xp33_ASAP7_75t_SL g4551 ( 
.A1(n_4480),
.A2(n_4475),
.B(n_4507),
.Y(n_4551)
);

AOI211xp5_ASAP7_75t_L g4552 ( 
.A1(n_4469),
.A2(n_3785),
.B(n_3816),
.C(n_4094),
.Y(n_4552)
);

NOR2xp33_ASAP7_75t_L g4553 ( 
.A(n_4468),
.B(n_3850),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_4491),
.Y(n_4554)
);

OAI21xp33_ASAP7_75t_L g4555 ( 
.A1(n_4508),
.A2(n_4519),
.B(n_4497),
.Y(n_4555)
);

NAND2xp5_ASAP7_75t_SL g4556 ( 
.A(n_4496),
.B(n_3848),
.Y(n_4556)
);

NAND2xp5_ASAP7_75t_L g4557 ( 
.A(n_4555),
.B(n_4472),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_L g4558 ( 
.A(n_4523),
.B(n_4477),
.Y(n_4558)
);

AO22x2_ASAP7_75t_L g4559 ( 
.A1(n_4537),
.A2(n_4482),
.B1(n_4478),
.B2(n_4484),
.Y(n_4559)
);

NOR3xp33_ASAP7_75t_L g4560 ( 
.A(n_4551),
.B(n_4503),
.C(n_4499),
.Y(n_4560)
);

AOI22xp5_ASAP7_75t_L g4561 ( 
.A1(n_4551),
.A2(n_4521),
.B1(n_4484),
.B2(n_4513),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4532),
.Y(n_4562)
);

INVxp67_ASAP7_75t_L g4563 ( 
.A(n_4529),
.Y(n_4563)
);

AOI22xp33_ASAP7_75t_L g4564 ( 
.A1(n_4524),
.A2(n_4479),
.B1(n_4510),
.B2(n_4511),
.Y(n_4564)
);

AND2x2_ASAP7_75t_L g4565 ( 
.A(n_4526),
.B(n_4493),
.Y(n_4565)
);

AOI211xp5_ASAP7_75t_L g4566 ( 
.A1(n_4530),
.A2(n_4547),
.B(n_4540),
.C(n_4533),
.Y(n_4566)
);

AOI21xp5_ASAP7_75t_L g4567 ( 
.A1(n_4556),
.A2(n_4483),
.B(n_4492),
.Y(n_4567)
);

INVxp67_ASAP7_75t_SL g4568 ( 
.A(n_4528),
.Y(n_4568)
);

OAI21xp33_ASAP7_75t_SL g4569 ( 
.A1(n_4546),
.A2(n_4509),
.B(n_3947),
.Y(n_4569)
);

AOI21xp5_ASAP7_75t_L g4570 ( 
.A1(n_4525),
.A2(n_3983),
.B(n_4094),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4538),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4541),
.Y(n_4572)
);

NOR2x1_ASAP7_75t_L g4573 ( 
.A(n_4548),
.B(n_4553),
.Y(n_4573)
);

INVxp67_ASAP7_75t_L g4574 ( 
.A(n_4549),
.Y(n_4574)
);

NOR3xp33_ASAP7_75t_L g4575 ( 
.A(n_4535),
.B(n_3125),
.C(n_3875),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4531),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_L g4577 ( 
.A(n_4522),
.B(n_3901),
.Y(n_4577)
);

AOI21xp5_ASAP7_75t_L g4578 ( 
.A1(n_4527),
.A2(n_4101),
.B(n_4098),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4550),
.Y(n_4579)
);

AOI21xp33_ASAP7_75t_L g4580 ( 
.A1(n_4554),
.A2(n_757),
.B(n_758),
.Y(n_4580)
);

NOR3xp33_ASAP7_75t_L g4581 ( 
.A(n_4542),
.B(n_4101),
.C(n_4098),
.Y(n_4581)
);

AO22x2_ASAP7_75t_L g4582 ( 
.A1(n_4534),
.A2(n_4060),
.B1(n_4061),
.B2(n_4046),
.Y(n_4582)
);

AOI211xp5_ASAP7_75t_SL g4583 ( 
.A1(n_4552),
.A2(n_4106),
.B(n_4113),
.C(n_4102),
.Y(n_4583)
);

O2A1O1Ixp33_ASAP7_75t_L g4584 ( 
.A1(n_4560),
.A2(n_4566),
.B(n_4558),
.C(n_4563),
.Y(n_4584)
);

OAI21xp5_ASAP7_75t_L g4585 ( 
.A1(n_4561),
.A2(n_4545),
.B(n_4539),
.Y(n_4585)
);

AOI322xp5_ASAP7_75t_L g4586 ( 
.A1(n_4564),
.A2(n_4557),
.A3(n_4573),
.B1(n_4568),
.B2(n_4569),
.C1(n_4565),
.C2(n_4576),
.Y(n_4586)
);

NOR2xp33_ASAP7_75t_R g4587 ( 
.A(n_4579),
.B(n_759),
.Y(n_4587)
);

AOI221xp5_ASAP7_75t_L g4588 ( 
.A1(n_4559),
.A2(n_4544),
.B1(n_4543),
.B2(n_4536),
.C(n_4113),
.Y(n_4588)
);

OAI221xp5_ASAP7_75t_SL g4589 ( 
.A1(n_4575),
.A2(n_4106),
.B1(n_4102),
.B2(n_3864),
.C(n_3851),
.Y(n_4589)
);

AOI21xp5_ASAP7_75t_L g4590 ( 
.A1(n_4559),
.A2(n_3780),
.B(n_3767),
.Y(n_4590)
);

AOI211xp5_ASAP7_75t_SL g4591 ( 
.A1(n_4580),
.A2(n_762),
.B(n_760),
.C(n_761),
.Y(n_4591)
);

AOI211xp5_ASAP7_75t_L g4592 ( 
.A1(n_4574),
.A2(n_4053),
.B(n_3953),
.C(n_3954),
.Y(n_4592)
);

AOI21xp33_ASAP7_75t_SL g4593 ( 
.A1(n_4582),
.A2(n_4572),
.B(n_4562),
.Y(n_4593)
);

NAND3xp33_ASAP7_75t_L g4594 ( 
.A(n_4583),
.B(n_2815),
.C(n_2791),
.Y(n_4594)
);

OAI211xp5_ASAP7_75t_L g4595 ( 
.A1(n_4567),
.A2(n_3283),
.B(n_4079),
.C(n_4065),
.Y(n_4595)
);

AOI211xp5_ASAP7_75t_SL g4596 ( 
.A1(n_4571),
.A2(n_764),
.B(n_762),
.C(n_763),
.Y(n_4596)
);

AOI21xp5_ASAP7_75t_L g4597 ( 
.A1(n_4582),
.A2(n_4578),
.B(n_4570),
.Y(n_4597)
);

AOI221xp5_ASAP7_75t_SL g4598 ( 
.A1(n_4577),
.A2(n_3954),
.B1(n_3975),
.B2(n_3953),
.C(n_3947),
.Y(n_4598)
);

AOI31xp33_ASAP7_75t_L g4599 ( 
.A1(n_4581),
.A2(n_4085),
.A3(n_4097),
.B(n_4093),
.Y(n_4599)
);

AOI22xp5_ASAP7_75t_L g4600 ( 
.A1(n_4560),
.A2(n_4053),
.B1(n_3981),
.B2(n_3991),
.Y(n_4600)
);

AOI322xp5_ASAP7_75t_L g4601 ( 
.A1(n_4560),
.A2(n_3975),
.A3(n_3981),
.B1(n_3991),
.B2(n_3998),
.C1(n_3996),
.C2(n_3999),
.Y(n_4601)
);

O2A1O1Ixp33_ASAP7_75t_SL g4602 ( 
.A1(n_4566),
.A2(n_4099),
.B(n_4112),
.C(n_4105),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_4560),
.B(n_3961),
.Y(n_4603)
);

OAI22xp5_ASAP7_75t_L g4604 ( 
.A1(n_4564),
.A2(n_4080),
.B1(n_4111),
.B2(n_4088),
.Y(n_4604)
);

XNOR2xp5_ASAP7_75t_L g4605 ( 
.A(n_4565),
.B(n_763),
.Y(n_4605)
);

AOI221xp5_ASAP7_75t_L g4606 ( 
.A1(n_4560),
.A2(n_3961),
.B1(n_4059),
.B2(n_4066),
.C(n_4058),
.Y(n_4606)
);

NOR2xp33_ASAP7_75t_SL g4607 ( 
.A(n_4584),
.B(n_4125),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4603),
.Y(n_4608)
);

AOI31xp33_ASAP7_75t_L g4609 ( 
.A1(n_4605),
.A2(n_766),
.A3(n_764),
.B(n_765),
.Y(n_4609)
);

AND2x2_ASAP7_75t_L g4610 ( 
.A(n_4585),
.B(n_3963),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4604),
.Y(n_4611)
);

NOR2xp33_ASAP7_75t_L g4612 ( 
.A(n_4593),
.B(n_767),
.Y(n_4612)
);

AOI22xp5_ASAP7_75t_L g4613 ( 
.A1(n_4600),
.A2(n_3918),
.B1(n_3968),
.B2(n_3967),
.Y(n_4613)
);

NOR2x1_ASAP7_75t_L g4614 ( 
.A(n_4597),
.B(n_3283),
.Y(n_4614)
);

NOR2xp67_ASAP7_75t_L g4615 ( 
.A(n_4590),
.B(n_767),
.Y(n_4615)
);

NOR2x1_ASAP7_75t_L g4616 ( 
.A(n_4595),
.B(n_768),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_4586),
.B(n_3973),
.Y(n_4617)
);

NOR2x1_ASAP7_75t_L g4618 ( 
.A(n_4587),
.B(n_768),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4599),
.Y(n_4619)
);

INVx2_ASAP7_75t_L g4620 ( 
.A(n_4594),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4602),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4592),
.Y(n_4622)
);

NAND2xp5_ASAP7_75t_L g4623 ( 
.A(n_4596),
.B(n_769),
.Y(n_4623)
);

NOR2x1_ASAP7_75t_L g4624 ( 
.A(n_4591),
.B(n_4601),
.Y(n_4624)
);

OAI221xp5_ASAP7_75t_L g4625 ( 
.A1(n_4612),
.A2(n_4618),
.B1(n_4624),
.B2(n_4607),
.C(n_4623),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4610),
.Y(n_4626)
);

AND2x2_ASAP7_75t_SL g4627 ( 
.A(n_4620),
.B(n_4588),
.Y(n_4627)
);

NAND4xp75_ASAP7_75t_L g4628 ( 
.A(n_4616),
.B(n_4598),
.C(n_4589),
.D(n_4606),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4608),
.Y(n_4629)
);

BUFx2_ASAP7_75t_L g4630 ( 
.A(n_4621),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4611),
.Y(n_4631)
);

CKINVDCx20_ASAP7_75t_R g4632 ( 
.A(n_4619),
.Y(n_4632)
);

HB1xp67_ASAP7_75t_L g4633 ( 
.A(n_4615),
.Y(n_4633)
);

XOR2xp5_ASAP7_75t_L g4634 ( 
.A(n_4622),
.B(n_769),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4609),
.Y(n_4635)
);

NAND4xp75_ASAP7_75t_L g4636 ( 
.A(n_4617),
.B(n_772),
.C(n_770),
.D(n_771),
.Y(n_4636)
);

NAND2xp33_ASAP7_75t_SL g4637 ( 
.A(n_4615),
.B(n_3447),
.Y(n_4637)
);

CKINVDCx16_ASAP7_75t_R g4638 ( 
.A(n_4632),
.Y(n_4638)
);

CKINVDCx20_ASAP7_75t_R g4639 ( 
.A(n_4634),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4626),
.Y(n_4640)
);

CKINVDCx5p33_ASAP7_75t_R g4641 ( 
.A(n_4630),
.Y(n_4641)
);

CKINVDCx20_ASAP7_75t_R g4642 ( 
.A(n_4635),
.Y(n_4642)
);

HB1xp67_ASAP7_75t_L g4643 ( 
.A(n_4629),
.Y(n_4643)
);

CKINVDCx5p33_ASAP7_75t_R g4644 ( 
.A(n_4631),
.Y(n_4644)
);

NOR2xp33_ASAP7_75t_L g4645 ( 
.A(n_4625),
.B(n_4614),
.Y(n_4645)
);

INVx2_ASAP7_75t_L g4646 ( 
.A(n_4638),
.Y(n_4646)
);

AOI22xp5_ASAP7_75t_L g4647 ( 
.A1(n_4642),
.A2(n_4625),
.B1(n_4636),
.B2(n_4628),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4641),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_4646),
.B(n_4627),
.Y(n_4649)
);

INVx2_ASAP7_75t_L g4650 ( 
.A(n_4648),
.Y(n_4650)
);

CKINVDCx20_ASAP7_75t_R g4651 ( 
.A(n_4647),
.Y(n_4651)
);

INVx2_ASAP7_75t_L g4652 ( 
.A(n_4650),
.Y(n_4652)
);

AOI22x1_ASAP7_75t_L g4653 ( 
.A1(n_4652),
.A2(n_4644),
.B1(n_4643),
.B2(n_4640),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_L g4654 ( 
.A(n_4653),
.B(n_4645),
.Y(n_4654)
);

AOI22xp33_ASAP7_75t_SL g4655 ( 
.A1(n_4654),
.A2(n_4651),
.B1(n_4639),
.B2(n_4649),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_L g4656 ( 
.A(n_4655),
.B(n_4633),
.Y(n_4656)
);

AOI31xp33_ASAP7_75t_L g4657 ( 
.A1(n_4656),
.A2(n_4637),
.A3(n_4613),
.B(n_774),
.Y(n_4657)
);


endmodule