module real_jpeg_1020_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_SL g12 ( 
.A(n_0),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_15),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_0),
.B(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g9 ( 
.A(n_1),
.Y(n_9)
);

OR2x4_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_1),
.B(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_4),
.B(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_18),
.Y(n_17)
);

NAND2x1_ASAP7_75t_SL g19 ( 
.A(n_4),
.B(n_18),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_9),
.Y(n_8)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_26),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_10),
.B1(n_20),
.B2(n_22),
.Y(n_7)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_9),
.B(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_13),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_12),
.B(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_12),
.B(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

OA21x2_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_17),
.B(n_19),
.Y(n_15)
);

OA21x2_ASAP7_75t_L g32 ( 
.A1(n_16),
.A2(n_33),
.B(n_34),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_19),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI211xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B(n_36),
.C(n_38),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);


endmodule