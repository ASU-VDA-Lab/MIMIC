module real_jpeg_25469_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_1),
.A2(n_51),
.B1(n_52),
.B2(n_58),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_1),
.A2(n_25),
.B1(n_29),
.B2(n_58),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_3),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_79),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_5),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_5),
.A2(n_51),
.B1(n_52),
.B2(n_79),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_5),
.A2(n_25),
.B1(n_29),
.B2(n_79),
.Y(n_145)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_61),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_9),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_9),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_9),
.A2(n_61),
.B1(n_93),
.B2(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_9),
.A2(n_25),
.B1(n_29),
.B2(n_61),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_10),
.A2(n_25),
.B1(n_29),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_10),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_11),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_11),
.B(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_11),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_11),
.B(n_52),
.C(n_54),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_96),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_11),
.B(n_77),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_96),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_11),
.B(n_25),
.C(n_85),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_11),
.A2(n_24),
.B(n_146),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_13),
.A2(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_14),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_121),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_119),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_101),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_18),
.B(n_101),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_72),
.B2(n_73),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_48),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.B1(n_31),
.B2(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_23),
.A2(n_158),
.B1(n_160),
.B2(n_162),
.Y(n_157)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_24),
.A2(n_28),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_24),
.B(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_24),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_25),
.A2(n_29),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_26),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_29),
.B(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_31),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI32xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.A3(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_38),
.B1(n_54),
.B2(n_55),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_67)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_38),
.B(n_114),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_41),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_93),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_65),
.C(n_68),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_56),
.B(n_59),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_52),
.B1(n_84),
.B2(n_85),
.Y(n_88)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_52),
.B(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_62),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_60),
.B(n_77),
.Y(n_131)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_63),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_71),
.A2(n_159),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_90),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_81),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_86),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_83),
.A2(n_86),
.B(n_127),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_83),
.B(n_96),
.Y(n_167)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_109),
.B1(n_111),
.B2(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_95),
.B(n_98),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_96),
.B(n_161),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.C(n_112),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_103),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_112),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B(n_110),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_110),
.B(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_113),
.B(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_135),
.B(n_183),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_132),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_123),
.B(n_132),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.C(n_128),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_124),
.B(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_125),
.A2(n_128),
.B1(n_129),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_177),
.B(n_182),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_155),
.B(n_176),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_149),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_149),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_144),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_143),
.C(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_165),
.B(n_175),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_163),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_170),
.B(n_174),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_181),
.Y(n_182)
);


endmodule