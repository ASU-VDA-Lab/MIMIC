module fake_jpeg_22141_n_163 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_163);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_15),
.Y(n_54)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_0),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_24),
.Y(n_45)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_57),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_31),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_17),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_15),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_65),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_60),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_16),
.Y(n_62)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_31),
.B1(n_29),
.B2(n_25),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_68),
.B1(n_27),
.B2(n_22),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_42),
.B1(n_29),
.B2(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_35),
.A2(n_28),
.B1(n_27),
.B2(n_22),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_70),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_93)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_75),
.Y(n_98)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_80),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2x1_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_0),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_83),
.B(n_85),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_1),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_89),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_1),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_91),
.Y(n_104)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_16),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_82),
.B(n_21),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_52),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_100),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_49),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_103),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_105),
.B(n_108),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_74),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_85),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_55),
.B1(n_65),
.B2(n_51),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_80),
.B1(n_90),
.B2(n_81),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_60),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_51),
.B1(n_69),
.B2(n_71),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_84),
.B1(n_72),
.B2(n_58),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_87),
.B1(n_78),
.B2(n_76),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_117),
.B(n_63),
.Y(n_135)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_121),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_85),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_123),
.C(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_100),
.C(n_106),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_125),
.B(n_77),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_133),
.C(n_137),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_99),
.B(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_130),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_92),
.A3(n_104),
.B1(n_111),
.B2(n_110),
.C1(n_103),
.C2(n_102),
.Y(n_132)
);

OAI322xp33_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_114),
.A3(n_119),
.B1(n_125),
.B2(n_19),
.C1(n_120),
.C2(n_121),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_59),
.C(n_97),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_136),
.B(n_113),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_61),
.C(n_63),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_134),
.B(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_112),
.B1(n_119),
.B2(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_143),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_123),
.C(n_115),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_133),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_144),
.A2(n_136),
.B1(n_137),
.B2(n_56),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_89),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_75),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_151),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_150),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_152),
.B(n_144),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_155),
.C(n_149),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_141),
.A3(n_142),
.B1(n_138),
.B2(n_11),
.C1(n_13),
.C2(n_8),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_156),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_1),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_138),
.C(n_147),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_159),
.B1(n_2),
.B2(n_4),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_153),
.A2(n_151),
.B(n_12),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_160),
.A2(n_161),
.B(n_5),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_6),
.Y(n_163)
);


endmodule