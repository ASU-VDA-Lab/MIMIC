module fake_jpeg_13269_n_168 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_35),
.B(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_36),
.B(n_38),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g38 ( 
.A(n_12),
.B(n_0),
.C(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_6),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_17),
.Y(n_62)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_13),
.B(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_53),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_16),
.B(n_4),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_58),
.Y(n_83)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_56),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_12),
.B(n_5),
.C(n_6),
.Y(n_57)
);

FAx1_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_5),
.CI(n_31),
.CON(n_61),
.SN(n_61)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_18),
.B1(n_23),
.B2(n_31),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_59),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_62),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_18),
.B(n_23),
.C(n_31),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_63),
.A2(n_77),
.B(n_65),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_5),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_58),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_21),
.B1(n_24),
.B2(n_17),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_87),
.B(n_82),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_49),
.B1(n_47),
.B2(n_43),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_21),
.B1(n_24),
.B2(n_38),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_53),
.B1(n_54),
.B2(n_19),
.Y(n_71)
);

AOI32xp33_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_54),
.A3(n_38),
.B1(n_35),
.B2(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_50),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_95),
.Y(n_129)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_83),
.B1(n_80),
.B2(n_88),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_110),
.B1(n_102),
.B2(n_99),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_106),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_72),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_104),
.Y(n_127)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

NOR2x1_ASAP7_75t_SL g105 ( 
.A(n_63),
.B(n_59),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_80),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_72),
.A2(n_74),
.B1(n_63),
.B2(n_79),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_101),
.B1(n_109),
.B2(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_111),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_100),
.B(n_108),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_65),
.B1(n_70),
.B2(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_62),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_92),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_98),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_116),
.B(n_125),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_119),
.A2(n_126),
.B(n_113),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_120),
.A2(n_122),
.B1(n_125),
.B2(n_103),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_91),
.B(n_101),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_93),
.B1(n_111),
.B2(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_112),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_96),
.B1(n_106),
.B2(n_92),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_90),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_95),
.B1(n_120),
.B2(n_122),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_137),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_115),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_114),
.A3(n_127),
.B1(n_129),
.B2(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_139),
.B(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_116),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_140),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_129),
.C(n_121),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_146),
.C(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_148),
.B(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_151),
.A2(n_155),
.B(n_145),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_153),
.B(n_137),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_143),
.A2(n_134),
.B1(n_135),
.B2(n_119),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_158),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_151),
.C(n_155),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_150),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_158),
.B(n_149),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_149),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_160),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_166),
.C(n_144),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_144),
.Y(n_168)
);


endmodule