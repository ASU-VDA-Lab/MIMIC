module real_jpeg_22915_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_249;
wire n_286;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_200;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_2),
.A2(n_20),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_2),
.A2(n_30),
.B1(n_32),
.B2(n_59),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_2),
.A2(n_51),
.B1(n_53),
.B2(n_59),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_2),
.A2(n_59),
.B1(n_72),
.B2(n_73),
.Y(n_196)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_6),
.A2(n_18),
.B1(n_21),
.B2(n_24),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_6),
.A2(n_24),
.B1(n_30),
.B2(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_24),
.B1(n_51),
.B2(n_53),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_6),
.A2(n_24),
.B1(n_72),
.B2(n_73),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_18),
.B1(n_21),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_7),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_7),
.A2(n_34),
.B1(n_51),
.B2(n_53),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_7),
.A2(n_34),
.B1(n_72),
.B2(n_73),
.Y(n_90)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_8),
.A2(n_9),
.B1(n_18),
.B2(n_41),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_9),
.A2(n_41),
.B1(n_51),
.B2(n_53),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_9),
.A2(n_30),
.B1(n_32),
.B2(n_41),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_9),
.A2(n_41),
.B1(n_72),
.B2(n_73),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_9),
.B(n_28),
.C(n_32),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_9),
.B(n_29),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_9),
.B(n_48),
.C(n_51),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_9),
.B(n_69),
.C(n_72),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_9),
.B(n_11),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_9),
.B(n_105),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_9),
.B(n_62),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_11),
.Y(n_89)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_11),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_11),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_77),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_75),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_35),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_15),
.B(n_35),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_25),
.B1(n_29),
.B2(n_33),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_17),
.A2(n_38),
.B(n_39),
.Y(n_37)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_19),
.B(n_192),
.Y(n_191)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_25),
.A2(n_29),
.B1(n_40),
.B2(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_25),
.B(n_29),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

AO22x1_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_29)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_30),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_32),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_32),
.B(n_225),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_36),
.B(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_36),
.B(n_293),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_42),
.CI(n_54),
.CON(n_36),
.SN(n_36)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_38),
.A2(n_39),
.B(n_57),
.Y(n_114)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_46),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_45),
.A2(n_50),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_46),
.A2(n_62),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_46),
.B(n_110),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OA22x2_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_50),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_50),
.A2(n_109),
.B(n_120),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_53),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_51),
.B(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.C(n_63),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_SL g127 ( 
.A(n_55),
.B(n_128),
.C(n_136),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_55),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_55),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_55),
.A2(n_136),
.B1(n_137),
.B2(n_150),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_55),
.A2(n_107),
.B1(n_150),
.B2(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_55),
.B(n_107),
.C(n_189),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_60),
.A2(n_63),
.B1(n_117),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_60),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_63),
.A2(n_117),
.B1(n_118),
.B2(n_121),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_63),
.B(n_113),
.C(n_118),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_74),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_65),
.B(n_95),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_67),
.A2(n_95),
.B1(n_105),
.B2(n_135),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_71),
.A2(n_94),
.B(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_72),
.B(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_292),
.B(n_294),
.Y(n_77)
);

OAI211xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_138),
.B(n_152),
.C(n_291),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_122),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_80),
.B(n_122),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_100),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_81),
.B(n_102),
.C(n_111),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_91),
.B(n_96),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_82),
.A2(n_96),
.B1(n_97),
.B2(n_125),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_82),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_82),
.A2(n_92),
.B1(n_125),
.B2(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_90),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_84),
.B(n_197),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_85),
.A2(n_90),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_85),
.B(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_85),
.Y(n_195)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_91),
.B(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_92),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_111),
.B2(n_112),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_103),
.B(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_107),
.B(n_209),
.C(n_211),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_107),
.A2(n_199),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_110),
.Y(n_172)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_114),
.B1(n_146),
.B2(n_151),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_113),
.B(n_136),
.C(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_113),
.A2(n_114),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_113),
.A2(n_114),
.B1(n_171),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_162),
.C(n_171),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_114),
.B(n_142),
.C(n_146),
.Y(n_293)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_118),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.C(n_127),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_126),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_129),
.A2(n_133),
.B1(n_134),
.B2(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_129),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_130),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_133),
.A2(n_134),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_133),
.A2(n_134),
.B1(n_222),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_134),
.B(n_216),
.C(n_222),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_134),
.B(n_194),
.C(n_253),
.Y(n_257)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_136),
.A2(n_137),
.B1(n_185),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_136),
.A2(n_137),
.B1(n_169),
.B2(n_182),
.Y(n_259)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_137),
.B(n_169),
.C(n_260),
.Y(n_263)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_153),
.C(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_140),
.B(n_141),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_175),
.B(n_290),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_173),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_156),
.B(n_173),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.C(n_161),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_157),
.B(n_159),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_161),
.B(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_162),
.A2(n_163),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_169),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_164),
.Y(n_183)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_167),
.A2(n_196),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_169),
.A2(n_182),
.B1(n_237),
.B2(n_239),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_169),
.B(n_239),
.Y(n_249)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_171),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_285),
.B(n_289),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_212),
.B(n_271),
.C(n_284),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_201),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_178),
.B(n_201),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_188),
.B2(n_200),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_181),
.B(n_187),
.C(n_200),
.Y(n_272)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_198),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_193),
.A2(n_194),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_194),
.B(n_245),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.C(n_208),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_202),
.A2(n_203),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_208),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_211),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_209),
.B(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_211),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_270),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_231),
.B(n_269),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_228),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_215),
.B(n_228),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_216),
.A2(n_217),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_221),
.B(n_236),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_262),
.B(n_268),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_256),
.B(n_261),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_248),
.B(n_255),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_240),
.B(n_247),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_237),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_244),
.B(n_246),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_249),
.B(n_250),
.Y(n_255)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_253),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_258),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_263),
.B(n_264),
.Y(n_268)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_273),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_283),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_280),
.B2(n_281),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_281),
.C(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_287),
.Y(n_289)
);


endmodule