module fake_jpeg_17205_n_296 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_26),
.C(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_26),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_51),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_29),
.B1(n_30),
.B2(n_25),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_29),
.B1(n_22),
.B2(n_24),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_45),
.B1(n_49),
.B2(n_53),
.Y(n_73)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_29),
.B1(n_32),
.B2(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_21),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_16),
.B1(n_17),
.B2(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_57),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_16),
.B1(n_17),
.B2(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_26),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_16),
.B1(n_19),
.B2(n_30),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_21),
.B1(n_19),
.B2(n_30),
.Y(n_74)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_65),
.A2(n_68),
.B1(n_74),
.B2(n_86),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_52),
.B(n_57),
.C(n_48),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_69),
.B1(n_43),
.B2(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_33),
.B1(n_35),
.B2(n_34),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_24),
.B1(n_23),
.B2(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_23),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_77),
.B(n_81),
.C(n_58),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_83),
.Y(n_95)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_33),
.CI(n_38),
.CON(n_77),
.SN(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_78),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_24),
.B(n_28),
.C(n_21),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_37),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_37),
.C(n_35),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_42),
.A2(n_28),
.B1(n_38),
.B2(n_22),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_89),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_51),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_108),
.C(n_117),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_98),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_48),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_56),
.B1(n_46),
.B2(n_47),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_64),
.B(n_61),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_101),
.B(n_80),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_61),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_87),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_59),
.B1(n_47),
.B2(n_35),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_111),
.B1(n_115),
.B2(n_88),
.Y(n_121)
);

AO21x2_ASAP7_75t_L g107 ( 
.A1(n_71),
.A2(n_35),
.B(n_34),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_60),
.B1(n_75),
.B2(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_59),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_113),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_59),
.B1(n_34),
.B2(n_56),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_34),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_27),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_27),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_73),
.A2(n_46),
.B1(n_22),
.B2(n_37),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_27),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_124),
.B1(n_131),
.B2(n_133),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_114),
.A2(n_67),
.B(n_79),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_122),
.A2(n_123),
.B(n_130),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_79),
.B(n_73),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_65),
.B1(n_79),
.B2(n_68),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_109),
.B1(n_115),
.B2(n_98),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_80),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_138),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_107),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_137),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_69),
.B1(n_74),
.B2(n_81),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_132),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_116),
.B(n_106),
.C(n_96),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_117),
.B(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_135),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_76),
.B(n_64),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_95),
.B(n_107),
.Y(n_147)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_82),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_95),
.B(n_22),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_87),
.B1(n_78),
.B2(n_18),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_167)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_91),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_1),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_147),
.A2(n_148),
.B1(n_167),
.B2(n_120),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_93),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_150),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_108),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_157),
.C(n_164),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_134),
.B1(n_121),
.B2(n_130),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_111),
.C(n_103),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_154),
.B(n_156),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_92),
.C(n_78),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_18),
.B(n_27),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_163),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_166),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_27),
.B(n_2),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_91),
.C(n_9),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_9),
.Y(n_165)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_176),
.CI(n_14),
.CON(n_197),
.SN(n_197)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_14),
.C(n_13),
.Y(n_166)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_175),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_14),
.C(n_12),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_11),
.Y(n_203)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_151),
.A2(n_129),
.B1(n_145),
.B2(n_134),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_184),
.B1(n_185),
.B2(n_191),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_181),
.B(n_186),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_134),
.A3(n_146),
.B1(n_143),
.B2(n_140),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_151),
.A2(n_134),
.B1(n_136),
.B2(n_127),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_155),
.B(n_138),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_162),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_189),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_193),
.B1(n_194),
.B2(n_200),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_149),
.A2(n_157),
.B1(n_164),
.B2(n_177),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_118),
.B1(n_135),
.B2(n_132),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_148),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_15),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_147),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_15),
.C(n_12),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_203),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_168),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_156),
.B(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_160),
.Y(n_206)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_152),
.C(n_150),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_217),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_173),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_210),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_195),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_165),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_216),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_166),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_158),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_163),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_221),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_176),
.C(n_171),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_224),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_169),
.B(n_175),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_220),
.A2(n_182),
.B1(n_188),
.B2(n_185),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_167),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_170),
.C(n_3),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_223),
.B(n_191),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_228),
.B(n_223),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_215),
.B(n_197),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_183),
.B1(n_184),
.B2(n_180),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_231),
.A2(n_236),
.B1(n_213),
.B2(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_239),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_222),
.B(n_203),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_234),
.B(n_205),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_224),
.A2(n_194),
.B1(n_179),
.B2(n_197),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_209),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_179),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_213),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_208),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_219),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_249),
.C(n_250),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_227),
.B1(n_244),
.B2(n_235),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_247),
.A2(n_231),
.B1(n_240),
.B2(n_237),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_217),
.C(n_226),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_253),
.C(n_254),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_252),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_220),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_228),
.B(n_212),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_10),
.C(n_11),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_225),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_258),
.A2(n_242),
.B(n_232),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_264),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_243),
.B(n_205),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_265),
.B(n_266),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_243),
.Y(n_264)
);

NOR3xp33_ASAP7_75t_SL g265 ( 
.A(n_251),
.B(n_236),
.C(n_218),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_210),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_216),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_267),
.A2(n_1),
.B(n_4),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_270),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_260),
.A2(n_253),
.B(n_248),
.Y(n_273)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_246),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_275),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_265),
.A2(n_250),
.B(n_255),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_270),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_278),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_259),
.B(n_263),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_283),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_4),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_286),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_5),
.C(n_6),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_288),
.A2(n_289),
.B1(n_287),
.B2(n_7),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_277),
.B(n_274),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_285),
.B(n_283),
.C(n_7),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_292),
.C(n_5),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_5),
.C(n_6),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_295),
.Y(n_296)
);


endmodule