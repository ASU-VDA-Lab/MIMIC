module fake_jpeg_14076_n_531 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_531);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_531;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_12),
.B(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_60),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_61),
.Y(n_191)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_62),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_10),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_63),
.B(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_10),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_83),
.Y(n_124)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_65),
.Y(n_200)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_66),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g68 ( 
.A(n_22),
.Y(n_68)
);

CKINVDCx6p67_ASAP7_75t_R g143 ( 
.A(n_68),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_10),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_74),
.B(n_81),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_76),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_77),
.Y(n_177)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_80),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_10),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_21),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_89),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_28),
.B(n_9),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_90),
.B(n_93),
.Y(n_134)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_28),
.B(n_9),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_94),
.Y(n_193)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_95),
.Y(n_197)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_96),
.Y(n_198)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_97),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_30),
.B(n_17),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_103),
.Y(n_202)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_18),
.Y(n_104)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_30),
.B(n_9),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_106),
.B(n_109),
.Y(n_145)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_107),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_39),
.B(n_34),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_18),
.Y(n_117)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_39),
.B(n_8),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_118),
.B(n_13),
.Y(n_186)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_32),
.Y(n_119)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_32),
.Y(n_120)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_18),
.Y(n_122)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_31),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_34),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_47),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_128),
.B(n_131),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_130),
.B(n_42),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_47),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_71),
.A2(n_23),
.B1(n_32),
.B2(n_54),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_135),
.A2(n_139),
.B1(n_146),
.B2(n_165),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_59),
.A2(n_56),
.B1(n_44),
.B2(n_46),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_137),
.A2(n_21),
.B1(n_1),
.B2(n_0),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_65),
.A2(n_44),
.B1(n_46),
.B2(n_56),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_138),
.A2(n_70),
.B1(n_113),
.B2(n_112),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_84),
.A2(n_54),
.B1(n_44),
.B2(n_46),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_54),
.B1(n_42),
.B2(n_18),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_55),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_147),
.B(n_152),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_97),
.B(n_55),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_48),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_154),
.B(n_160),
.Y(n_214)
);

BUFx2_ASAP7_75t_R g158 ( 
.A(n_62),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_158),
.B(n_114),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_69),
.B(n_48),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_76),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_68),
.B(n_41),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_170),
.B(n_173),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_80),
.B(n_45),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_85),
.B(n_45),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_175),
.B(n_186),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_121),
.A2(n_42),
.B1(n_38),
.B2(n_35),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_176),
.A2(n_180),
.B1(n_0),
.B2(n_1),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_116),
.A2(n_42),
.B1(n_35),
.B2(n_2),
.Y(n_180)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_60),
.Y(n_199)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_61),
.Y(n_203)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx4_ASAP7_75t_SL g307 ( 
.A(n_205),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_206),
.B(n_212),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_133),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_207),
.B(n_219),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_129),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_208),
.Y(n_282)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_209),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_149),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_210),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_211),
.A2(n_228),
.B1(n_162),
.B2(n_177),
.Y(n_292)
);

AO22x1_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_72),
.B1(n_110),
.B2(n_108),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_215),
.Y(n_284)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_216),
.Y(n_300)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_144),
.Y(n_217)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_217),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_125),
.A2(n_16),
.B(n_15),
.C(n_3),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_172),
.Y(n_220)
);

BUFx24_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_221),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_222),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_163),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_153),
.Y(n_227)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_227),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_138),
.A2(n_103),
.B1(n_99),
.B2(n_89),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_229),
.Y(n_273)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_230),
.Y(n_318)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_231),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_135),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_232),
.B(n_251),
.Y(n_289)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_233),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_234),
.Y(n_285)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_235),
.Y(n_294)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_236),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_124),
.B(n_145),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_238),
.B(n_247),
.Y(n_312)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_167),
.Y(n_239)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_239),
.Y(n_323)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_241),
.Y(n_286)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_140),
.Y(n_242)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_242),
.Y(n_308)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_140),
.Y(n_244)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_244),
.Y(n_320)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_171),
.Y(n_245)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_245),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_134),
.B(n_77),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_153),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_143),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_248),
.B(n_250),
.Y(n_322)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_197),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_249),
.Y(n_303)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_127),
.B(n_67),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_196),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_253),
.Y(n_291)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

AO22x1_ASAP7_75t_SL g254 ( 
.A1(n_136),
.A2(n_0),
.B1(n_1),
.B2(n_21),
.Y(n_254)
);

AO22x1_ASAP7_75t_SL g314 ( 
.A1(n_254),
.A2(n_164),
.B1(n_202),
.B2(n_204),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_141),
.B(n_11),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_256),
.B(n_258),
.Y(n_315)
);

AND2x2_ASAP7_75t_SL g257 ( 
.A(n_148),
.B(n_0),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_257),
.B(n_132),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_159),
.B(n_168),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_166),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_259),
.B(n_260),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_126),
.Y(n_260)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_191),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_261),
.B(n_262),
.Y(n_316)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_196),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_183),
.A2(n_21),
.B1(n_8),
.B2(n_3),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_266),
.B1(n_180),
.B2(n_139),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_143),
.B(n_14),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_264),
.B(n_265),
.Y(n_319)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_192),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_161),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_267),
.Y(n_279)
);

INVx3_ASAP7_75t_SL g268 ( 
.A(n_142),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_268),
.A2(n_270),
.B1(n_271),
.B2(n_182),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_143),
.B(n_155),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_272),
.Y(n_275)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_150),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_169),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_126),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_281),
.A2(n_317),
.B(n_257),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_205),
.A2(n_146),
.B(n_176),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_290),
.A2(n_245),
.B(n_250),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_292),
.A2(n_310),
.B1(n_266),
.B2(n_237),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_265),
.B1(n_259),
.B2(n_234),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_232),
.A2(n_156),
.B1(n_157),
.B2(n_192),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_246),
.A2(n_202),
.B1(n_204),
.B2(n_187),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_298),
.A2(n_222),
.B(n_223),
.Y(n_332)
);

XNOR2x1_ASAP7_75t_L g333 ( 
.A(n_301),
.B(n_257),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_251),
.A2(n_142),
.B1(n_177),
.B2(n_162),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_254),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_225),
.A2(n_182),
.B(n_200),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_237),
.A2(n_187),
.B1(n_183),
.B2(n_164),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_330),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_289),
.A2(n_271),
.B1(n_214),
.B2(n_255),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_226),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_328),
.B(n_341),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_292),
.A2(n_263),
.B1(n_254),
.B2(n_212),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_290),
.A2(n_191),
.B1(n_151),
.B2(n_200),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_339),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_332),
.A2(n_285),
.B1(n_293),
.B2(n_313),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_333),
.B(n_276),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_276),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_347),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_304),
.A2(n_219),
.B(n_208),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_335),
.A2(n_336),
.B(n_351),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_288),
.A2(n_268),
.B1(n_213),
.B2(n_233),
.Y(n_336)
);

AOI32xp33_ASAP7_75t_L g337 ( 
.A1(n_288),
.A2(n_188),
.A3(n_221),
.B1(n_240),
.B2(n_242),
.Y(n_337)
);

AOI32xp33_ASAP7_75t_L g375 ( 
.A1(n_337),
.A2(n_277),
.A3(n_274),
.B1(n_307),
.B2(n_276),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_315),
.B(n_229),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_281),
.B(n_253),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_342),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_343),
.A2(n_349),
.B1(n_298),
.B2(n_277),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_344),
.A2(n_332),
.B(n_338),
.Y(n_392)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_306),
.Y(n_345)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_345),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_322),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_287),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_295),
.A2(n_151),
.B1(n_231),
.B2(n_224),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_281),
.B(n_216),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_274),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_302),
.A2(n_260),
.B(n_220),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_287),
.Y(n_352)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_352),
.Y(n_381)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_316),
.Y(n_353)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_280),
.Y(n_354)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_301),
.B(n_244),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_357),
.C(n_329),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_314),
.A2(n_218),
.B1(n_261),
.B2(n_227),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_356),
.B(n_358),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_281),
.A2(n_275),
.B(n_319),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_357),
.A2(n_282),
.B(n_307),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_314),
.A2(n_247),
.B1(n_188),
.B2(n_0),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_317),
.B(n_1),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_359),
.B(n_360),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_310),
.A2(n_188),
.B1(n_8),
.B2(n_15),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_309),
.Y(n_361)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_361),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_275),
.B(n_291),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_362),
.B(n_364),
.Y(n_376)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_280),
.Y(n_363)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_363),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_279),
.B(n_6),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_365),
.A2(n_356),
.B1(n_358),
.B2(n_346),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_367),
.B(n_385),
.C(n_388),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_278),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_368),
.B(n_378),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_362),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_371),
.B(n_294),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_375),
.A2(n_396),
.B1(n_331),
.B2(n_340),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_382),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_333),
.B(n_311),
.C(n_318),
.Y(n_385)
);

AO22x1_ASAP7_75t_L g386 ( 
.A1(n_335),
.A2(n_284),
.B1(n_323),
.B2(n_286),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_386),
.B(n_394),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_333),
.B(n_305),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_391),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_344),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_347),
.B(n_299),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_325),
.A2(n_309),
.B1(n_324),
.B2(n_294),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_397),
.A2(n_406),
.B1(n_411),
.B2(n_412),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_353),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_399),
.B(n_402),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_401),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_328),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_374),
.A2(n_343),
.B1(n_349),
.B2(n_351),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_403),
.A2(n_404),
.B1(n_408),
.B2(n_414),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_374),
.A2(n_351),
.B1(n_359),
.B2(n_326),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_339),
.Y(n_407)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_407),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_366),
.A2(n_341),
.B1(n_350),
.B2(n_330),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_327),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_409),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_336),
.C(n_342),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_419),
.C(n_423),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_366),
.A2(n_360),
.B1(n_337),
.B2(n_334),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_389),
.A2(n_361),
.B1(n_345),
.B2(n_354),
.Y(n_412)
);

BUFx24_ASAP7_75t_SL g413 ( 
.A(n_395),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_413),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_389),
.A2(n_364),
.B1(n_361),
.B2(n_363),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_367),
.B(n_286),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_415),
.B(n_398),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_387),
.A2(n_352),
.B1(n_348),
.B2(n_293),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_416),
.A2(n_418),
.B1(n_372),
.B2(n_384),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_387),
.A2(n_313),
.B1(n_285),
.B2(n_324),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_368),
.B(n_303),
.C(n_308),
.Y(n_419)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_421),
.Y(n_428)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_372),
.Y(n_422)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_422),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_373),
.B(n_378),
.C(n_385),
.Y(n_423)
);

MAJx2_ASAP7_75t_L g424 ( 
.A(n_376),
.B(n_299),
.C(n_273),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_424),
.B(n_386),
.Y(n_441)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_425),
.Y(n_451)
);

AOI331xp33_ASAP7_75t_L g429 ( 
.A1(n_420),
.A2(n_386),
.A3(n_395),
.B1(n_379),
.B2(n_380),
.B3(n_370),
.C1(n_376),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_429),
.B(n_420),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_370),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_439),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_404),
.A2(n_403),
.B1(n_408),
.B2(n_417),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_421),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_438),
.B(n_407),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_405),
.B(n_379),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_441),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_417),
.A2(n_365),
.B1(n_396),
.B2(n_375),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_422),
.Y(n_443)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_414),
.A2(n_392),
.B1(n_390),
.B2(n_393),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_398),
.B(n_382),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_445),
.B(n_446),
.C(n_447),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_415),
.B(n_393),
.C(n_384),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_377),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_410),
.B(n_377),
.C(n_381),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_412),
.C(n_416),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_449),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_450),
.B(n_463),
.Y(n_477)
);

AO21x1_ASAP7_75t_L g483 ( 
.A1(n_452),
.A2(n_426),
.B(n_427),
.Y(n_483)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_455),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_430),
.A2(n_401),
.B(n_400),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_456),
.A2(n_458),
.B(n_428),
.Y(n_481)
);

FAx1_ASAP7_75t_SL g459 ( 
.A(n_429),
.B(n_400),
.CI(n_419),
.CON(n_459),
.SN(n_459)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_460),
.Y(n_471)
);

FAx1_ASAP7_75t_SL g460 ( 
.A(n_445),
.B(n_400),
.CI(n_424),
.CON(n_460),
.SN(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_433),
.A2(n_397),
.B1(n_411),
.B2(n_424),
.Y(n_461)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_461),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_369),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_465),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_434),
.C(n_447),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_381),
.C(n_418),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_467),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_436),
.B(n_390),
.C(n_320),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_438),
.Y(n_474)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_474),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_462),
.Y(n_476)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_476),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_458),
.A2(n_435),
.B(n_442),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_478),
.B(n_480),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_426),
.Y(n_479)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_479),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_454),
.Y(n_480)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_481),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_454),
.B(n_448),
.Y(n_482)
);

XNOR2x1_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_453),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_483),
.A2(n_484),
.B1(n_444),
.B2(n_427),
.Y(n_494)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_457),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_480),
.C(n_472),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_473),
.A2(n_469),
.B1(n_428),
.B2(n_464),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_490),
.A2(n_495),
.B1(n_496),
.B2(n_492),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_466),
.C(n_467),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_491),
.B(n_493),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_453),
.C(n_446),
.Y(n_493)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_494),
.Y(n_504)
);

OAI221xp5_ASAP7_75t_L g495 ( 
.A1(n_470),
.A2(n_459),
.B1(n_460),
.B2(n_456),
.C(n_431),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_473),
.A2(n_471),
.B1(n_470),
.B2(n_474),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_498),
.A2(n_503),
.B1(n_443),
.B2(n_437),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_485),
.A2(n_481),
.B1(n_479),
.B2(n_471),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_499),
.A2(n_502),
.B1(n_506),
.B2(n_460),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_440),
.C(n_484),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_491),
.B(n_472),
.C(n_482),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_501),
.A2(n_468),
.B(n_441),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_488),
.A2(n_483),
.B1(n_477),
.B2(n_425),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_496),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_431),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_505),
.B(n_486),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_493),
.A2(n_459),
.B1(n_478),
.B2(n_461),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_507),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_487),
.C(n_489),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_510),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_509),
.B(n_514),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_487),
.C(n_468),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_511),
.A2(n_512),
.B(n_513),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_499),
.B(n_437),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_504),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_516),
.A2(n_519),
.B(n_369),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_508),
.A2(n_503),
.B(n_500),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_517),
.A2(n_506),
.B(n_502),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_521),
.A2(n_522),
.B(n_523),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_518),
.A2(n_369),
.B(n_300),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_515),
.C(n_320),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_300),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_525),
.A2(n_283),
.B(n_303),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_527),
.B(n_526),
.C(n_283),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_308),
.B(n_273),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_6),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_6),
.B(n_16),
.Y(n_531)
);


endmodule