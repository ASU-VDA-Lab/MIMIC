module fake_netlist_1_8584_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVxp67_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_3), .B(n_7), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_5), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_8), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_6), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_10), .B(n_0), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_11), .B(n_0), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_11), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_11), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_15), .Y(n_21) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_17), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_18), .A2(n_10), .B1(n_12), .B2(n_14), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_18), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_24), .B(n_18), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_23), .B(n_18), .Y(n_26) );
NAND3xp33_ASAP7_75t_L g27 ( .A(n_23), .B(n_13), .C(n_16), .Y(n_27) );
OAI221xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_14), .B1(n_15), .B2(n_20), .C(n_19), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_22), .B1(n_12), .B2(n_15), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_25), .B1(n_12), .B2(n_21), .Y(n_30) );
AOI21xp33_ASAP7_75t_SL g31 ( .A1(n_29), .A2(n_0), .B(n_1), .Y(n_31) );
OAI321xp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_21), .A3(n_25), .B1(n_1), .B2(n_2), .C(n_4), .Y(n_32) );
A2O1A1Ixp33_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_12), .B(n_2), .C(n_1), .Y(n_33) );
INVx2_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
AOI22xp33_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_33), .B1(n_8), .B2(n_9), .Y(n_35) );
endmodule