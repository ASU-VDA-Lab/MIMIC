module fake_jpeg_14785_n_124 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_124);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_4),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_5),
.Y(n_15)
);

AND2x2_ASAP7_75t_SL g16 ( 
.A(n_6),
.B(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx9p33_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_13),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_1),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_2),
.C(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_21),
.B(n_2),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_6),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_36),
.B(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_19),
.B(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_10),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_24),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_18),
.B(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_18),
.B(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_46),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_20),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_29),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_25),
.B1(n_17),
.B2(n_22),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_67),
.B1(n_51),
.B2(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_14),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_22),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_29),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_35),
.A2(n_23),
.B1(n_34),
.B2(n_39),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_78),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_32),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_68),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_34),
.B1(n_39),
.B2(n_59),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_57),
.B(n_55),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_79),
.B(n_65),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_46),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_87),
.B(n_69),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_55),
.B(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_53),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_94),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_47),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_80),
.B(n_72),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_78),
.B1(n_76),
.B2(n_72),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_102),
.B(n_104),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_83),
.C(n_74),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_89),
.C(n_85),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_80),
.B1(n_73),
.B2(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_92),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_88),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_109),
.C(n_110),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_91),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_100),
.B(n_94),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_112),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_93),
.C(n_87),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_103),
.B(n_99),
.C(n_106),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_116),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_106),
.B(n_47),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_117),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_111),
.C(n_47),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_119),
.C(n_114),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_121),
.Y(n_124)
);


endmodule