module fake_aes_12611_n_722 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_39, n_722);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_39;
output n_722;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g94 ( .A(n_12), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_14), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_32), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_52), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_24), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_53), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_73), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_93), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_80), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_46), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_70), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_71), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_82), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_14), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_72), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_47), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_69), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_63), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_78), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_85), .Y(n_113) );
BUFx10_ASAP7_75t_L g114 ( .A(n_13), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_37), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_2), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_40), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_35), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_65), .Y(n_119) );
INVxp33_ASAP7_75t_L g120 ( .A(n_48), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_75), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_91), .Y(n_122) );
CKINVDCx14_ASAP7_75t_R g123 ( .A(n_87), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_3), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_60), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_76), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_30), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_68), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_10), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_27), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_28), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_15), .B(n_83), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_105), .Y(n_133) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_110), .A2(n_42), .B(n_90), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_119), .B(n_0), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_130), .B(n_0), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_129), .B(n_1), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_112), .Y(n_138) );
NOR2xp33_ASAP7_75t_SL g139 ( .A(n_109), .B(n_20), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_95), .B(n_1), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_130), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_130), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_105), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_130), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_130), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_129), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_95), .B(n_2), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_110), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_96), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_94), .B(n_3), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_116), .B(n_4), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_98), .Y(n_152) );
OR2x2_ASAP7_75t_L g153 ( .A(n_135), .B(n_111), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_137), .Y(n_154) );
INVx2_ASAP7_75t_SL g155 ( .A(n_133), .Y(n_155) );
OR2x2_ASAP7_75t_L g156 ( .A(n_135), .B(n_115), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_133), .B(n_99), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_142), .Y(n_158) );
BUFx6f_ASAP7_75t_SL g159 ( .A(n_137), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_142), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_143), .B(n_123), .Y(n_161) );
INVxp67_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_148), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_143), .B(n_100), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_148), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_137), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_149), .B(n_103), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_137), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_149), .B(n_102), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_150), .Y(n_171) );
INVx4_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_142), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_134), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_152), .B(n_104), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
BUFx10_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_150), .A2(n_124), .B1(n_107), .B2(n_108), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_152), .B(n_102), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_141), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_138), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_163), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_162), .B(n_139), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_162), .A2(n_139), .B1(n_151), .B2(n_147), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_165), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_165), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_161), .B(n_146), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_153), .A2(n_146), .B(n_136), .C(n_108), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_161), .B(n_114), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_177), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_180), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_161), .B(n_118), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_167), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_155), .B(n_118), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_153), .A2(n_113), .B(n_117), .C(n_106), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_153), .B(n_156), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_156), .B(n_121), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_156), .B(n_121), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_172), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_155), .B(n_122), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_180), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_178), .B(n_114), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_155), .B(n_122), .Y(n_206) );
AND2x6_ASAP7_75t_SL g207 ( .A(n_183), .B(n_132), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_167), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_172), .B(n_125), .Y(n_209) );
NOR2x1p5_ASAP7_75t_L g210 ( .A(n_168), .B(n_116), .Y(n_210) );
AND2x6_ASAP7_75t_SL g211 ( .A(n_168), .B(n_126), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_172), .B(n_125), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_154), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_181), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_170), .B(n_120), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_159), .A2(n_114), .B1(n_128), .B2(n_127), .Y(n_216) );
INVx6_ASAP7_75t_L g217 ( .A(n_177), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_178), .A2(n_131), .B1(n_128), .B2(n_97), .Y(n_218) );
INVx8_ASAP7_75t_L g219 ( .A(n_159), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_171), .A2(n_101), .B(n_144), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_174), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_177), .B(n_131), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_199), .B(n_171), .Y(n_223) );
O2A1O1Ixp5_ASAP7_75t_L g224 ( .A1(n_186), .A2(n_166), .B(n_154), .C(n_169), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_221), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_193), .B(n_177), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_213), .A2(n_182), .B(n_174), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_219), .A2(n_169), .B1(n_154), .B2(n_166), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_200), .B(n_179), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_219), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_201), .B(n_172), .Y(n_231) );
OAI21x1_ASAP7_75t_L g232 ( .A1(n_184), .A2(n_154), .B(n_166), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_218), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_205), .B(n_159), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_192), .B(n_175), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_213), .A2(n_182), .B(n_174), .Y(n_236) );
INVx1_ASAP7_75t_SL g237 ( .A(n_192), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_205), .B(n_166), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_194), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_209), .A2(n_182), .B(n_157), .Y(n_240) );
AOI21x1_ASAP7_75t_L g241 ( .A1(n_184), .A2(n_157), .B(n_164), .Y(n_241) );
INVx4_ASAP7_75t_L g242 ( .A(n_219), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_185), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_193), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_212), .A2(n_164), .B(n_175), .Y(n_245) );
BUFx4f_ASAP7_75t_L g246 ( .A(n_219), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_185), .B(n_177), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_194), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_221), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_198), .A2(n_181), .B(n_141), .C(n_145), .Y(n_250) );
AO22x1_ASAP7_75t_L g251 ( .A1(n_221), .A2(n_159), .B1(n_144), .B2(n_145), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_221), .B(n_142), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_217), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_221), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_235), .B(n_187), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_236), .A2(n_206), .B(n_203), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_246), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_SL g258 ( .A1(n_243), .A2(n_196), .B(n_188), .C(n_189), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_227), .A2(n_190), .B(n_220), .Y(n_259) );
NOR2xp67_ASAP7_75t_L g260 ( .A(n_242), .B(n_188), .Y(n_260) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_232), .A2(n_196), .B(n_189), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_242), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_233), .A2(n_210), .B1(n_195), .B2(n_215), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_SL g264 ( .A1(n_243), .A2(n_208), .B(n_204), .C(n_214), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_237), .B(n_211), .Y(n_265) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_232), .A2(n_208), .B(n_214), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_238), .B(n_191), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_240), .A2(n_222), .B(n_197), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_245), .A2(n_202), .B(n_204), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_238), .B(n_202), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_223), .A2(n_202), .B(n_216), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_246), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_246), .Y(n_273) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_241), .A2(n_158), .B(n_176), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_247), .B(n_217), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_239), .Y(n_276) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_274), .A2(n_224), .B(n_241), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_265), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_262), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_276), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_274), .A2(n_252), .B(n_239), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_260), .B(n_248), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_276), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_255), .B(n_248), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_267), .B(n_234), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_266), .A2(n_228), .B(n_244), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_262), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g288 ( .A1(n_259), .A2(n_250), .B(n_231), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_267), .B(n_247), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_270), .B(n_229), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_266), .A2(n_244), .B(n_253), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_258), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_263), .A2(n_233), .B1(n_242), .B2(n_230), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_264), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_270), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_275), .B(n_230), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_261), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_260), .B(n_244), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_273), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_283), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_279), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_283), .B(n_261), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_279), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_280), .Y(n_304) );
INVx3_ASAP7_75t_SL g305 ( .A(n_299), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_280), .B(n_275), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_287), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_280), .Y(n_308) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_288), .A2(n_271), .B(n_269), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_297), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_292), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_295), .B(n_273), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_296), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_297), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_292), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_284), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_284), .B(n_273), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_291), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_277), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_299), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_294), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_277), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_285), .B(n_144), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_294), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_285), .B(n_257), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_277), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_289), .B(n_257), .Y(n_329) );
OA21x2_ASAP7_75t_L g330 ( .A1(n_286), .A2(n_256), .B(n_268), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_286), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_277), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_310), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_302), .B(n_298), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_310), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_304), .B(n_289), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_302), .B(n_288), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_304), .B(n_298), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_317), .B(n_290), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_308), .B(n_290), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_313), .B(n_278), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_310), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_329), .A2(n_293), .B1(n_296), .B2(n_282), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_308), .B(n_145), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_314), .B(n_281), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_308), .B(n_281), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_314), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_313), .B(n_293), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_314), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_324), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_300), .Y(n_351) );
AOI22xp33_ASAP7_75t_SL g352 ( .A1(n_307), .A2(n_272), .B1(n_225), .B2(n_249), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_305), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_316), .B(n_5), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_316), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_311), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_317), .B(n_5), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_307), .B(n_6), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_301), .B(n_6), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_321), .B(n_142), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_306), .B(n_225), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_306), .B(n_225), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_324), .Y(n_363) );
OAI22xp5_ASAP7_75t_SL g364 ( .A1(n_305), .A2(n_207), .B1(n_8), .B2(n_9), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_318), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_301), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_319), .B(n_7), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_319), .B(n_225), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_324), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_301), .B(n_7), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_328), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_303), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_328), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_321), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_318), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_311), .B(n_225), .Y(n_376) );
INVx2_ASAP7_75t_R g377 ( .A(n_331), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_315), .B(n_8), .Y(n_378) );
INVx2_ASAP7_75t_SL g379 ( .A(n_322), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_315), .B(n_9), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_329), .A2(n_254), .B1(n_249), .B2(n_253), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_323), .B(n_249), .Y(n_382) );
OR2x6_ASAP7_75t_L g383 ( .A(n_309), .B(n_251), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_323), .Y(n_384) );
NOR2x1_ASAP7_75t_SL g385 ( .A(n_322), .B(n_249), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_326), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_318), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_337), .B(n_332), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_350), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_351), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_337), .B(n_332), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_351), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_356), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_356), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_336), .B(n_325), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_353), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_384), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_353), .B(n_305), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_355), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_337), .B(n_328), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_334), .B(n_332), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_334), .B(n_331), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_336), .B(n_325), .Y(n_403) );
INVx4_ASAP7_75t_L g404 ( .A(n_353), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_350), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_372), .B(n_326), .Y(n_406) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_358), .B(n_322), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_355), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_341), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_341), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_350), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_334), .B(n_320), .Y(n_412) );
AND2x4_ASAP7_75t_SL g413 ( .A(n_370), .B(n_312), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_384), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_334), .B(n_320), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_370), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_386), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_363), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_366), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_363), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_338), .B(n_320), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_338), .B(n_309), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_367), .B(n_312), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_342), .B(n_330), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_342), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_363), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_347), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_347), .B(n_330), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_372), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_358), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_359), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_349), .B(n_333), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_359), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_349), .B(n_330), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_369), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_366), .B(n_330), .Y(n_438) );
INVx4_ASAP7_75t_L g439 ( .A(n_379), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_333), .B(n_330), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_354), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_333), .B(n_327), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_374), .Y(n_443) );
INVx3_ASAP7_75t_R g444 ( .A(n_382), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_369), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_374), .B(n_327), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_335), .B(n_10), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_335), .B(n_11), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_335), .B(n_11), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_369), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_379), .B(n_56), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_360), .B(n_12), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_340), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_360), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_360), .B(n_13), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_371), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_371), .B(n_15), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_371), .B(n_16), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_373), .Y(n_459) );
BUFx2_ASAP7_75t_L g460 ( .A(n_373), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_373), .B(n_17), .Y(n_461) );
BUFx2_ASAP7_75t_L g462 ( .A(n_345), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_346), .B(n_17), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_346), .B(n_18), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_352), .B(n_254), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_454), .B(n_348), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_390), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_390), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_392), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_443), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_404), .B(n_439), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_460), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_420), .Y(n_473) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_404), .B(n_357), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_402), .B(n_345), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_409), .B(n_368), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_392), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_424), .A2(n_364), .B1(n_343), .B2(n_383), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_410), .B(n_368), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_417), .B(n_413), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_413), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_460), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_420), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_393), .Y(n_484) );
NAND2x1p5_ASAP7_75t_L g485 ( .A(n_451), .B(n_357), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_404), .B(n_352), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_402), .B(n_345), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_432), .B(n_340), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_393), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_389), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_394), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_389), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_452), .A2(n_364), .B1(n_343), .B2(n_455), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_453), .B(n_378), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_405), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_405), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_402), .B(n_345), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_394), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_439), .B(n_385), .Y(n_499) );
INVx2_ASAP7_75t_SL g500 ( .A(n_396), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_397), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_439), .B(n_385), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_442), .B(n_339), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_397), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_396), .B(n_378), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_418), .Y(n_506) );
OR2x6_ASAP7_75t_L g507 ( .A(n_465), .B(n_383), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_446), .B(n_361), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_421), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_446), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_418), .B(n_339), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_411), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_400), .B(n_380), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_388), .B(n_361), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_399), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_408), .Y(n_516) );
AOI21xp33_ASAP7_75t_L g517 ( .A1(n_452), .A2(n_380), .B(n_381), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_400), .B(n_377), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_427), .B(n_429), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_427), .B(n_365), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_414), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_388), .B(n_362), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_401), .B(n_377), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_401), .B(n_377), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_442), .B(n_382), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_424), .B(n_382), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_415), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_407), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_424), .B(n_382), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_429), .B(n_365), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_391), .B(n_362), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_451), .B(n_381), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_434), .B(n_387), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_391), .B(n_375), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_431), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_463), .B(n_387), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_395), .B(n_375), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_403), .B(n_375), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_434), .B(n_426), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_406), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_421), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_426), .B(n_387), .Y(n_542) );
NAND3xp33_ASAP7_75t_L g543 ( .A(n_455), .B(n_344), .C(n_376), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_419), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_412), .B(n_387), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_406), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_433), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_430), .B(n_375), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_441), .A2(n_383), .B1(n_376), .B2(n_344), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_463), .B(n_365), .Y(n_550) );
NAND2x1p5_ASAP7_75t_L g551 ( .A(n_451), .B(n_249), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_435), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_464), .B(n_365), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_398), .Y(n_554) );
INVxp33_ASAP7_75t_L g555 ( .A(n_474), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_480), .B(n_412), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_510), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_519), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_547), .B(n_430), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_519), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_540), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_473), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_546), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_515), .Y(n_564) );
NOR2x2_ASAP7_75t_L g565 ( .A(n_507), .B(n_444), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_516), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_473), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_466), .B(n_416), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_539), .B(n_462), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_521), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_527), .Y(n_571) );
AOI21xp33_ASAP7_75t_SL g572 ( .A1(n_471), .A2(n_486), .B(n_481), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_534), .Y(n_573) );
INVxp33_ASAP7_75t_L g574 ( .A(n_474), .Y(n_574) );
CKINVDCx16_ASAP7_75t_R g575 ( .A(n_513), .Y(n_575) );
AND2x2_ASAP7_75t_SL g576 ( .A(n_499), .B(n_462), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_535), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_526), .B(n_416), .Y(n_578) );
AOI32xp33_ASAP7_75t_L g579 ( .A1(n_478), .A2(n_461), .A3(n_457), .B1(n_458), .B2(n_448), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_467), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_468), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_483), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_469), .Y(n_583) );
NAND3xp33_ASAP7_75t_L g584 ( .A(n_493), .B(n_461), .C(n_457), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_477), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_493), .A2(n_425), .B1(n_423), .B2(n_458), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_552), .B(n_436), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_484), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_472), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_500), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_470), .B(n_444), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_482), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_489), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_539), .B(n_436), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_509), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_554), .B(n_423), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_511), .B(n_491), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_529), .B(n_423), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_517), .A2(n_448), .B1(n_449), .B2(n_447), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_498), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_541), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_494), .B(n_440), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_514), .B(n_438), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_501), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_488), .B(n_18), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_511), .B(n_440), .Y(n_606) );
NOR3xp33_ASAP7_75t_L g607 ( .A(n_528), .B(n_449), .C(n_459), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_499), .Y(n_608) );
AND2x4_ASAP7_75t_L g609 ( .A(n_502), .B(n_459), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_522), .B(n_456), .Y(n_610) );
BUFx2_ASAP7_75t_L g611 ( .A(n_502), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_525), .B(n_456), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_523), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_504), .Y(n_614) );
INVx3_ASAP7_75t_L g615 ( .A(n_475), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_475), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_503), .B(n_19), .Y(n_617) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_542), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_506), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_531), .B(n_450), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_476), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_508), .B(n_450), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_536), .B(n_445), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_537), .B(n_445), .Y(n_624) );
AOI222xp33_ASAP7_75t_L g625 ( .A1(n_543), .A2(n_428), .B1(n_422), .B2(n_437), .C1(n_19), .C2(n_251), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_609), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_558), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_590), .Y(n_628) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_584), .A2(n_507), .B1(n_485), .B2(n_532), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_560), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_609), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_590), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_575), .B(n_487), .Y(n_633) );
NAND2x1_ASAP7_75t_L g634 ( .A(n_611), .B(n_507), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_557), .B(n_548), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_555), .A2(n_479), .B(n_505), .Y(n_636) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_572), .A2(n_517), .B(n_551), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_584), .A2(n_497), .B1(n_487), .B2(n_549), .Y(n_638) );
OAI21xp5_ASAP7_75t_L g639 ( .A1(n_625), .A2(n_549), .B(n_550), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_595), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_567), .Y(n_641) );
OA21x2_ASAP7_75t_L g642 ( .A1(n_597), .A2(n_548), .B(n_520), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_618), .B(n_538), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_586), .A2(n_545), .B1(n_497), .B2(n_518), .Y(n_644) );
NOR2xp67_ASAP7_75t_L g645 ( .A(n_608), .B(n_533), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_625), .A2(n_553), .B1(n_545), .B2(n_524), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_616), .B(n_533), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_596), .A2(n_520), .B1(n_530), .B2(n_544), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_615), .B(n_490), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_562), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_561), .B(n_496), .Y(n_651) );
OAI31xp33_ASAP7_75t_L g652 ( .A1(n_574), .A2(n_512), .A3(n_495), .B(n_492), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_559), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_559), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_587), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_576), .A2(n_383), .B1(n_428), .B2(n_422), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_617), .B(n_253), .C(n_173), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_587), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_607), .A2(n_383), .B1(n_254), .B2(n_226), .Y(n_659) );
INVxp67_ASAP7_75t_L g660 ( .A(n_582), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_621), .A2(n_383), .B1(n_254), .B2(n_173), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_605), .A2(n_160), .B1(n_254), .B2(n_23), .C(n_25), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_597), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_603), .B(n_160), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_615), .B(n_21), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_567), .B(n_22), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_663), .B(n_563), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_633), .B(n_556), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_627), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_639), .A2(n_591), .B1(n_599), .B2(n_601), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_646), .A2(n_569), .B1(n_613), .B2(n_594), .Y(n_671) );
AOI21xp33_ASAP7_75t_SL g672 ( .A1(n_629), .A2(n_579), .B(n_565), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_637), .A2(n_613), .B1(n_577), .B2(n_606), .C(n_570), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g674 ( .A1(n_637), .A2(n_594), .B(n_602), .C(n_606), .Y(n_674) );
NOR4xp25_ASAP7_75t_L g675 ( .A(n_632), .B(n_564), .C(n_566), .D(n_571), .Y(n_675) );
AOI211xp5_ASAP7_75t_SL g676 ( .A1(n_638), .A2(n_593), .B(n_580), .C(n_588), .Y(n_676) );
NAND4xp25_ASAP7_75t_SL g677 ( .A(n_644), .B(n_598), .C(n_568), .D(n_612), .Y(n_677) );
AND4x1_ASAP7_75t_L g678 ( .A(n_639), .B(n_578), .C(n_623), .D(n_600), .Y(n_678) );
AOI222xp33_ASAP7_75t_L g679 ( .A1(n_632), .A2(n_628), .B1(n_641), .B2(n_655), .C1(n_654), .C2(n_658), .Y(n_679) );
AOI322xp5_ASAP7_75t_L g680 ( .A1(n_634), .A2(n_573), .A3(n_604), .B1(n_583), .B2(n_619), .C1(n_614), .C2(n_585), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_653), .B(n_581), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_657), .A2(n_592), .B1(n_589), .B2(n_610), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_645), .A2(n_622), .B1(n_620), .B2(n_624), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_640), .A2(n_217), .B1(n_29), .B2(n_31), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_636), .A2(n_26), .B1(n_33), .B2(n_34), .C(n_36), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g686 ( .A1(n_652), .A2(n_38), .B(n_39), .Y(n_686) );
INVx1_ASAP7_75t_SL g687 ( .A(n_641), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_652), .A2(n_217), .B1(n_43), .B2(n_44), .C(n_45), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_630), .A2(n_41), .B1(n_49), .B2(n_50), .C(n_51), .Y(n_689) );
OAI21xp33_ASAP7_75t_L g690 ( .A1(n_648), .A2(n_54), .B(n_55), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_SL g691 ( .A1(n_665), .A2(n_57), .B(n_58), .C(n_59), .Y(n_691) );
OAI322xp33_ASAP7_75t_SL g692 ( .A1(n_635), .A2(n_61), .A3(n_62), .B1(n_64), .B2(n_66), .C1(n_67), .C2(n_74), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_651), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_664), .B(n_77), .C(n_79), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_660), .A2(n_81), .B1(n_84), .B2(n_86), .C(n_88), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g696 ( .A1(n_659), .A2(n_89), .B(n_92), .C(n_656), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_666), .A2(n_642), .B(n_631), .Y(n_697) );
AOI211xp5_ASAP7_75t_L g698 ( .A1(n_662), .A2(n_626), .B(n_647), .C(n_643), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_642), .B(n_650), .Y(n_699) );
NAND4xp25_ASAP7_75t_L g700 ( .A(n_661), .B(n_493), .C(n_478), .D(n_637), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_700), .B(n_672), .C(n_673), .Y(n_701) );
NOR2x1_ASAP7_75t_L g702 ( .A(n_674), .B(n_677), .Y(n_702) );
NAND4xp25_ASAP7_75t_L g703 ( .A(n_670), .B(n_676), .C(n_679), .D(n_686), .Y(n_703) );
AOI321xp33_ASAP7_75t_L g704 ( .A1(n_671), .A2(n_675), .A3(n_698), .B1(n_697), .B2(n_682), .C(n_688), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_687), .A2(n_693), .B1(n_699), .B2(n_692), .C(n_669), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_683), .A2(n_682), .B1(n_678), .B2(n_668), .Y(n_706) );
NOR3xp33_ASAP7_75t_L g707 ( .A(n_701), .B(n_685), .C(n_696), .Y(n_707) );
XNOR2xp5_ASAP7_75t_L g708 ( .A(n_703), .B(n_684), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g709 ( .A(n_704), .B(n_684), .C(n_690), .D(n_680), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_702), .B(n_667), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_710), .Y(n_711) );
INVx3_ASAP7_75t_L g712 ( .A(n_708), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_709), .B(n_706), .Y(n_713) );
NOR2x1_ASAP7_75t_L g714 ( .A(n_712), .B(n_707), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_711), .Y(n_715) );
OAI22xp33_ASAP7_75t_SL g716 ( .A1(n_715), .A2(n_713), .B1(n_712), .B2(n_681), .Y(n_716) );
AND2x4_ASAP7_75t_L g717 ( .A(n_714), .B(n_649), .Y(n_717) );
BUFx2_ASAP7_75t_L g718 ( .A(n_717), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_716), .B(n_705), .Y(n_719) );
OA21x2_ASAP7_75t_L g720 ( .A1(n_719), .A2(n_695), .B(n_689), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_720), .Y(n_721) );
AOI21xp33_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_691), .B(n_694), .Y(n_722) );
endmodule