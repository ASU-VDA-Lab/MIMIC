module fake_jpeg_12406_n_424 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_424);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_424;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_6),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_46),
.B(n_51),
.Y(n_104)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_52),
.B(n_86),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_53),
.Y(n_142)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_54),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx5_ASAP7_75t_SL g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_60),
.Y(n_111)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g134 ( 
.A(n_65),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

NAND2x1_ASAP7_75t_L g74 ( 
.A(n_24),
.B(n_0),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_74),
.B(n_23),
.C(n_30),
.Y(n_138)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_16),
.B(n_8),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_83),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_18),
.B(n_45),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_39),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_32),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_20),
.B(n_40),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_39),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_90),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_89),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_18),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_95),
.A2(n_4),
.B(n_6),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_32),
.B1(n_44),
.B2(n_17),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_99),
.A2(n_114),
.B1(n_120),
.B2(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_41),
.B1(n_44),
.B2(n_21),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_100),
.A2(n_124),
.B1(n_129),
.B2(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_61),
.B(n_33),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_113),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_50),
.B(n_34),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_79),
.A2(n_44),
.B1(n_17),
.B2(n_38),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_44),
.B1(n_38),
.B2(n_37),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_87),
.A2(n_21),
.B1(n_34),
.B2(n_36),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_21),
.B1(n_36),
.B2(n_37),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_35),
.B1(n_43),
.B2(n_45),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_126),
.A2(n_133),
.B1(n_65),
.B2(n_60),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_64),
.A2(n_36),
.B1(n_43),
.B2(n_25),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_60),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_69),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_66),
.A2(n_35),
.B1(n_25),
.B2(n_36),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_72),
.A2(n_36),
.B1(n_23),
.B2(n_10),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_74),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_67),
.A2(n_23),
.B1(n_30),
.B2(n_3),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_141),
.A2(n_49),
.B1(n_57),
.B2(n_53),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_143),
.B(n_151),
.Y(n_204)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_106),
.B(n_54),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_146),
.B(n_184),
.Y(n_213)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_147),
.Y(n_212)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_148),
.Y(n_216)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_134),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_153),
.B(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_154),
.Y(n_229)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

OAI22x1_ASAP7_75t_L g205 ( 
.A1(n_157),
.A2(n_169),
.B1(n_180),
.B2(n_185),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_113),
.A2(n_55),
.B1(n_58),
.B2(n_63),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_158),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_134),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_168),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_91),
.Y(n_162)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_163),
.Y(n_202)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g166 ( 
.A1(n_114),
.A2(n_48),
.B1(n_73),
.B2(n_56),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_166),
.A2(n_171),
.B1(n_145),
.B2(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_117),
.A2(n_69),
.B1(n_59),
.B2(n_65),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_9),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_174),
.B(n_183),
.Y(n_220)
);

OR2x2_ASAP7_75t_SL g175 ( 
.A(n_97),
.B(n_15),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_187),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_92),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_177),
.Y(n_201)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_182),
.Y(n_225)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_117),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_180)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_181),
.Y(n_207)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_116),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_92),
.B(n_10),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_142),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_120),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_186),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_122),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_10),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_136),
.Y(n_222)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_93),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_152),
.A2(n_99),
.B1(n_133),
.B2(n_103),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_193),
.A2(n_227),
.B1(n_231),
.B2(n_156),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_125),
.B(n_122),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_203),
.A2(n_202),
.B(n_205),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_94),
.C(n_127),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_211),
.C(n_221),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_209),
.A2(n_215),
.B1(n_233),
.B2(n_232),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_150),
.B(n_107),
.Y(n_211)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_187),
.B(n_107),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_214),
.B(n_227),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_171),
.A2(n_123),
.B1(n_93),
.B2(n_94),
.Y(n_215)
);

NOR2x1p5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_135),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_217),
.B(n_194),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_164),
.B(n_144),
.C(n_147),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_183),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_152),
.A2(n_123),
.B1(n_127),
.B2(n_121),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_166),
.A2(n_121),
.B1(n_136),
.B2(n_81),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_172),
.A2(n_4),
.B1(n_12),
.B2(n_13),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_149),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_250),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_235),
.A2(n_246),
.B1(n_247),
.B2(n_268),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_237),
.B(n_242),
.Y(n_295)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_214),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_239),
.B(n_245),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_178),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_240),
.A2(n_266),
.B(n_207),
.Y(n_287)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_175),
.C(n_15),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_251),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_196),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_221),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_243),
.B(n_249),
.Y(n_298)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_244),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_177),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_193),
.A2(n_191),
.B1(n_162),
.B2(n_161),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_208),
.A2(n_188),
.B1(n_160),
.B2(n_148),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_248),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_226),
.B(n_182),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_181),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_253),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_170),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_256),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

BUFx24_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_170),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_223),
.Y(n_257)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_258),
.A2(n_262),
.B1(n_229),
.B2(n_213),
.Y(n_283)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_200),
.Y(n_260)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

INVx8_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_209),
.A2(n_232),
.B1(n_215),
.B2(n_203),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_198),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_264),
.Y(n_296)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_200),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_220),
.B(n_222),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_226),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_267),
.A2(n_270),
.B(n_217),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_231),
.A2(n_205),
.B1(n_229),
.B2(n_195),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_219),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_270),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_273),
.B(n_278),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_276),
.A2(n_264),
.B(n_260),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_240),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_245),
.A2(n_239),
.B(n_267),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_279),
.A2(n_282),
.B(n_287),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_267),
.A2(n_195),
.B(n_194),
.Y(n_282)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_240),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_288),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_262),
.A2(n_266),
.B1(n_236),
.B2(n_235),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_292),
.B1(n_300),
.B2(n_240),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_268),
.A2(n_199),
.B1(n_228),
.B2(n_230),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_234),
.B(n_192),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_250),
.C(n_254),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_246),
.A2(n_199),
.B1(n_230),
.B2(n_212),
.Y(n_300)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_236),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_307),
.C(n_310),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_265),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_319),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_309),
.A2(n_321),
.B1(n_317),
.B2(n_312),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_299),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_293),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_313),
.C(n_314),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_256),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_252),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_296),
.Y(n_315)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_315),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_290),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_318),
.Y(n_338)
);

FAx1_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_272),
.CI(n_274),
.CON(n_348),
.SN(n_348)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_257),
.C(n_248),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_295),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_294),
.A2(n_261),
.B1(n_238),
.B2(n_244),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_322),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_271),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_323),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_281),
.B(n_269),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_328),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_271),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_325),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_216),
.Y(n_326)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_326),
.Y(n_350)
);

OAI21x1_ASAP7_75t_L g327 ( 
.A1(n_282),
.A2(n_210),
.B(n_255),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_276),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_287),
.B(n_219),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_271),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_329),
.Y(n_349)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_330),
.Y(n_358)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_320),
.Y(n_333)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_333),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_334),
.A2(n_348),
.B(n_307),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_306),
.A2(n_292),
.B1(n_300),
.B2(n_283),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_345),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_301),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_337),
.Y(n_357)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_346),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_344),
.A2(n_284),
.B1(n_313),
.B2(n_210),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_306),
.A2(n_291),
.B1(n_272),
.B2(n_289),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_291),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_312),
.A2(n_280),
.B(n_297),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_351),
.A2(n_303),
.B(n_328),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_316),
.A2(n_297),
.B1(n_284),
.B2(n_216),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_309),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_304),
.C(n_310),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_360),
.C(n_366),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_342),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_355),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_311),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_359),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_324),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_347),
.C(n_337),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_362),
.A2(n_365),
.B(n_368),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_363),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_343),
.B(n_347),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_364),
.B(n_365),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_343),
.B(n_314),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_341),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_367),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_368),
.A2(n_352),
.B(n_346),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_212),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_339),
.C(n_344),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_336),
.B(n_349),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_350),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_376),
.B(n_378),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_361),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_383),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_357),
.B(n_345),
.Y(n_381)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_381),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g382 ( 
.A(n_362),
.B(n_348),
.CI(n_351),
.CON(n_382),
.SN(n_382)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_385),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_340),
.C(n_335),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_384),
.B(n_386),
.Y(n_393)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_384),
.B(n_360),
.C(n_359),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_392),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_380),
.B(n_358),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_389),
.B(n_397),
.Y(n_406)
);

XNOR2x1_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_366),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_398),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_375),
.B(n_356),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_386),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_381),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_333),
.Y(n_397)
);

XNOR2x1_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_364),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_377),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_400),
.B(n_401),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_375),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_395),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_402),
.B(n_407),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_376),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_403),
.B(n_404),
.Y(n_412)
);

MAJx2_ASAP7_75t_L g404 ( 
.A(n_388),
.B(n_379),
.C(n_378),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_399),
.B(n_394),
.C(n_391),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_413),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_406),
.B(n_390),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_411),
.A2(n_379),
.B1(n_385),
.B2(n_372),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_405),
.B(n_373),
.Y(n_413)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_414),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_412),
.B(n_405),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_415),
.A2(n_416),
.B(n_408),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_413),
.B(n_404),
.C(n_398),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_418),
.B(n_417),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_420),
.A2(n_419),
.B1(n_411),
.B2(n_410),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_421),
.Y(n_422)
);

A2O1A1Ixp33_ASAP7_75t_L g423 ( 
.A1(n_422),
.A2(n_416),
.B(n_382),
.C(n_348),
.Y(n_423)
);

OAI321xp33_ASAP7_75t_L g424 ( 
.A1(n_423),
.A2(n_353),
.A3(n_363),
.B1(n_370),
.B2(n_382),
.C(n_407),
.Y(n_424)
);


endmodule