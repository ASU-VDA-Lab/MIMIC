module fake_jpeg_19377_n_319 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_23),
.A2(n_0),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_0),
.Y(n_73)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_30),
.Y(n_62)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_19),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_54),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_63),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_61),
.B(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_18),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_17),
.B1(n_36),
.B2(n_33),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_44),
.B1(n_40),
.B2(n_22),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_30),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_33),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_66),
.Y(n_115)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_20),
.C(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_43),
.B(n_27),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_40),
.A2(n_17),
.B1(n_35),
.B2(n_27),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_48),
.B1(n_46),
.B2(n_41),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_82),
.B(n_42),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_40),
.B1(n_45),
.B2(n_44),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_84),
.A2(n_86),
.B1(n_88),
.B2(n_96),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_35),
.B1(n_25),
.B2(n_32),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_76),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_32),
.B1(n_25),
.B2(n_20),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_90),
.A2(n_38),
.B(n_21),
.Y(n_129)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_40),
.B1(n_48),
.B2(n_46),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_48),
.B1(n_46),
.B2(n_39),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_98),
.A2(n_101),
.B1(n_107),
.B2(n_117),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_29),
.B1(n_28),
.B2(n_26),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_102),
.B1(n_104),
.B2(n_108),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_51),
.A2(n_29),
.B1(n_26),
.B2(n_24),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_48),
.B1(n_46),
.B2(n_39),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_57),
.A2(n_41),
.B1(n_42),
.B2(n_24),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_67),
.A2(n_68),
.B1(n_74),
.B2(n_61),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_29),
.B1(n_26),
.B2(n_31),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_114),
.B1(n_116),
.B2(n_53),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_74),
.A2(n_60),
.B1(n_75),
.B2(n_76),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_74),
.A2(n_41),
.B1(n_42),
.B2(n_31),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_21),
.B1(n_31),
.B2(n_26),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_56),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_125),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_81),
.B1(n_83),
.B2(n_85),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_127),
.B1(n_139),
.B2(n_151),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_75),
.B1(n_76),
.B2(n_72),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_126),
.B(n_129),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_56),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_60),
.B(n_53),
.C(n_41),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_31),
.B1(n_21),
.B2(n_56),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_38),
.B(n_12),
.C(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_135),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_38),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_150),
.C(n_153),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_69),
.Y(n_135)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_148),
.Y(n_156)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_42),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_116),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_11),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_144),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_80),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_142),
.B(n_147),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_11),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_90),
.B(n_10),
.C(n_16),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_3),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_97),
.B(n_12),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_93),
.A2(n_69),
.B(n_1),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_108),
.A2(n_69),
.B1(n_0),
.B2(n_4),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_3),
.C(n_4),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_158),
.A2(n_164),
.B(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_163),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_149),
.A2(n_87),
.B1(n_92),
.B2(n_91),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_182),
.B1(n_148),
.B2(n_133),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_87),
.B(n_80),
.C(n_107),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_167),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_123),
.A2(n_111),
.B1(n_113),
.B2(n_97),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_186),
.B1(n_140),
.B2(n_139),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_82),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_112),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_173),
.B(n_176),
.Y(n_204)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_113),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_122),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_138),
.B(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_149),
.A2(n_140),
.B1(n_123),
.B2(n_126),
.Y(n_182)
);

BUFx24_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

INVx5_ASAP7_75t_SL g195 ( 
.A(n_184),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_130),
.B(n_94),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_185),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_128),
.A2(n_100),
.B1(n_110),
.B2(n_89),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_135),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_208),
.Y(n_227)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_140),
.B(n_129),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g229 ( 
.A1(n_190),
.A2(n_194),
.B1(n_196),
.B2(n_205),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_182),
.B1(n_158),
.B2(n_161),
.Y(n_216)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_151),
.B1(n_150),
.B2(n_143),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_162),
.A2(n_148),
.B(n_132),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_199),
.A2(n_205),
.B(n_206),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_130),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_203),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_153),
.Y(n_203)
);

AND2x4_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_119),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_94),
.C(n_7),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_154),
.C(n_175),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_6),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_94),
.B(n_7),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_211),
.B(n_12),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_162),
.A2(n_6),
.B(n_7),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_8),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_214),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_157),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_189),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_220),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_158),
.B1(n_164),
.B2(n_155),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_223),
.Y(n_251)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_155),
.B1(n_169),
.B2(n_179),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_224),
.A2(n_238),
.B(n_197),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_225),
.A2(n_229),
.B1(n_205),
.B2(n_207),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_174),
.C(n_165),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_234),
.C(n_236),
.Y(n_244)
);

MAJx2_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_183),
.C(n_178),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_230),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_186),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_204),
.A2(n_211),
.B(n_191),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_159),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_209),
.B(n_176),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_171),
.C(n_160),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_202),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_214),
.C(n_213),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_198),
.B1(n_205),
.B2(n_194),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_187),
.B(n_171),
.C(n_183),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_206),
.C(n_190),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_240),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_235),
.B1(n_224),
.B2(n_231),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_191),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_253),
.C(n_258),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_252),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_232),
.B(n_208),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_226),
.C(n_230),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_218),
.C(n_229),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_256),
.A2(n_231),
.B1(n_216),
.B2(n_221),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_197),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_234),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_227),
.B(n_239),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_260),
.A2(n_261),
.B1(n_265),
.B2(n_248),
.Y(n_283)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_242),
.A2(n_229),
.B1(n_228),
.B2(n_194),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_212),
.Y(n_266)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_244),
.B(n_241),
.Y(n_285)
);

INVx11_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_275),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_244),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_212),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_229),
.C(n_190),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_252),
.C(n_250),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_194),
.B1(n_202),
.B2(n_210),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_257),
.B1(n_256),
.B2(n_249),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_210),
.Y(n_275)
);

INVxp33_ASAP7_75t_SL g276 ( 
.A(n_268),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_276),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_281),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_265),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_284),
.B1(n_267),
.B2(n_272),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_246),
.B1(n_258),
.B2(n_250),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_269),
.C(n_262),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_184),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_292),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_288),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_296),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_274),
.Y(n_295)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_259),
.C(n_273),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_297),
.A2(n_285),
.B(n_279),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_303),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_304),
.B(n_305),
.Y(n_306)
);

OAI321xp33_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_266),
.A3(n_270),
.B1(n_276),
.B2(n_275),
.C(n_274),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_259),
.B(n_286),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_263),
.Y(n_305)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_287),
.Y(n_307)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_184),
.B(n_195),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_305),
.B(n_294),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_294),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_302),
.A2(n_296),
.B1(n_278),
.B2(n_264),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_301),
.C(n_184),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_312),
.Y(n_314)
);

OAI21x1_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_306),
.B(n_307),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_306),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_308),
.A3(n_314),
.B1(n_195),
.B2(n_168),
.C1(n_16),
.C2(n_15),
.Y(n_317)
);

OAI321xp33_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_168),
.C(n_240),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_14),
.Y(n_319)
);


endmodule