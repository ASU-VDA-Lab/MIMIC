module fake_jpeg_14685_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_27),
.C(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_19),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_32),
.C(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_54),
.Y(n_63)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_16),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_19),
.B1(n_30),
.B2(n_16),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_19),
.B1(n_23),
.B2(n_30),
.Y(n_65)
);

NAND2x1_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_20),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_38),
.Y(n_76)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_67),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_68),
.Y(n_84)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_23),
.B(n_21),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_74),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_32),
.C(n_37),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_73),
.Y(n_86)
);

AO22x1_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_44),
.B1(n_32),
.B2(n_20),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_34),
.B1(n_48),
.B2(n_50),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_37),
.C(n_34),
.Y(n_77)
);

AOI22x1_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_39),
.B1(n_20),
.B2(n_37),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_58),
.B1(n_55),
.B2(n_34),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_51),
.B(n_29),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_96),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_91),
.B(n_99),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_68),
.B(n_21),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_90),
.Y(n_118)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_94),
.Y(n_107)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_87),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_47),
.B1(n_18),
.B2(n_26),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_72),
.B(n_28),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_47),
.B1(n_53),
.B2(n_42),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_66),
.B1(n_78),
.B2(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_42),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_63),
.B(n_27),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_37),
.C(n_17),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_28),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_84),
.B(n_96),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_103),
.A2(n_89),
.B(n_90),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_108),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_84),
.B1(n_86),
.B2(n_99),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_111),
.B1(n_80),
.B2(n_89),
.Y(n_126)
);

BUFx24_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_78),
.B1(n_64),
.B2(n_60),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_95),
.B1(n_87),
.B2(n_81),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_64),
.B1(n_53),
.B2(n_75),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_97),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_28),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_120),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_126),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_82),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_118),
.B(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_134),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_26),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_138),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_26),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_113),
.B(n_107),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_17),
.C(n_18),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_139),
.C(n_110),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_17),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_52),
.C(n_22),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_145),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_116),
.B(n_117),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_147),
.B1(n_151),
.B2(n_153),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_116),
.B(n_117),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_125),
.A2(n_111),
.B1(n_119),
.B2(n_108),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_154),
.B1(n_127),
.B2(n_133),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_105),
.B(n_102),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_104),
.B(n_121),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_102),
.C(n_109),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_124),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_158),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_151),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_162),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_152),
.A2(n_135),
.B1(n_129),
.B2(n_123),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_137),
.B1(n_139),
.B2(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_124),
.B1(n_138),
.B2(n_136),
.Y(n_163)
);

BUFx12_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_148),
.Y(n_174)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_166),
.Y(n_173)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_156),
.C(n_163),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_146),
.A2(n_114),
.B1(n_109),
.B2(n_52),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_140),
.Y(n_175)
);

OAI211xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_147),
.B(n_142),
.C(n_141),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_164),
.A3(n_109),
.B1(n_14),
.B2(n_13),
.C1(n_12),
.C2(n_7),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_149),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_176),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_1),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_1),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_154),
.B(n_145),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_168),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_158),
.B1(n_164),
.B2(n_161),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_190)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_14),
.B1(n_12),
.B2(n_4),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_22),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_175),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_2),
.Y(n_187)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_184),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_196)
);

AOI321xp33_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_173),
.A3(n_169),
.B1(n_172),
.B2(n_22),
.C(n_8),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_5),
.B(n_6),
.Y(n_195)
);

OAI321xp33_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_186),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_2),
.Y(n_194)
);

OAI21x1_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_196),
.B(n_191),
.Y(n_198)
);

OAI21x1_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_9),
.B(n_11),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_198),
.B(n_200),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_197),
.A2(n_188),
.B(n_11),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_193),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_9),
.B(n_22),
.C(n_201),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_22),
.Y(n_204)
);


endmodule