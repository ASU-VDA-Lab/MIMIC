module fake_jpeg_22031_n_228 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_0),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_38),
.B(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_2),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_5),
.Y(n_76)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_23),
.A2(n_2),
.B(n_3),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_3),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_5),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_29),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_19),
.B1(n_23),
.B2(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_49),
.B(n_82),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_72),
.B1(n_8),
.B2(n_9),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_19),
.B1(n_27),
.B2(n_32),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_54),
.B1(n_62),
.B2(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_46),
.B1(n_20),
.B2(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_28),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_60),
.Y(n_96)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_35),
.B1(n_18),
.B2(n_33),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_22),
.B1(n_20),
.B2(n_35),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_69),
.B1(n_53),
.B2(n_77),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_22),
.B1(n_28),
.B2(n_31),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_24),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_15),
.Y(n_106)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_78),
.Y(n_102)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_7),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_36),
.A2(n_25),
.B1(n_34),
.B2(n_21),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_97)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_104),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_34),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_95),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_21),
.B1(n_8),
.B2(n_7),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_98),
.B1(n_105),
.B2(n_103),
.Y(n_126)
);

OR2x2_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_8),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_90),
.B(n_106),
.Y(n_128)
);

OAI22x1_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_69),
.B1(n_61),
.B2(n_59),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_11),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_97),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_14),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_105),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_15),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_78),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_60),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_70),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_64),
.B(n_61),
.C(n_73),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_86),
.B(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_80),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_121),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_130),
.Y(n_139)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_51),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_129),
.Y(n_158)
);

INVx5_ASAP7_75t_SL g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_124),
.B(n_128),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_95),
.B1(n_99),
.B2(n_87),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_101),
.B1(n_106),
.B2(n_85),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_127),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_88),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_90),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_85),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_149),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_127),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_94),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_150),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_94),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_156),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_145),
.B1(n_157),
.B2(n_152),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_101),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_154),
.Y(n_159)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_101),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_131),
.B(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_157),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_125),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_126),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_128),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_161),
.C(n_166),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_119),
.C(n_112),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_165),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_110),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_122),
.C(n_129),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_169),
.B(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_174),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_143),
.B(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_181),
.B(n_170),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_143),
.B(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_184),
.Y(n_192)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_155),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_185),
.B(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_188),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_142),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_187),
.B(n_189),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_168),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_174),
.B(n_159),
.C(n_164),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_185),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_193),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_167),
.B(n_154),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_184),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_138),
.Y(n_196)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_149),
.B1(n_135),
.B2(n_133),
.Y(n_199)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_183),
.Y(n_202)
);

OAI21x1_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_190),
.B(n_198),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_205),
.B(n_137),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_197),
.B(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_211),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_191),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g217 ( 
.A(n_212),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_199),
.B(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_214),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_178),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_165),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_222),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_207),
.B(n_202),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_213),
.C(n_217),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_224),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_226),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_227),
.B(n_216),
.Y(n_228)
);


endmodule