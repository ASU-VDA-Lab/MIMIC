module fake_jpeg_4029_n_270 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

BUFx12f_ASAP7_75t_SL g36 ( 
.A(n_18),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_19),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_0),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_47),
.B(n_53),
.Y(n_89)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_55),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_57),
.Y(n_94)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_17),
.B(n_29),
.C(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_59),
.B(n_60),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_21),
.B1(n_17),
.B2(n_29),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_68),
.B(n_31),
.C(n_25),
.Y(n_92)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_72),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_21),
.B1(n_26),
.B2(n_19),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_70),
.B1(n_12),
.B2(n_14),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_28),
.B1(n_33),
.B2(n_30),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_67),
.B1(n_32),
.B2(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_66),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_30),
.B1(n_33),
.B2(n_22),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_36),
.A2(n_18),
.B(n_27),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_36),
.A2(n_26),
.B1(n_22),
.B2(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_41),
.B(n_26),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_85),
.B1(n_86),
.B2(n_72),
.Y(n_106)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_77),
.B(n_92),
.Y(n_113)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_81),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_31),
.B1(n_25),
.B2(n_24),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_95),
.B1(n_48),
.B2(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_27),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_65),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_67),
.B1(n_51),
.B2(n_59),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_34),
.B(n_23),
.C(n_27),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_62),
.B(n_65),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_27),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_45),
.C(n_52),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_48),
.A2(n_31),
.B1(n_25),
.B2(n_24),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_69),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_104),
.B(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_51),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_103),
.Y(n_135)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_61),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_109),
.B1(n_112),
.B2(n_118),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_122),
.B1(n_95),
.B2(n_93),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_117),
.B1(n_120),
.B2(n_88),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_111),
.Y(n_136)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_60),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_74),
.B(n_46),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_121),
.C(n_97),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_71),
.B1(n_55),
.B2(n_56),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_79),
.B1(n_82),
.B2(n_90),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_57),
.B1(n_66),
.B2(n_23),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_50),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_50),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_58),
.B1(n_23),
.B2(n_34),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_123),
.B(n_141),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_114),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_107),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_132),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_114),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_126),
.A2(n_50),
.B(n_18),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_148),
.B1(n_122),
.B2(n_119),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_88),
.B(n_93),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_115),
.B(n_101),
.Y(n_161)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_140),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_109),
.B1(n_78),
.B2(n_34),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_85),
.B1(n_75),
.B2(n_87),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_144),
.B1(n_147),
.B2(n_101),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_78),
.C(n_18),
.Y(n_171)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_142),
.B(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_75),
.B1(n_87),
.B2(n_81),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_116),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_149),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_87),
.B1(n_90),
.B2(n_84),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_110),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_97),
.A2(n_82),
.B1(n_79),
.B2(n_31),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_151),
.B(n_156),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_106),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_164),
.C(n_171),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_157),
.B1(n_175),
.B2(n_145),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_97),
.A3(n_115),
.B1(n_118),
.B2(n_112),
.C1(n_105),
.C2(n_102),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_155),
.B(n_143),
.C(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_160),
.Y(n_194)
);

BUFx12_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_167),
.B(n_170),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_166),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_34),
.A3(n_23),
.B1(n_24),
.B2(n_18),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_150),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_78),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_131),
.B1(n_130),
.B2(n_125),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_127),
.A2(n_27),
.B(n_82),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_176),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_96),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_178),
.C(n_179),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_109),
.B1(n_10),
.B2(n_11),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_96),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_9),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_137),
.B1(n_141),
.B2(n_128),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_184),
.B1(n_191),
.B2(n_162),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_142),
.B1(n_133),
.B2(n_136),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_160),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_160),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_162),
.A2(n_149),
.B1(n_131),
.B2(n_127),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_132),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_172),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_203),
.B1(n_16),
.B2(n_8),
.Y(n_221)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

OA21x2_ASAP7_75t_SL g216 ( 
.A1(n_201),
.A2(n_178),
.B(n_163),
.Y(n_216)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_204),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_123),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_1),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_217),
.B1(n_198),
.B2(n_185),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_212),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_174),
.C(n_152),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_219),
.C(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_164),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_218),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_184),
.B(n_179),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_215),
.B(n_216),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_204),
.A2(n_167),
.B1(n_170),
.B2(n_171),
.Y(n_217)
);

AOI321xp33_ASAP7_75t_L g218 ( 
.A1(n_195),
.A2(n_170),
.A3(n_169),
.B1(n_156),
.B2(n_160),
.C(n_11),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_1),
.C(n_2),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_220),
.A2(n_180),
.B(n_188),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_2),
.C(n_3),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_223),
.A2(n_181),
.B1(n_186),
.B2(n_191),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_205),
.C(n_182),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_217),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_232),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_196),
.B1(n_203),
.B2(n_187),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_203),
.B1(n_187),
.B2(n_183),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_189),
.B(n_199),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_231),
.B1(n_223),
.B2(n_222),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_202),
.B(n_201),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_221),
.Y(n_243)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_213),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_238),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_218),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_226),
.A2(n_206),
.B1(n_220),
.B2(n_208),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_240),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_236),
.B(n_215),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_243),
.C(n_225),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_245),
.B1(n_233),
.B2(n_225),
.Y(n_251)
);

O2A1O1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_219),
.B(n_4),
.C(n_5),
.Y(n_245)
);

INVxp33_ASAP7_75t_SL g247 ( 
.A(n_241),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_250),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_239),
.A2(n_227),
.B(n_228),
.Y(n_248)
);

OAI21x1_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_238),
.B(n_234),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_245),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_233),
.C(n_12),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_256),
.B(n_258),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_255),
.C(n_6),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_2),
.C(n_4),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_4),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_13),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_257),
.A2(n_248),
.B1(n_252),
.B2(n_7),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_259),
.B(n_260),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_5),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_14),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_6),
.C(n_10),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_16),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_266),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_260),
.Y(n_268)
);

OAI31xp33_ASAP7_75t_SL g269 ( 
.A1(n_268),
.A2(n_263),
.A3(n_265),
.B(n_15),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_267),
.Y(n_270)
);


endmodule