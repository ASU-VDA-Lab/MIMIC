module fake_jpeg_29461_n_552 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_552);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_552;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVxp33_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_22),
.B(n_18),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_53),
.B(n_1),
.Y(n_166)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_55),
.Y(n_156)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_56),
.Y(n_152)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_58),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_59),
.B(n_50),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_62),
.Y(n_116)
);

NOR4xp25_ASAP7_75t_L g61 ( 
.A(n_30),
.B(n_17),
.C(n_16),
.D(n_2),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_61),
.A2(n_51),
.B(n_42),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_69),
.Y(n_165)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_80),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_82),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_85),
.Y(n_137)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_87),
.Y(n_145)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

NOR2xp67_ASAP7_75t_L g90 ( 
.A(n_40),
.B(n_16),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_90),
.B(n_0),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_95),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_32),
.B(n_0),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_96),
.B(n_97),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_25),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_32),
.B(n_50),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_98),
.B(n_104),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_38),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_107),
.B(n_133),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_108),
.B(n_41),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_53),
.B(n_39),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_110),
.B(n_117),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_39),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_120),
.B(n_126),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_124),
.B(n_43),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_51),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_42),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_128),
.B(n_146),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_102),
.B(n_27),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_68),
.B(n_33),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_135),
.B(n_143),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_55),
.A2(n_38),
.B1(n_33),
.B2(n_27),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_138),
.A2(n_155),
.B1(n_73),
.B2(n_101),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_103),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_93),
.B(n_47),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_52),
.Y(n_151)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_69),
.A2(n_43),
.B1(n_47),
.B2(n_41),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_76),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_159),
.B(n_161),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_100),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_167),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_78),
.B(n_37),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_171),
.Y(n_246)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_174),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_176),
.B(n_191),
.Y(n_241)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_113),
.Y(n_177)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_177),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_67),
.B1(n_85),
.B2(n_77),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_179),
.Y(n_236)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_183),
.Y(n_259)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_184),
.Y(n_238)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_64),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_193),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_190),
.A2(n_163),
.B1(n_157),
.B2(n_165),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_192),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_131),
.B(n_150),
.Y(n_193)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_195),
.Y(n_277)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_105),
.Y(n_196)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_196),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_118),
.B(n_56),
.C(n_92),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_220),
.C(n_229),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_147),
.A2(n_99),
.B1(n_75),
.B2(n_74),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

CKINVDCx12_ASAP7_75t_R g199 ( 
.A(n_111),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_199),
.Y(n_255)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_200),
.Y(n_252)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_201),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_148),
.A2(n_58),
.B1(n_65),
.B2(n_47),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_130),
.B1(n_163),
.B2(n_157),
.Y(n_237)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_203),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_125),
.B(n_166),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_204),
.B(n_210),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_122),
.A2(n_47),
.B1(n_41),
.B2(n_25),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_205),
.A2(n_218),
.B1(n_137),
.B2(n_144),
.Y(n_249)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_136),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_209),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_145),
.A2(n_47),
.B1(n_41),
.B2(n_25),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_225),
.B1(n_141),
.B2(n_130),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_132),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_208),
.B(n_219),
.Y(n_270)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_139),
.B(n_47),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_139),
.B(n_142),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_211),
.B(n_206),
.Y(n_275)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_212),
.Y(n_272)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_111),
.Y(n_215)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

INVx4_ASAP7_75t_SL g216 ( 
.A(n_123),
.Y(n_216)
);

NAND2xp33_ASAP7_75t_SL g278 ( 
.A(n_216),
.B(n_151),
.Y(n_278)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_142),
.A2(n_41),
.B1(n_25),
.B2(n_37),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_108),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_108),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_221),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_116),
.B(n_34),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_158),
.B(n_34),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_224),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_115),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_223),
.A2(n_141),
.B1(n_112),
.B2(n_151),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_158),
.B(n_149),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_145),
.A2(n_41),
.B1(n_37),
.B2(n_34),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_106),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_226),
.Y(n_260)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_228),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_106),
.B(n_2),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_152),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_235),
.B(n_247),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g310 ( 
.A1(n_237),
.A2(n_209),
.B1(n_201),
.B2(n_185),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_149),
.B1(n_144),
.B2(n_109),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_242),
.A2(n_261),
.B1(n_265),
.B2(n_211),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_179),
.A2(n_137),
.B(n_152),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_248),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_249),
.A2(n_202),
.B1(n_248),
.B2(n_232),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_187),
.B(n_160),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_253),
.B(n_263),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_219),
.A2(n_109),
.B1(n_165),
.B2(n_156),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_197),
.B(n_229),
.C(n_210),
.Y(n_263)
);

AND2x2_ASAP7_75t_SL g303 ( 
.A(n_264),
.B(n_203),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_191),
.A2(n_2),
.B(n_3),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_271),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_213),
.A2(n_2),
.B(n_3),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_189),
.B(n_123),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_280),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_180),
.Y(n_315)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_182),
.B(n_34),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_204),
.B(n_156),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_282),
.B(n_4),
.Y(n_323)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_254),
.Y(n_286)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_286),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_240),
.Y(n_287)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_287),
.Y(n_350)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_288),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_289),
.A2(n_318),
.B1(n_324),
.B2(n_328),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_230),
.B(n_176),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_290),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_208),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_291),
.B(n_293),
.Y(n_362)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_241),
.B(n_169),
.C(n_172),
.Y(n_293)
);

AND2x6_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_194),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_294),
.A2(n_238),
.B(n_245),
.Y(n_337)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_295),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_236),
.A2(n_174),
.B1(n_227),
.B2(n_217),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_297),
.A2(n_300),
.B1(n_313),
.B2(n_314),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_268),
.A2(n_200),
.B1(n_181),
.B2(n_192),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_298),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_266),
.B(n_175),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_299),
.B(n_302),
.Y(n_367)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_234),
.Y(n_301)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_301),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_253),
.B(n_212),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_303),
.B(n_310),
.Y(n_349)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_259),
.Y(n_305)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_305),
.Y(n_372)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_276),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_306),
.B(n_308),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_244),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_309),
.Y(n_354)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_244),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_311),
.B(n_312),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_262),
.B(n_177),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_232),
.A2(n_186),
.B1(n_223),
.B2(n_170),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_268),
.A2(n_195),
.B1(n_171),
.B2(n_183),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_323),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_244),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_316),
.Y(n_361)
);

OAI222xp33_ASAP7_75t_L g317 ( 
.A1(n_256),
.A2(n_216),
.B1(n_112),
.B2(n_196),
.C1(n_184),
.C2(n_226),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_317),
.B(n_322),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_256),
.A2(n_148),
.B1(n_173),
.B2(n_112),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_246),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_233),
.A2(n_173),
.B1(n_215),
.B2(n_34),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_233),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_275),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_263),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_282),
.B(n_247),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_326),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_267),
.B(n_4),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_271),
.B(n_5),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_327),
.B(n_330),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_237),
.A2(n_20),
.B1(n_7),
.B2(n_8),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_264),
.B(n_5),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_261),
.Y(n_343)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_264),
.C(n_242),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_331),
.B(n_336),
.C(n_370),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_296),
.A2(n_322),
.B1(n_300),
.B2(n_317),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_335),
.A2(n_348),
.B1(n_356),
.B2(n_358),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_325),
.C(n_292),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_SL g396 ( 
.A(n_337),
.B(n_357),
.C(n_309),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_292),
.A2(n_296),
.B(n_285),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_340),
.A2(n_351),
.B(n_355),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_346),
.Y(n_374)
);

OA21x2_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_249),
.B(n_260),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_345),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_323),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_292),
.A2(n_257),
.B1(n_238),
.B2(n_239),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_285),
.A2(n_307),
.B(n_312),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_289),
.A2(n_257),
.B1(n_245),
.B2(n_279),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_353),
.A2(n_309),
.B1(n_310),
.B2(n_295),
.Y(n_387)
);

AOI22x1_ASAP7_75t_SL g355 ( 
.A1(n_284),
.A2(n_252),
.B1(n_272),
.B2(n_255),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_294),
.A2(n_252),
.B1(n_272),
.B2(n_273),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_307),
.A2(n_279),
.B(n_276),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_308),
.A2(n_239),
.B1(n_273),
.B2(n_250),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_316),
.A2(n_277),
.B1(n_251),
.B2(n_250),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_359),
.A2(n_305),
.B1(n_330),
.B2(n_310),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_314),
.A2(n_277),
.B1(n_251),
.B2(n_246),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_360),
.B(n_369),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_326),
.A2(n_258),
.B(n_231),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_329),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_286),
.B(n_231),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_303),
.B(n_20),
.C(n_7),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_318),
.B(n_20),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_371),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_283),
.Y(n_373)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

INVxp33_ASAP7_75t_L g376 ( 
.A(n_368),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_408),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_324),
.Y(n_377)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_377),
.Y(n_420)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_350),
.Y(n_378)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_378),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_381),
.Y(n_437)
);

OAI22x1_ASAP7_75t_L g382 ( 
.A1(n_355),
.A2(n_284),
.B1(n_303),
.B2(n_310),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_382),
.A2(n_396),
.B(n_348),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_288),
.Y(n_383)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_301),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_384),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_385),
.A2(n_387),
.B1(n_400),
.B2(n_402),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_333),
.B(n_327),
.Y(n_388)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_388),
.Y(n_436)
);

INVx13_ASAP7_75t_L g389 ( 
.A(n_355),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_389),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_333),
.B(n_319),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_393),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_350),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_391),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_336),
.B(n_328),
.C(n_306),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_406),
.C(n_363),
.Y(n_414)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_369),
.Y(n_393)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_344),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_398),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_362),
.B(n_5),
.Y(n_397)
);

NAND3xp33_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_363),
.C(n_354),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_338),
.B(n_287),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_342),
.A2(n_287),
.B1(n_20),
.B2(n_10),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_338),
.B(n_346),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_345),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_342),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_347),
.B(n_9),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_404),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_11),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_367),
.B(n_362),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_405),
.B(n_407),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_340),
.B(n_11),
.C(n_13),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_366),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_368),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_414),
.B(n_425),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_380),
.A2(n_347),
.B(n_335),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_415),
.A2(n_382),
.B(n_403),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_417),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_394),
.A2(n_353),
.B1(n_339),
.B2(n_332),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_419),
.A2(n_423),
.B1(n_432),
.B2(n_385),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_339),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_424),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_375),
.B(n_331),
.C(n_351),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_427),
.C(n_438),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_394),
.A2(n_365),
.B1(n_343),
.B2(n_349),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_337),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_349),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_392),
.B(n_371),
.C(n_359),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_429),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_396),
.A2(n_341),
.B1(n_371),
.B2(n_358),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_431),
.A2(n_404),
.B1(n_386),
.B2(n_389),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_379),
.A2(n_345),
.B1(n_341),
.B2(n_364),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_381),
.B(n_345),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_374),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_401),
.B(n_370),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_434),
.B(n_372),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_399),
.B(n_357),
.C(n_344),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_360),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_441),
.A2(n_449),
.B(n_460),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_SL g442 ( 
.A(n_434),
.B(n_408),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_442),
.A2(n_448),
.B1(n_459),
.B2(n_418),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_380),
.C(n_393),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_444),
.B(n_464),
.C(n_437),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_446),
.B(n_461),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_374),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_447),
.B(n_465),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_423),
.B(n_390),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_415),
.A2(n_379),
.B(n_404),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_450),
.A2(n_458),
.B1(n_416),
.B2(n_431),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_451),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_398),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_453),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_411),
.B(n_384),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_454),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_428),
.B(n_383),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_456),
.B(n_463),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_436),
.B(n_386),
.Y(n_457)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_457),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_419),
.A2(n_387),
.B1(n_400),
.B2(n_399),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_439),
.A2(n_389),
.B(n_406),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_402),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_409),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_437),
.B(n_407),
.C(n_395),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_364),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_466),
.B(n_436),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_391),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_468),
.B(n_475),
.Y(n_494)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_469),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_452),
.A2(n_417),
.B(n_438),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_471),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_472),
.A2(n_478),
.B1(n_485),
.B2(n_458),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_459),
.A2(n_432),
.B1(n_412),
.B2(n_420),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_473),
.A2(n_483),
.B1(n_489),
.B2(n_460),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_414),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_476),
.B(n_467),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_455),
.A2(n_416),
.B1(n_412),
.B2(n_418),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_457),
.B(n_410),
.Y(n_480)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_480),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_461),
.A2(n_435),
.B1(n_430),
.B2(n_413),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_450),
.A2(n_410),
.B1(n_413),
.B2(n_430),
.Y(n_485)
);

AOI21xp33_ASAP7_75t_L g486 ( 
.A1(n_462),
.A2(n_372),
.B(n_366),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_486),
.B(n_441),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_487),
.B(n_464),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_448),
.A2(n_378),
.B1(n_391),
.B2(n_354),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_496),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_443),
.C(n_445),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_498),
.C(n_507),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_470),
.Y(n_495)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_495),
.Y(n_510)
);

CKINVDCx14_ASAP7_75t_R g513 ( 
.A(n_497),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_443),
.C(n_445),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_469),
.Y(n_499)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_499),
.Y(n_512)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_484),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_506),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_501),
.B(n_504),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_L g502 ( 
.A(n_479),
.B(n_444),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_502),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_477),
.B(n_447),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_505),
.B(n_474),
.Y(n_521)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_480),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_477),
.B(n_446),
.C(n_449),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_503),
.A2(n_482),
.B1(n_475),
.B2(n_473),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_514),
.B(n_517),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_490),
.B(n_488),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_515),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_503),
.A2(n_481),
.B(n_471),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_516),
.B(n_519),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_491),
.A2(n_481),
.B(n_488),
.Y(n_517)
);

AND2x2_ASAP7_75t_SL g518 ( 
.A(n_507),
.B(n_483),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_518),
.B(n_521),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_494),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_513),
.A2(n_472),
.B1(n_485),
.B2(n_494),
.Y(n_524)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_524),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_493),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_525),
.B(n_527),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_498),
.C(n_492),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_512),
.A2(n_487),
.B1(n_489),
.B2(n_504),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_530),
.B(n_533),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_509),
.B(n_505),
.C(n_474),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_518),
.C(n_522),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_517),
.A2(n_352),
.B1(n_14),
.B2(n_15),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_532),
.A2(n_352),
.B1(n_516),
.B2(n_515),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_510),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_535),
.B(n_536),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_508),
.C(n_522),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_537),
.B(n_532),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_523),
.B(n_511),
.Y(n_538)
);

AOI31xp67_ASAP7_75t_SL g542 ( 
.A1(n_538),
.A2(n_528),
.A3(n_526),
.B(n_511),
.Y(n_542)
);

NOR3x1_ASAP7_75t_SL g546 ( 
.A(n_542),
.B(n_539),
.C(n_529),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_534),
.B(n_531),
.C(n_508),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_543),
.B(n_544),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_539),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_541),
.C(n_545),
.Y(n_548)
);

AOI21x1_ASAP7_75t_L g549 ( 
.A1(n_548),
.A2(n_540),
.B(n_518),
.Y(n_549)
);

OAI32xp33_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_524),
.A3(n_530),
.B1(n_352),
.B2(n_13),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_13),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_15),
.Y(n_552)
);


endmodule