module fake_jpeg_4649_n_78 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx16f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx10_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_20),
.B(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_16),
.B(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_14),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_14),
.Y(n_34)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_33),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_32),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_8),
.B(n_17),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_8),
.C(n_10),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_11),
.B1(n_12),
.B2(n_9),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_41),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_25),
.C(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_31),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_30),
.C(n_37),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_52),
.Y(n_60)
);

AOI322xp5_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_29),
.A3(n_8),
.B1(n_10),
.B2(n_23),
.C1(n_26),
.C2(n_14),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_20),
.C(n_8),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_55),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_23),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_13),
.B(n_23),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_61),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_13),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_20),
.C(n_26),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_10),
.C(n_14),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_23),
.B(n_14),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_10),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_56),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_10),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_69),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_3),
.C(n_5),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_10),
.B(n_1),
.C(n_0),
.Y(n_69)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_64),
.C(n_0),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_6),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_73),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_75),
.Y(n_78)
);


endmodule