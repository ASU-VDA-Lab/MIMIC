module fake_jpeg_25688_n_126 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_126);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx8_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_7),
.B(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_15),
.B1(n_18),
.B2(n_25),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_15),
.B1(n_18),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_28),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_27),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_32),
.B1(n_37),
.B2(n_45),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_62),
.B1(n_38),
.B2(n_45),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_33),
.B(n_23),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_38),
.B(n_14),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_56),
.Y(n_80)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_11),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_60),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx2_ASAP7_75t_SL g77 ( 
.A(n_58),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_64),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_20),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_66),
.B(n_56),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_57),
.B1(n_62),
.B2(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_22),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_19),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_83),
.Y(n_89)
);

BUFx24_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_73),
.B(n_2),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_92),
.B1(n_94),
.B2(n_21),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_55),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_87),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_70),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_56),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_91),
.C(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_67),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_65),
.B1(n_67),
.B2(n_16),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_17),
.B1(n_16),
.B2(n_19),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_77),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_97),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_75),
.B(n_78),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_101),
.B(n_102),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_73),
.C(n_81),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_88),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_2),
.B(n_17),
.Y(n_102)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_21),
.B(n_14),
.C(n_27),
.D(n_24),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_79),
.B1(n_21),
.B2(n_14),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_105),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_108),
.B(n_106),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_95),
.B1(n_92),
.B2(n_93),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_4),
.B(n_5),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_5),
.B(n_8),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_115),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_110),
.Y(n_115)
);

AOI21x1_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_103),
.B(n_21),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_116),
.A2(n_117),
.B(n_112),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_113),
.C(n_79),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_12),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_47),
.Y(n_123)
);

AO21x1_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_123),
.B(n_47),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_125),
.Y(n_126)
);


endmodule