module fake_jpeg_24722_n_243 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_14),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_28),
.B1(n_30),
.B2(n_21),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_45),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_37),
.B1(n_34),
.B2(n_18),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_23),
.B1(n_15),
.B2(n_17),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_19),
.B1(n_18),
.B2(n_29),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_59),
.B1(n_62),
.B2(n_31),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_27),
.B1(n_25),
.B2(n_15),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_18),
.B1(n_20),
.B2(n_26),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_38),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_20),
.B1(n_29),
.B2(n_26),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_33),
.A2(n_29),
.B1(n_20),
.B2(n_26),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_76),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_74),
.B1(n_82),
.B2(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_21),
.B1(n_23),
.B2(n_30),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_75),
.B1(n_80),
.B2(n_81),
.Y(n_94)
);

AOI22x1_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_42),
.B1(n_36),
.B2(n_32),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_23),
.B1(n_21),
.B2(n_27),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_79),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_42),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_31),
.B1(n_17),
.B2(n_15),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_33),
.B1(n_40),
.B2(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_32),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_35),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_46),
.Y(n_89)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_52),
.B1(n_48),
.B2(n_59),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_42),
.B1(n_36),
.B2(n_67),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_103),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_52),
.Y(n_97)
);

XOR2x2_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_104),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_47),
.B1(n_69),
.B2(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_51),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_17),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_1),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_65),
.B1(n_31),
.B2(n_17),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_112),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_113),
.B1(n_122),
.B2(n_97),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_98),
.B1(n_86),
.B2(n_128),
.Y(n_131)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_65),
.B1(n_40),
.B2(n_39),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_36),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_126),
.C(n_93),
.Y(n_129)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_104),
.A3(n_94),
.B1(n_90),
.B2(n_91),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_124),
.B(n_15),
.Y(n_149)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_127),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_87),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_120),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_85),
.B(n_25),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_88),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_129),
.B(n_110),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_93),
.B1(n_101),
.B2(n_86),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_149),
.B(n_150),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_95),
.C(n_103),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_132),
.B(n_144),
.Y(n_162)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_85),
.Y(n_136)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_87),
.Y(n_138)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_109),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_145),
.B(n_147),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_97),
.B1(n_105),
.B2(n_35),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_13),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_25),
.B1(n_3),
.B2(n_4),
.Y(n_150)
);

XNOR2x2_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_116),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_168),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_159),
.Y(n_175)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_123),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_145),
.C(n_134),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_166),
.C(n_133),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_107),
.B(n_112),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_124),
.Y(n_166)
);

NAND2x1_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_124),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_130),
.B1(n_137),
.B2(n_141),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_172),
.B1(n_151),
.B2(n_167),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_137),
.B1(n_141),
.B2(n_131),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_135),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_177),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_181),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_146),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_150),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_185),
.C(n_161),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_170),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_162),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_183),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_158),
.B(n_144),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_140),
.C(n_139),
.Y(n_185)
);

FAx1_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_25),
.CI(n_4),
.CON(n_186),
.SN(n_186)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_159),
.B(n_167),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_173),
.B1(n_156),
.B2(n_177),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_187),
.B1(n_186),
.B2(n_155),
.Y(n_204)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_201),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_165),
.Y(n_210)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_196),
.B(n_199),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_198),
.C(n_200),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_153),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_192),
.A2(n_160),
.B(n_186),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_205),
.A2(n_203),
.B(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_207),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_165),
.B1(n_184),
.B2(n_153),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_210),
.C(n_211),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_2),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_213),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_197),
.C(n_195),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_209),
.C(n_5),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_219),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_200),
.B(n_191),
.Y(n_219)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_191),
.B(n_4),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_2),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_210),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_7),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_225),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_227),
.A2(n_228),
.B(n_229),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_2),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_7),
.B(n_8),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_216),
.B1(n_222),
.B2(n_220),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_232),
.C(n_226),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_236)
);

OAI311xp33_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_234),
.A3(n_231),
.B1(n_11),
.C1(n_12),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_238),
.B(n_10),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_233),
.A2(n_9),
.B(n_10),
.Y(n_238)
);

BUFx24_ASAP7_75t_SL g241 ( 
.A(n_240),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_239),
.C(n_11),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_12),
.Y(n_243)
);


endmodule