module real_jpeg_25991_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_215;
wire n_288;
wire n_286;
wire n_292;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_299;
wire n_173;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_293;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_195;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_216;
wire n_179;
wire n_295;
wire n_167;
wire n_133;
wire n_244;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_21),
.B1(n_22),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_2),
.A2(n_29),
.B1(n_31),
.B2(n_68),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_2),
.A2(n_61),
.B1(n_63),
.B2(n_68),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_2),
.A2(n_68),
.B1(n_81),
.B2(n_82),
.Y(n_201)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_15),
.B(n_301),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_4),
.B(n_302),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_6),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_8),
.A2(n_20),
.B1(n_29),
.B2(n_31),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_8),
.A2(n_20),
.B1(n_61),
.B2(n_63),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_8),
.A2(n_20),
.B1(n_81),
.B2(n_82),
.Y(n_97)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_22),
.B1(n_28),
.B2(n_32),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_10),
.A2(n_23),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_10),
.A2(n_29),
.B1(n_31),
.B2(n_40),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_10),
.A2(n_40),
.B1(n_61),
.B2(n_63),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_10),
.A2(n_40),
.B1(n_81),
.B2(n_82),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_11),
.A2(n_22),
.B1(n_39),
.B2(n_51),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_11),
.A2(n_51),
.B1(n_61),
.B2(n_63),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_11),
.A2(n_29),
.B1(n_31),
.B2(n_51),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_11),
.A2(n_51),
.B1(n_81),
.B2(n_82),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_11),
.B(n_28),
.C(n_31),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_11),
.B(n_27),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_11),
.B(n_58),
.C(n_61),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_11),
.B(n_78),
.C(n_81),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_11),
.B(n_95),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_11),
.B(n_111),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_11),
.B(n_71),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_13),
.Y(n_93)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_13),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_43),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_41),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_35),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_19),
.A2(n_27),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_21),
.B(n_197),
.Y(n_196)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_26),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_27),
.A2(n_33),
.B1(n_50),
.B2(n_66),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_29),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_29),
.A2(n_31),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_31),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_36),
.B(n_45),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_48),
.B(n_49),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_84),
.B(n_300),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_46),
.B(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_46),
.B(n_298),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_52),
.CI(n_64),
.CON(n_46),
.SN(n_46)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_48),
.A2(n_49),
.B(n_67),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_56),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_60),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_55),
.A2(n_60),
.B(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_56),
.A2(n_71),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_56),
.B(n_116),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OA22x2_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_60),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_60),
.A2(n_115),
.B(n_126),
.Y(n_143)
);

INVx5_ASAP7_75t_SL g63 ( 
.A(n_61),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_63),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_61),
.B(n_243),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.C(n_72),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_65),
.B(n_134),
.C(n_142),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_65),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_65),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_65),
.A2(n_142),
.B1(n_143),
.B2(n_156),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_65),
.A2(n_113),
.B1(n_156),
.B2(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_65),
.B(n_113),
.C(n_194),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_69),
.A2(n_72),
.B1(n_123),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_69),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_72),
.A2(n_123),
.B1(n_124),
.B2(n_127),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_72),
.B(n_119),
.C(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_83),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_74),
.B(n_102),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_76),
.A2(n_102),
.B1(n_111),
.B2(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_80),
.A2(n_101),
.B(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_81),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_81),
.B(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_297),
.B(n_299),
.Y(n_84)
);

OAI211xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_144),
.B(n_158),
.C(n_296),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_128),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_87),
.B(n_128),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_106),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_88),
.B(n_108),
.C(n_117),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_98),
.B(n_103),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_89),
.A2(n_103),
.B1(n_104),
.B2(n_131),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_89),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_89),
.A2(n_99),
.B1(n_131),
.B2(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_97),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_91),
.B(n_202),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_97),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_92),
.B(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_92),
.Y(n_200)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_96),
.A2(n_136),
.B(n_171),
.Y(n_170)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_96),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_99),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_117),
.B2(n_118),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_109),
.B(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_113),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_113),
.B(n_214),
.C(n_216),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_113),
.A2(n_204),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_120),
.B1(n_152),
.B2(n_157),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_142),
.C(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_119),
.A2(n_120),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_119),
.A2(n_120),
.B1(n_176),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_120),
.B(n_168),
.C(n_176),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_120),
.B(n_148),
.C(n_152),
.Y(n_298)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_124),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.C(n_133),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_129),
.B(n_132),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_135),
.A2(n_139),
.B1(n_140),
.B2(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_135),
.Y(n_287)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_139),
.A2(n_140),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_139),
.A2(n_140),
.B1(n_227),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_140),
.B(n_221),
.C(n_227),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_140),
.B(n_199),
.C(n_258),
.Y(n_262)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_142),
.A2(n_143),
.B1(n_190),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_142),
.A2(n_143),
.B1(n_174),
.B2(n_187),
.Y(n_264)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_143),
.B(n_174),
.C(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_SL g158 ( 
.A(n_145),
.B(n_159),
.C(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_146),
.B(n_147),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_153),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_180),
.B(n_295),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_178),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_162),
.B(n_178),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_167),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_163),
.B(n_165),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_167),
.B(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_168),
.A2(n_169),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_174),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_170),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_172),
.A2(n_201),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_174),
.A2(n_187),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_174),
.B(n_244),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_176),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_290),
.B(n_294),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_217),
.B(n_276),
.C(n_289),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_206),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_183),
.B(n_206),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_193),
.B2(n_205),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_186),
.B(n_192),
.C(n_205),
.Y(n_277)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_203),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_198),
.A2(n_199),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_199),
.B(n_250),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_212),
.C(n_213),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_207),
.A2(n_208),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_213),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_216),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_214),
.B(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_216),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_275),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_236),
.B(n_274),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_233),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_220),
.B(n_233),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_221),
.A2(n_222),
.B1(n_270),
.B2(n_272),
.Y(n_269)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_226),
.B(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_227),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_267),
.B(n_273),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_261),
.B(n_266),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_253),
.B(n_260),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_245),
.B(n_252),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_242),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_249),
.B(n_251),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_254),
.B(n_255),
.Y(n_260)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_258),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_268),
.B(n_269),
.Y(n_273)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_270),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_278),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_288),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_285),
.B2(n_286),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_286),
.C(n_288),
.Y(n_291)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);


endmodule