module fake_ariane_3037_n_1953 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1953);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1953;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1865;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g185 ( 
.A(n_4),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_128),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_129),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_57),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_0),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_133),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_138),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_62),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_26),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_18),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_36),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_34),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_36),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_44),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_7),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_38),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_135),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_92),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_21),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_19),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_146),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_43),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_181),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_143),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_120),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_65),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_39),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_145),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_55),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_10),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_122),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_68),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_153),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_134),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_28),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_109),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_78),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_79),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_90),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_98),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_117),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_148),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_70),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_126),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_176),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_184),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_1),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_157),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_72),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_93),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_21),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_11),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_32),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_30),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_104),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_33),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_31),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_23),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_94),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_39),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_7),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_69),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_141),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_144),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_64),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_1),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_165),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_162),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_156),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_106),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_63),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_42),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_41),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_42),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_114),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_47),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_26),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_147),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_40),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_74),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_182),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_10),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_84),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_100),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_52),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_46),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_52),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_8),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_127),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_85),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_11),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_53),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_61),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_45),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_116),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_172),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_33),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_103),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_108),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_140),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_161),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_53),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_9),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_8),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_6),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_80),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_150),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_163),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_16),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_46),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_51),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_169),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_30),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_178),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_20),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_54),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_3),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_152),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_43),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_183),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_14),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_166),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_99),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_137),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_124),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_164),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_17),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_97),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_18),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_168),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_171),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_48),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_83),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_41),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_37),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_158),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_16),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_9),
.Y(n_325)
);

BUFx5_ASAP7_75t_L g326 ( 
.A(n_48),
.Y(n_326)
);

BUFx10_ASAP7_75t_L g327 ( 
.A(n_75),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_89),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_86),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_111),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_160),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_76),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_32),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_22),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_73),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_110),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_173),
.Y(n_337)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_132),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_24),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_6),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_149),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_151),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_22),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_31),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_20),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_4),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_5),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_17),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_67),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_77),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_27),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_5),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_60),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_91),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_37),
.Y(n_355)
);

CKINVDCx11_ASAP7_75t_R g356 ( 
.A(n_101),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_130),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_24),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_82),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_25),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_34),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_29),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_55),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_115),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_136),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_139),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_38),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_246),
.B(n_0),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_356),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_326),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_306),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_292),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_326),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_195),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_206),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_306),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_247),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_326),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_186),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_326),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

INVxp33_ASAP7_75t_SL g383 ( 
.A(n_198),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_247),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_247),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_326),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_247),
.Y(n_387)
);

INVxp33_ASAP7_75t_SL g388 ( 
.A(n_198),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_253),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_253),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_253),
.Y(n_391)
);

INVxp33_ASAP7_75t_SL g392 ( 
.A(n_200),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_186),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_214),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_253),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_266),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_R g397 ( 
.A(n_191),
.B(n_71),
.Y(n_397)
);

BUFx6f_ASAP7_75t_SL g398 ( 
.A(n_221),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_204),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_191),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_197),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_266),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_288),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_200),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_266),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_217),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_222),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_266),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_197),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_199),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_199),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_241),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_210),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_210),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_305),
.B(n_2),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_234),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_194),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_241),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_239),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_298),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_218),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_205),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_243),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_L g424 ( 
.A(n_216),
.B(n_2),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_196),
.B(n_3),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_298),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_244),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_224),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_248),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_224),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_185),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_225),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_260),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_261),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_218),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_263),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_215),
.B(n_12),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_225),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_269),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_189),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_277),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_272),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_277),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_223),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_252),
.B(n_12),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_201),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_209),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_295),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_273),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_295),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_232),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_268),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_262),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_265),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_L g455 ( 
.A(n_238),
.B(n_13),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_317),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_267),
.B(n_13),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_285),
.B(n_14),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_377),
.B(n_336),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_379),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_370),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_369),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_R g464 ( 
.A(n_374),
.B(n_202),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_393),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_400),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_373),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_413),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_414),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_373),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_447),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_384),
.B(n_293),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_399),
.B(n_221),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_385),
.B(n_294),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_421),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_378),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_435),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_378),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_417),
.B(n_444),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_447),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_451),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_380),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_380),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_381),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_447),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_452),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_418),
.B(n_205),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_381),
.A2(n_337),
.B(n_317),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_382),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_382),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_386),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_428),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_R g494 ( 
.A(n_394),
.B(n_268),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_428),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_430),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_430),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_406),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_407),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_417),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_389),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_395),
.B(n_299),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_372),
.B(n_328),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_404),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_440),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_432),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_432),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_438),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_399),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_441),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_416),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_419),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_R g514 ( 
.A(n_423),
.B(n_331),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_441),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_443),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_398),
.B(n_301),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_389),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_427),
.Y(n_519)
);

OA21x2_ASAP7_75t_L g520 ( 
.A1(n_445),
.A2(n_309),
.B(n_307),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_403),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_444),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_443),
.B(n_337),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_387),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_371),
.B(n_205),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_448),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_376),
.B(n_274),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_387),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_390),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_450),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_450),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_429),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_390),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_433),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_459),
.B(n_405),
.Y(n_537)
);

INVxp33_ASAP7_75t_L g538 ( 
.A(n_505),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_459),
.B(n_403),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_520),
.A2(n_500),
.B1(n_479),
.B2(n_375),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_471),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_480),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_536),
.B(n_422),
.Y(n_543)
);

BUFx10_ASAP7_75t_L g544 ( 
.A(n_498),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_480),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_499),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_467),
.B(n_478),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_500),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_500),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_480),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_536),
.B(n_415),
.Y(n_551)
);

INVx4_ASAP7_75t_SL g552 ( 
.A(n_523),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_471),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_471),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_467),
.B(n_478),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_479),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_494),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_517),
.B(n_434),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_514),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_504),
.B(n_436),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_479),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_487),
.B(n_439),
.Y(n_562)
);

CKINVDCx6p67_ASAP7_75t_R g563 ( 
.A(n_510),
.Y(n_563)
);

AND2x6_ASAP7_75t_L g564 ( 
.A(n_487),
.B(n_366),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_483),
.B(n_398),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_512),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_480),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_485),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_483),
.B(n_398),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_484),
.B(n_442),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_484),
.B(n_449),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_489),
.B(n_383),
.Y(n_572)
);

BUFx10_ASAP7_75t_L g573 ( 
.A(n_513),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_527),
.B(n_401),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_460),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_489),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_491),
.B(n_388),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_465),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_479),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_527),
.B(n_409),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_491),
.B(n_392),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_519),
.B(n_331),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_485),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_471),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_492),
.B(n_471),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_485),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_529),
.B(n_431),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_493),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_493),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_485),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_492),
.B(n_311),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_495),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_461),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_521),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_L g595 ( 
.A(n_461),
.B(n_397),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_529),
.B(n_453),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_503),
.B(n_472),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_495),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_461),
.Y(n_599)
);

BUFx10_ASAP7_75t_L g600 ( 
.A(n_463),
.Y(n_600)
);

INVxp67_ASAP7_75t_SL g601 ( 
.A(n_471),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_534),
.B(n_446),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_462),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_496),
.Y(n_604)
);

OAI22xp33_ASAP7_75t_L g605 ( 
.A1(n_464),
.A2(n_322),
.B1(n_189),
.B2(n_275),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_462),
.B(n_315),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_518),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_462),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_520),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_473),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_472),
.B(n_424),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_470),
.B(n_323),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_470),
.Y(n_613)
);

AND2x6_ASAP7_75t_L g614 ( 
.A(n_470),
.B(n_366),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_476),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_466),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_476),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_496),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_468),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_474),
.B(n_398),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_497),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_476),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_469),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_482),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_518),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_477),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_520),
.Y(n_627)
);

AND2x2_ASAP7_75t_SL g628 ( 
.A(n_520),
.B(n_368),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_482),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_482),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_497),
.Y(n_631)
);

BUFx6f_ASAP7_75t_SL g632 ( 
.A(n_523),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_474),
.B(n_454),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_502),
.B(n_454),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_490),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_522),
.B(n_410),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_490),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_502),
.B(n_456),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_490),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_475),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_522),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_522),
.Y(n_642)
);

INVx4_ASAP7_75t_SL g643 ( 
.A(n_523),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_506),
.Y(n_644)
);

INVx4_ASAP7_75t_SL g645 ( 
.A(n_523),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_522),
.B(n_424),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_525),
.B(n_341),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_524),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_525),
.B(n_455),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_525),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_524),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_506),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_518),
.Y(n_653)
);

BUFx8_ASAP7_75t_SL g654 ( 
.A(n_486),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_525),
.B(n_353),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_507),
.Y(n_656)
);

AND2x6_ASAP7_75t_L g657 ( 
.A(n_507),
.B(n_359),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_508),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_524),
.Y(n_659)
);

AND2x2_ASAP7_75t_SL g660 ( 
.A(n_508),
.B(n_425),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_523),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_509),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_509),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_511),
.B(n_515),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_511),
.B(n_455),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_523),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_515),
.B(n_203),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_516),
.B(n_410),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_516),
.A2(n_458),
.B1(n_457),
.B2(n_437),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g670 ( 
.A(n_526),
.B(n_208),
.C(n_202),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_526),
.B(n_411),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_528),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_528),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_481),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_532),
.B(n_456),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_518),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_532),
.B(n_533),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_533),
.B(n_203),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_531),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_523),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_523),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_531),
.B(n_411),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_488),
.B(n_207),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_531),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_535),
.B(n_391),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_488),
.B(n_207),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_518),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_488),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_628),
.B(n_354),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_560),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_597),
.B(n_270),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_633),
.B(n_312),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_582),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_562),
.B(n_354),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_566),
.B(n_535),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_633),
.B(n_320),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_570),
.B(n_281),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_654),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_628),
.A2(n_275),
.B1(n_322),
.B2(n_348),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_565),
.B(n_357),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_613),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_564),
.A2(n_357),
.B1(n_348),
.B2(n_361),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_537),
.B(n_611),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_613),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_611),
.B(n_535),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_575),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_565),
.B(n_209),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_601),
.A2(n_501),
.B(n_188),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_569),
.B(n_209),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_611),
.B(n_289),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_620),
.B(n_297),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_539),
.B(n_193),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_622),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_572),
.B(n_264),
.C(n_259),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_620),
.B(n_303),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_555),
.A2(n_501),
.B(n_190),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_569),
.B(n_209),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_576),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_638),
.B(n_304),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_576),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_622),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_615),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_615),
.Y(n_723)
);

NOR3xp33_ASAP7_75t_L g724 ( 
.A(n_572),
.B(n_351),
.C(n_245),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_636),
.Y(n_725)
);

NOR2xp67_ASAP7_75t_L g726 ( 
.A(n_616),
.B(n_412),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_654),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_638),
.B(n_316),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_543),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_602),
.B(n_558),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_564),
.A2(n_251),
.B1(n_280),
.B2(n_365),
.Y(n_731)
);

OR2x6_ASAP7_75t_L g732 ( 
.A(n_619),
.B(n_420),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_664),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_615),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_557),
.B(n_208),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_564),
.B(n_319),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_571),
.B(n_291),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_617),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_564),
.B(n_334),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_544),
.B(n_291),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_595),
.B(n_581),
.C(n_577),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_564),
.B(n_340),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_617),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_657),
.A2(n_339),
.B1(n_333),
.B2(n_325),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_617),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_554),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_661),
.B(n_209),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_596),
.B(n_343),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_661),
.B(n_209),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_634),
.B(n_344),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_660),
.B(n_346),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_660),
.B(n_347),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_574),
.B(n_274),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_593),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_538),
.B(n_274),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_577),
.B(n_352),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_661),
.B(n_209),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_593),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_581),
.B(n_240),
.C(n_278),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_587),
.B(n_362),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_666),
.B(n_338),
.Y(n_761)
);

BUFx5_ASAP7_75t_L g762 ( 
.A(n_688),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_610),
.B(n_363),
.Y(n_763)
);

BUFx5_ASAP7_75t_L g764 ( 
.A(n_688),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_657),
.A2(n_367),
.B1(n_321),
.B2(n_324),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_665),
.B(n_279),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_555),
.A2(n_585),
.B(n_547),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_554),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_585),
.A2(n_501),
.B(n_229),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_599),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_599),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_666),
.B(n_338),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_666),
.B(n_338),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_667),
.B(n_678),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_603),
.Y(n_775)
);

AO221x1_ASAP7_75t_L g776 ( 
.A1(n_605),
.A2(n_345),
.B1(n_314),
.B2(n_284),
.C(n_290),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_665),
.B(n_296),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_677),
.B(n_302),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_667),
.B(n_300),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_657),
.A2(n_308),
.B1(n_327),
.B2(n_221),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_680),
.B(n_338),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_548),
.Y(n_782)
);

AND2x6_ASAP7_75t_L g783 ( 
.A(n_603),
.B(n_518),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_538),
.B(n_420),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_677),
.B(n_300),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_669),
.A2(n_355),
.B1(n_358),
.B2(n_360),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_559),
.B(n_426),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_540),
.B(n_355),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_678),
.B(n_641),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_680),
.B(n_338),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_668),
.B(n_426),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_549),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_554),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_680),
.B(n_338),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_556),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_580),
.B(n_358),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_561),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_641),
.B(n_360),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_579),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_649),
.B(n_187),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_595),
.A2(n_212),
.B1(n_364),
.B2(n_350),
.Y(n_801)
);

NOR3xp33_ASAP7_75t_L g802 ( 
.A(n_626),
.B(n_391),
.C(n_408),
.Y(n_802)
);

BUFx8_ASAP7_75t_L g803 ( 
.A(n_594),
.Y(n_803)
);

OR2x6_ASAP7_75t_L g804 ( 
.A(n_543),
.B(n_530),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_608),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_641),
.B(n_276),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_L g807 ( 
.A(n_657),
.B(n_338),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_608),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_649),
.B(n_192),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_681),
.B(n_530),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_L g811 ( 
.A1(n_668),
.A2(n_408),
.B1(n_402),
.B2(n_396),
.Y(n_811)
);

A2O1A1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_547),
.A2(n_402),
.B(n_396),
.C(n_530),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_544),
.B(n_276),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_624),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_544),
.B(n_276),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_588),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_649),
.B(n_211),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_589),
.A2(n_15),
.B(n_19),
.C(n_25),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_592),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_642),
.B(n_327),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_646),
.B(n_213),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_600),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_624),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_578),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_657),
.A2(n_327),
.B1(n_530),
.B2(n_342),
.Y(n_825)
);

O2A1O1Ixp5_ASAP7_75t_L g826 ( 
.A1(n_683),
.A2(n_256),
.B(n_349),
.C(n_335),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_598),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_604),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_618),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_646),
.B(n_219),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_621),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_646),
.B(n_220),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_631),
.B(n_226),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_681),
.B(n_530),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_668),
.A2(n_257),
.B1(n_332),
.B2(n_330),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_644),
.B(n_227),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_551),
.A2(n_255),
.B1(n_329),
.B2(n_318),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_629),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_629),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_681),
.B(n_530),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_652),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_656),
.B(n_658),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_662),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_663),
.B(n_313),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_554),
.B(n_310),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_674),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_551),
.B(n_15),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_609),
.A2(n_287),
.B1(n_286),
.B2(n_283),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_672),
.B(n_282),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_673),
.B(n_271),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_642),
.B(n_258),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_675),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_671),
.B(n_254),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_630),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_642),
.B(n_250),
.Y(n_855)
);

NAND2x1_ASAP7_75t_L g856 ( 
.A(n_650),
.B(n_112),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_609),
.A2(n_249),
.B1(n_242),
.B2(n_237),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_630),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_774),
.A2(n_545),
.B(n_590),
.C(n_550),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_733),
.A2(n_551),
.B1(n_671),
.B2(n_650),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_767),
.A2(n_686),
.B(n_683),
.Y(n_861)
);

AND2x6_ASAP7_75t_L g862 ( 
.A(n_847),
.B(n_671),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_851),
.A2(n_686),
.B(n_584),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_732),
.Y(n_864)
);

OAI21x1_ASAP7_75t_L g865 ( 
.A1(n_856),
.A2(n_637),
.B(n_635),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_822),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_851),
.A2(n_584),
.B(n_553),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_855),
.A2(n_584),
.B(n_553),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_786),
.A2(n_591),
.B(n_545),
.C(n_550),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_795),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_804),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_699),
.A2(n_650),
.B1(n_542),
.B2(n_590),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_691),
.B(n_542),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_774),
.A2(n_567),
.B(n_586),
.C(n_583),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_779),
.A2(n_567),
.B(n_586),
.C(n_583),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_855),
.A2(n_553),
.B(n_541),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_747),
.A2(n_541),
.B(n_568),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_747),
.A2(n_541),
.B(n_568),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_749),
.A2(n_635),
.B(n_637),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_846),
.B(n_546),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_749),
.A2(n_761),
.B(n_757),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_746),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_692),
.B(n_546),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_696),
.B(n_546),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_741),
.A2(n_627),
.B(n_609),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_SL g886 ( 
.A1(n_789),
.A2(n_591),
.B(n_639),
.C(n_612),
.Y(n_886)
);

AO21x2_ASAP7_75t_L g887 ( 
.A1(n_707),
.A2(n_612),
.B(n_606),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_730),
.B(n_573),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_746),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_796),
.B(n_573),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_690),
.B(n_573),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_757),
.A2(n_639),
.B(n_687),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_712),
.B(n_682),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_701),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_761),
.A2(n_687),
.B(n_627),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_772),
.A2(n_687),
.B(n_627),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_753),
.B(n_600),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_712),
.B(n_682),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_719),
.B(n_679),
.Y(n_899)
);

CKINVDCx6p67_ASAP7_75t_R g900 ( 
.A(n_727),
.Y(n_900)
);

AO21x1_ASAP7_75t_L g901 ( 
.A1(n_707),
.A2(n_606),
.B(n_684),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_772),
.A2(n_647),
.B(n_655),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_824),
.Y(n_903)
);

NOR3xp33_ASAP7_75t_L g904 ( 
.A(n_756),
.B(n_640),
.C(n_623),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_773),
.A2(n_647),
.B(n_655),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_789),
.A2(n_670),
.B(n_659),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_732),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_791),
.B(n_643),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_700),
.B(n_600),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_702),
.B(n_625),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_746),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_728),
.B(n_651),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_703),
.B(n_651),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_746),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_704),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_773),
.A2(n_659),
.B(n_648),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_781),
.A2(n_648),
.B(n_676),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_781),
.A2(n_607),
.B(n_676),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_699),
.A2(n_685),
.B1(n_563),
.B2(n_632),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_784),
.B(n_552),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_790),
.A2(n_676),
.B(n_653),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_L g922 ( 
.A(n_756),
.B(n_676),
.C(n_653),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_732),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_852),
.B(n_653),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_804),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_785),
.B(n_653),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_797),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_725),
.B(n_625),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_755),
.B(n_645),
.Y(n_929)
);

INVx11_ASAP7_75t_L g930 ( 
.A(n_803),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_689),
.A2(n_779),
.B1(n_798),
.B2(n_820),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_791),
.B(n_607),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_790),
.A2(n_607),
.B(n_625),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_798),
.B(n_625),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_806),
.A2(n_607),
.B(n_228),
.C(n_235),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_711),
.B(n_614),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_794),
.A2(n_230),
.B(n_231),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_715),
.B(n_614),
.Y(n_938)
);

BUFx12f_ASAP7_75t_L g939 ( 
.A(n_698),
.Y(n_939)
);

INVx11_ASAP7_75t_L g940 ( 
.A(n_803),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_713),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_768),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_794),
.A2(n_236),
.B(n_233),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_787),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_729),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_693),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_750),
.B(n_614),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_806),
.B(n_614),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_820),
.B(n_614),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_816),
.B(n_645),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_694),
.B(n_632),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_751),
.A2(n_643),
.B(n_552),
.C(n_29),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_810),
.A2(n_643),
.B(n_552),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_810),
.A2(n_96),
.B(n_179),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_834),
.A2(n_95),
.B(n_177),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_834),
.A2(n_88),
.B(n_175),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_819),
.B(n_27),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_840),
.A2(n_87),
.B(n_174),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_752),
.B(n_28),
.Y(n_959)
);

BUFx4f_ASAP7_75t_L g960 ( 
.A(n_804),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_799),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_689),
.A2(n_35),
.B1(n_40),
.B2(n_44),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_737),
.B(n_35),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_840),
.A2(n_105),
.B(n_170),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_812),
.A2(n_826),
.B(n_842),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_709),
.A2(n_102),
.B(n_167),
.Y(n_966)
);

OAI321xp33_ASAP7_75t_L g967 ( 
.A1(n_780),
.A2(n_45),
.A3(n_47),
.B1(n_49),
.B2(n_50),
.C(n_51),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_722),
.A2(n_49),
.B(n_50),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_726),
.B(n_54),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_709),
.A2(n_717),
.B(n_743),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_768),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_723),
.A2(n_56),
.B(n_58),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_763),
.B(n_180),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_721),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_760),
.B(n_59),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_827),
.B(n_828),
.Y(n_976)
);

OAI21xp33_ASAP7_75t_L g977 ( 
.A1(n_778),
.A2(n_66),
.B(n_81),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_717),
.A2(n_107),
.B(n_113),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_748),
.A2(n_118),
.B(n_121),
.C(n_123),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_763),
.B(n_125),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_829),
.B(n_159),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_768),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_831),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_754),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_734),
.A2(n_142),
.B(n_154),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_695),
.B(n_835),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_762),
.B(n_764),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_740),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_738),
.A2(n_745),
.B(n_841),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_762),
.B(n_764),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_843),
.B(n_718),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_780),
.A2(n_724),
.B1(n_714),
.B2(n_857),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_762),
.B(n_764),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_818),
.A2(n_720),
.B(n_782),
.C(n_792),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_697),
.A2(n_844),
.B(n_836),
.C(n_833),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_788),
.A2(n_776),
.B1(n_744),
.B2(n_765),
.Y(n_996)
);

O2A1O1Ixp5_ASAP7_75t_L g997 ( 
.A1(n_845),
.A2(n_708),
.B(n_849),
.C(n_850),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_762),
.B(n_764),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_758),
.B(n_858),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_L g1000 ( 
.A(n_848),
.B(n_857),
.C(n_765),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_SL g1001 ( 
.A1(n_845),
.A2(n_853),
.B(n_742),
.C(n_739),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_766),
.B(n_777),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_744),
.A2(n_848),
.B1(n_825),
.B2(n_731),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_759),
.A2(n_710),
.B1(n_801),
.B2(n_821),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_770),
.B(n_854),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_768),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_735),
.B(n_813),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_830),
.A2(n_832),
.B(n_817),
.Y(n_1008)
);

AOI22x1_ASAP7_75t_L g1009 ( 
.A1(n_771),
.A2(n_805),
.B1(n_838),
.B2(n_823),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_716),
.A2(n_814),
.B(n_808),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_800),
.A2(n_809),
.B(n_807),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_825),
.A2(n_705),
.B1(n_837),
.B2(n_736),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_793),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_775),
.A2(n_839),
.B(n_793),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_811),
.B(n_802),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_793),
.A2(n_769),
.B(n_764),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_811),
.B(n_793),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_783),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_815),
.B(n_762),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_783),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_762),
.B(n_764),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_783),
.A2(n_767),
.B(n_851),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_783),
.A2(n_767),
.B(n_851),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_783),
.A2(n_733),
.B1(n_699),
.B2(n_774),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_706),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_795),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_691),
.B(n_597),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_767),
.A2(n_855),
.B(n_851),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_846),
.B(n_379),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_767),
.A2(n_686),
.B(n_683),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_691),
.B(n_597),
.Y(n_1031)
);

INVx4_ASAP7_75t_L g1032 ( 
.A(n_822),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_699),
.A2(n_689),
.B1(n_628),
.B2(n_702),
.Y(n_1033)
);

OAI22x1_ASAP7_75t_L g1034 ( 
.A1(n_702),
.A2(n_440),
.B1(n_847),
.B2(n_689),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_796),
.B(n_574),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_846),
.B(n_379),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_767),
.A2(n_855),
.B(n_851),
.Y(n_1037)
);

AO21x1_ASAP7_75t_L g1038 ( 
.A1(n_707),
.A2(n_717),
.B(n_709),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_822),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_767),
.A2(n_855),
.B(n_851),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_846),
.B(n_379),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_690),
.B(n_566),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_689),
.A2(n_700),
.B1(n_741),
.B2(n_712),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_846),
.B(n_379),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_691),
.B(n_597),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_767),
.A2(n_686),
.B(n_683),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_691),
.B(n_597),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_908),
.B(n_871),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_931),
.A2(n_973),
.B(n_959),
.C(n_1043),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_865),
.A2(n_1016),
.B(n_861),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_1021),
.A2(n_934),
.B(n_1028),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_987),
.A2(n_993),
.B(n_990),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_998),
.A2(n_1023),
.B(n_1022),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1027),
.B(n_1031),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1030),
.A2(n_1046),
.B(n_885),
.Y(n_1055)
);

AO31x2_ASAP7_75t_L g1056 ( 
.A1(n_901),
.A2(n_1038),
.A3(n_1012),
.B(n_1003),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_862),
.A2(n_880),
.B1(n_992),
.B2(n_909),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_SL g1058 ( 
.A(n_1000),
.B(n_960),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1030),
.A2(n_1046),
.B(n_885),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_970),
.A2(n_863),
.B(n_1010),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_1045),
.A2(n_1047),
.B(n_898),
.C(n_893),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_SL g1062 ( 
.A1(n_1033),
.A2(n_962),
.B(n_963),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1037),
.A2(n_1040),
.B(n_949),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1024),
.B(n_899),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_1010),
.A2(n_896),
.B(n_895),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_948),
.A2(n_912),
.B(n_995),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1024),
.A2(n_976),
.B1(n_1003),
.B2(n_980),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_960),
.B(n_871),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_1008),
.A2(n_1004),
.B(n_975),
.C(n_994),
.Y(n_1069)
);

AOI221x1_ASAP7_75t_L g1070 ( 
.A1(n_1012),
.A2(n_1034),
.B1(n_977),
.B2(n_860),
.C(n_968),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_900),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_913),
.B(n_862),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_991),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_859),
.A2(n_874),
.B(n_881),
.Y(n_1074)
);

AO31x2_ASAP7_75t_L g1075 ( 
.A1(n_875),
.A2(n_947),
.A3(n_936),
.B(n_938),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_879),
.A2(n_916),
.B(n_917),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_944),
.B(n_1035),
.Y(n_1077)
);

AND3x4_ASAP7_75t_L g1078 ( 
.A(n_904),
.B(n_940),
.C(n_930),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_918),
.A2(n_933),
.B(n_921),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_983),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_883),
.B(n_884),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_870),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_926),
.A2(n_1011),
.B(n_878),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_906),
.A2(n_892),
.B(n_877),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_864),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_927),
.Y(n_1086)
);

OR2x6_ASAP7_75t_L g1087 ( 
.A(n_908),
.B(n_925),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_984),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_867),
.A2(n_868),
.B(n_876),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_862),
.B(n_1002),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_1029),
.B(n_1036),
.Y(n_1091)
);

AOI21xp33_ASAP7_75t_L g1092 ( 
.A1(n_919),
.A2(n_1015),
.B(n_860),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_897),
.B(n_890),
.Y(n_1093)
);

BUFx8_ASAP7_75t_L g1094 ( 
.A(n_939),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1014),
.A2(n_1009),
.B(n_989),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_873),
.A2(n_1001),
.B(n_886),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_889),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_907),
.B(n_923),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_872),
.A2(n_952),
.A3(n_935),
.B(n_902),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1041),
.B(n_1044),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_989),
.A2(n_981),
.B(n_997),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_L g1102 ( 
.A1(n_986),
.A2(n_965),
.B(n_906),
.C(n_969),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_862),
.B(n_961),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_888),
.B(n_891),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_1007),
.A2(n_967),
.B(n_869),
.C(n_968),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_872),
.A2(n_905),
.A3(n_919),
.B(n_999),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_925),
.B(n_866),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_924),
.A2(n_928),
.B(n_965),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_1020),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_972),
.A2(n_922),
.B(n_950),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_862),
.B(n_1026),
.Y(n_1111)
);

OAI21xp33_ASAP7_75t_L g1112 ( 
.A1(n_957),
.A2(n_996),
.B(n_1042),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_999),
.A2(n_1005),
.A3(n_1017),
.B(n_966),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_972),
.A2(n_1019),
.B(n_882),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_979),
.A2(n_951),
.B(n_978),
.C(n_955),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1018),
.A2(n_954),
.B(n_956),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1018),
.A2(n_964),
.B(n_958),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_903),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_882),
.A2(n_942),
.B(n_1013),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_946),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_866),
.B(n_1039),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1005),
.A2(n_985),
.B(n_1013),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_932),
.A2(n_929),
.B(n_920),
.C(n_910),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_894),
.B(n_941),
.Y(n_1124)
);

BUFx12f_ASAP7_75t_L g1125 ( 
.A(n_1032),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_915),
.B(n_974),
.Y(n_1126)
);

INVx5_ASAP7_75t_L g1127 ( 
.A(n_1020),
.Y(n_1127)
);

NOR2x1_ASAP7_75t_L g1128 ( 
.A(n_1032),
.B(n_1039),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_945),
.B(n_988),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_971),
.A2(n_982),
.B(n_953),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_937),
.A2(n_943),
.B(n_1020),
.C(n_911),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_889),
.B(n_911),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_887),
.A2(n_889),
.B(n_911),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_914),
.A2(n_1021),
.B(n_934),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1006),
.B(n_944),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1006),
.B(n_944),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1021),
.A2(n_934),
.B(n_1028),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1025),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_901),
.A2(n_1038),
.A3(n_861),
.B(n_1021),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_865),
.A2(n_1016),
.B(n_861),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_944),
.B(n_1035),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_991),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_908),
.B(n_871),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_930),
.Y(n_1144)
);

AO21x1_ASAP7_75t_L g1145 ( 
.A1(n_931),
.A2(n_973),
.B(n_1003),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1021),
.A2(n_934),
.B(n_1028),
.Y(n_1146)
);

AO22x1_ASAP7_75t_L g1147 ( 
.A1(n_880),
.A2(n_616),
.B1(n_468),
.B2(n_469),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_865),
.A2(n_1016),
.B(n_861),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_991),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_865),
.A2(n_1016),
.B(n_861),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1027),
.B(n_1031),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_864),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_931),
.A2(n_893),
.B1(n_898),
.B2(n_1000),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_L g1154 ( 
.A1(n_1035),
.A2(n_605),
.B1(n_699),
.B2(n_786),
.C(n_375),
.Y(n_1154)
);

NOR3xp33_ASAP7_75t_L g1155 ( 
.A(n_883),
.B(n_566),
.C(n_536),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_1025),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_931),
.A2(n_973),
.B(n_959),
.C(n_774),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_862),
.A2(n_582),
.B1(n_566),
.B2(n_699),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_861),
.A2(n_1046),
.B(n_1030),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_930),
.Y(n_1160)
);

O2A1O1Ixp5_ASAP7_75t_L g1161 ( 
.A1(n_973),
.A2(n_959),
.B(n_1011),
.C(n_1028),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_944),
.B(n_1035),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_865),
.A2(n_1016),
.B(n_861),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_931),
.A2(n_973),
.B(n_959),
.C(n_774),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_991),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1021),
.A2(n_934),
.B(n_1028),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1021),
.A2(n_934),
.B(n_1028),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_931),
.A2(n_893),
.B1(n_898),
.B2(n_1000),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_880),
.B(n_582),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_960),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1027),
.B(n_379),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1021),
.A2(n_934),
.B(n_1028),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_960),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1027),
.B(n_379),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1027),
.B(n_379),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_861),
.A2(n_1046),
.B(n_1030),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1027),
.B(n_1031),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_865),
.A2(n_1016),
.B(n_861),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_SL g1179 ( 
.A1(n_931),
.A2(n_1033),
.B(n_699),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_984),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_944),
.B(n_1035),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1027),
.B(n_1031),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1027),
.B(n_1031),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_865),
.A2(n_1016),
.B(n_861),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_880),
.B(n_582),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_901),
.A2(n_1038),
.A3(n_861),
.B(n_1021),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1021),
.A2(n_934),
.B(n_1028),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1027),
.B(n_1031),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_865),
.A2(n_1016),
.B(n_861),
.Y(n_1189)
);

AOI21x1_ASAP7_75t_L g1190 ( 
.A1(n_861),
.A2(n_1037),
.B(n_1028),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1020),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1021),
.A2(n_934),
.B(n_1028),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_931),
.A2(n_973),
.B(n_959),
.C(n_774),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_865),
.A2(n_1016),
.B(n_861),
.Y(n_1194)
);

INVx2_ASAP7_75t_SL g1195 ( 
.A(n_930),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_861),
.A2(n_1046),
.B(n_1030),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_865),
.A2(n_1016),
.B(n_861),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_901),
.A2(n_1038),
.A3(n_861),
.B(n_1021),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_908),
.B(n_871),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_865),
.A2(n_1016),
.B(n_861),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1021),
.A2(n_934),
.B(n_1028),
.Y(n_1201)
);

AOI221xp5_ASAP7_75t_SL g1202 ( 
.A1(n_968),
.A2(n_1031),
.B1(n_1045),
.B2(n_1027),
.C(n_1047),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1020),
.Y(n_1203)
);

AO21x1_ASAP7_75t_L g1204 ( 
.A1(n_931),
.A2(n_973),
.B(n_1003),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_984),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1088),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1157),
.A2(n_1164),
.B1(n_1193),
.B2(n_1049),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1161),
.A2(n_1204),
.B(n_1145),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1153),
.A2(n_1168),
.B(n_1069),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1054),
.B(n_1151),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1153),
.A2(n_1168),
.B(n_1137),
.Y(n_1211)
);

NOR2xp67_ASAP7_75t_L g1212 ( 
.A(n_1144),
.B(n_1160),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1077),
.B(n_1141),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1051),
.A2(n_1166),
.B(n_1146),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1080),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1106),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1127),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1054),
.B(n_1151),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1180),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1162),
.B(n_1181),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1177),
.B(n_1182),
.Y(n_1221)
);

AND2x2_ASAP7_75t_SL g1222 ( 
.A(n_1058),
.B(n_1064),
.Y(n_1222)
);

BUFx12f_ASAP7_75t_L g1223 ( 
.A(n_1094),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1171),
.B(n_1174),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1082),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_1127),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_SL g1227 ( 
.A(n_1091),
.B(n_1100),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1167),
.A2(n_1187),
.B(n_1172),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1127),
.Y(n_1229)
);

INVx1_ASAP7_75t_SL g1230 ( 
.A(n_1156),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1177),
.B(n_1182),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1192),
.A2(n_1201),
.B(n_1063),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1183),
.B(n_1188),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1170),
.Y(n_1234)
);

AOI21xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1078),
.A2(n_1195),
.B(n_1147),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1183),
.B(n_1188),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1175),
.B(n_1093),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1086),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1124),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1106),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1105),
.A2(n_1061),
.B(n_1102),
.Y(n_1241)
);

BUFx12f_ASAP7_75t_L g1242 ( 
.A(n_1094),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1067),
.A2(n_1083),
.B(n_1089),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1179),
.A2(n_1158),
.B1(n_1067),
.B2(n_1057),
.Y(n_1244)
);

AOI222xp33_ASAP7_75t_L g1245 ( 
.A1(n_1154),
.A2(n_1179),
.B1(n_1062),
.B2(n_1185),
.C1(n_1169),
.C2(n_1064),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_1071),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1048),
.B(n_1143),
.Y(n_1247)
);

BUFx10_ASAP7_75t_L g1248 ( 
.A(n_1107),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1125),
.Y(n_1249)
);

INVx4_ASAP7_75t_L g1250 ( 
.A(n_1170),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1062),
.A2(n_1155),
.B1(n_1092),
.B2(n_1090),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1106),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1205),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1066),
.A2(n_1196),
.B(n_1159),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1097),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1073),
.B(n_1142),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1149),
.B(n_1165),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1173),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1097),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1129),
.B(n_1098),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1135),
.B(n_1136),
.Y(n_1261)
);

NOR2xp67_ASAP7_75t_L g1262 ( 
.A(n_1138),
.B(n_1107),
.Y(n_1262)
);

AND2x2_ASAP7_75t_SL g1263 ( 
.A(n_1058),
.B(n_1092),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_1120),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1118),
.A2(n_1112),
.B1(n_1111),
.B2(n_1103),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1085),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1156),
.B(n_1104),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1126),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1159),
.A2(n_1196),
.B(n_1176),
.Y(n_1269)
);

OR2x6_ASAP7_75t_L g1270 ( 
.A(n_1087),
.B(n_1173),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1152),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1121),
.Y(n_1272)
);

OR2x6_ASAP7_75t_L g1273 ( 
.A(n_1087),
.B(n_1068),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1081),
.B(n_1072),
.Y(n_1274)
);

OAI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1070),
.A2(n_1111),
.B1(n_1103),
.B2(n_1072),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1132),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1199),
.B(n_1087),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1202),
.B(n_1199),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1176),
.A2(n_1055),
.B(n_1059),
.Y(n_1279)
);

NAND2xp33_ASAP7_75t_L g1280 ( 
.A(n_1115),
.B(n_1055),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1132),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1097),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1059),
.A2(n_1108),
.B(n_1084),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1068),
.B(n_1128),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1202),
.A2(n_1074),
.B1(n_1114),
.B2(n_1056),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1109),
.B(n_1203),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1191),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1191),
.B(n_1203),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1123),
.B(n_1056),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1096),
.A2(n_1110),
.B(n_1074),
.C(n_1134),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1130),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1133),
.A2(n_1119),
.B1(n_1131),
.B2(n_1122),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1095),
.A2(n_1065),
.B(n_1053),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1084),
.A2(n_1133),
.B1(n_1190),
.B2(n_1099),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1056),
.B(n_1113),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1116),
.B(n_1117),
.Y(n_1296)
);

BUFx10_ASAP7_75t_L g1297 ( 
.A(n_1099),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1052),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1099),
.B(n_1198),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1139),
.B(n_1198),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1101),
.A2(n_1060),
.B(n_1050),
.Y(n_1301)
);

BUFx12f_ASAP7_75t_L g1302 ( 
.A(n_1139),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1140),
.A2(n_1178),
.B(n_1197),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1079),
.Y(n_1304)
);

BUFx10_ASAP7_75t_L g1305 ( 
.A(n_1139),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1186),
.B(n_1198),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1186),
.B(n_1075),
.Y(n_1307)
);

OR2x2_ASAP7_75t_SL g1308 ( 
.A(n_1186),
.B(n_1075),
.Y(n_1308)
);

NAND2x1p5_ASAP7_75t_L g1309 ( 
.A(n_1076),
.B(n_1184),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1148),
.A2(n_1150),
.B1(n_1163),
.B2(n_1189),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1194),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1200),
.B(n_1054),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1054),
.B(n_1151),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_SL g1314 ( 
.A1(n_1159),
.A2(n_1196),
.B(n_1176),
.C(n_1155),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1157),
.A2(n_1164),
.B(n_1193),
.C(n_1049),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1049),
.B(n_1157),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1120),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1080),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1088),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1049),
.A2(n_1164),
.B(n_1157),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1054),
.B(n_1151),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1048),
.B(n_1143),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1054),
.B(n_1151),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1080),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1145),
.A2(n_699),
.B1(n_1033),
.B2(n_689),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1077),
.B(n_1141),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1054),
.B(n_1151),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1095),
.A2(n_1065),
.B(n_1053),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1088),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1088),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1125),
.Y(n_1331)
);

BUFx12f_ASAP7_75t_L g1332 ( 
.A(n_1094),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1048),
.B(n_1143),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1127),
.Y(n_1334)
);

AOI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1096),
.A2(n_1137),
.B(n_1051),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1157),
.A2(n_1193),
.B(n_1164),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1127),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1125),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1048),
.B(n_1143),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1071),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1157),
.A2(n_1193),
.B(n_1164),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1125),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1054),
.B(n_1151),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1171),
.B(n_1174),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1125),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1088),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1127),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1125),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1080),
.Y(n_1349)
);

O2A1O1Ixp5_ASAP7_75t_L g1350 ( 
.A1(n_1145),
.A2(n_1204),
.B(n_1049),
.C(n_1164),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1054),
.B(n_1151),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1054),
.B(n_1151),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1127),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1077),
.B(n_1141),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1054),
.B(n_1151),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1125),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1106),
.Y(n_1357)
);

OAI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1227),
.A2(n_1344),
.B1(n_1244),
.B2(n_1327),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1247),
.Y(n_1359)
);

INVx5_ASAP7_75t_L g1360 ( 
.A(n_1273),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1209),
.A2(n_1207),
.B1(n_1344),
.B2(n_1320),
.Y(n_1361)
);

INVxp33_ASAP7_75t_L g1362 ( 
.A(n_1213),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1215),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1222),
.B(n_1263),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1225),
.Y(n_1365)
);

BUFx2_ASAP7_75t_R g1366 ( 
.A(n_1331),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1224),
.A2(n_1245),
.B1(n_1263),
.B2(n_1222),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1289),
.B(n_1210),
.Y(n_1368)
);

BUFx2_ASAP7_75t_R g1369 ( 
.A(n_1331),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1325),
.A2(n_1244),
.B1(n_1237),
.B2(n_1251),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1216),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1238),
.Y(n_1372)
);

AO21x1_ASAP7_75t_SL g1373 ( 
.A1(n_1241),
.A2(n_1240),
.B(n_1216),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1217),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1302),
.A2(n_1325),
.B1(n_1336),
.B2(n_1341),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1232),
.A2(n_1228),
.B(n_1214),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1266),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1316),
.A2(n_1326),
.B1(n_1220),
.B2(n_1354),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1260),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1271),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1351),
.A2(n_1206),
.B1(n_1329),
.B2(n_1330),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1253),
.A2(n_1346),
.B1(n_1355),
.B2(n_1352),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1308),
.Y(n_1383)
);

AO21x1_ASAP7_75t_L g1384 ( 
.A1(n_1315),
.A2(n_1211),
.B(n_1208),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1232),
.A2(n_1228),
.B(n_1214),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1217),
.Y(n_1386)
);

BUFx12f_ASAP7_75t_L g1387 ( 
.A(n_1223),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1218),
.B(n_1221),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1240),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1252),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1267),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1306),
.B(n_1276),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1252),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1231),
.B(n_1233),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1315),
.A2(n_1321),
.B1(n_1236),
.B2(n_1343),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1318),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1350),
.A2(n_1211),
.B(n_1208),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1324),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1261),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1349),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1281),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1230),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1219),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1300),
.B(n_1295),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1357),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1313),
.A2(n_1323),
.B1(n_1319),
.B2(n_1219),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1285),
.A2(n_1278),
.B1(n_1317),
.B2(n_1265),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1256),
.A2(n_1257),
.B1(n_1307),
.B2(n_1274),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1303),
.A2(n_1293),
.B(n_1328),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1287),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1235),
.A2(n_1285),
.B(n_1279),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1303),
.A2(n_1243),
.B(n_1335),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1299),
.B(n_1357),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1297),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1243),
.A2(n_1290),
.B(n_1301),
.Y(n_1415)
);

INVxp67_ASAP7_75t_SL g1416 ( 
.A(n_1312),
.Y(n_1416)
);

OAI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1273),
.A2(n_1272),
.B1(n_1264),
.B2(n_1270),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1280),
.A2(n_1268),
.B1(n_1239),
.B2(n_1277),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1340),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1286),
.Y(n_1420)
);

AO21x1_ASAP7_75t_L g1421 ( 
.A1(n_1275),
.A2(n_1294),
.B(n_1254),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1288),
.Y(n_1422)
);

BUFx8_ASAP7_75t_SL g1423 ( 
.A(n_1242),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1269),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1255),
.Y(n_1425)
);

INVxp67_ASAP7_75t_SL g1426 ( 
.A(n_1269),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1255),
.Y(n_1427)
);

AOI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1254),
.A2(n_1283),
.B(n_1311),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1259),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1322),
.B(n_1333),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1246),
.A2(n_1262),
.B1(n_1339),
.B2(n_1333),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1350),
.A2(n_1314),
.B(n_1279),
.Y(n_1432)
);

OR2x6_ASAP7_75t_L g1433 ( 
.A(n_1270),
.B(n_1322),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1339),
.B(n_1277),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1259),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1298),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1283),
.B(n_1305),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_SL g1438 ( 
.A(n_1338),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1305),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1217),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1284),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1248),
.Y(n_1442)
);

BUFx2_ASAP7_75t_SL g1443 ( 
.A(n_1217),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1234),
.B(n_1258),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1270),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1234),
.A2(n_1246),
.B1(n_1337),
.B2(n_1248),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1304),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1234),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1234),
.A2(n_1258),
.B1(n_1250),
.B2(n_1348),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1304),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1290),
.A2(n_1249),
.B(n_1314),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1304),
.Y(n_1452)
);

AO21x1_ASAP7_75t_L g1453 ( 
.A1(n_1292),
.A2(n_1296),
.B(n_1309),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1282),
.B(n_1353),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1309),
.A2(n_1296),
.B(n_1291),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1226),
.B(n_1229),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1310),
.A2(n_1304),
.B(n_1291),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1212),
.A2(n_1226),
.B(n_1229),
.Y(n_1458)
);

NAND2x1p5_ASAP7_75t_L g1459 ( 
.A(n_1337),
.B(n_1353),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1334),
.Y(n_1460)
);

AOI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1334),
.A2(n_1347),
.B(n_1250),
.Y(n_1461)
);

INVx8_ASAP7_75t_L g1462 ( 
.A(n_1332),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1347),
.B(n_1338),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1342),
.A2(n_1345),
.B1(n_1348),
.B2(n_1356),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1342),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1345),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1356),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1215),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1344),
.A2(n_699),
.B1(n_1033),
.B2(n_1325),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1215),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1215),
.Y(n_1471)
);

BUFx4f_ASAP7_75t_SL g1472 ( 
.A(n_1223),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1297),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1266),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1215),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1232),
.A2(n_1228),
.B(n_1214),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1215),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1344),
.A2(n_1227),
.B1(n_582),
.B2(n_1100),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1216),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1210),
.B(n_1327),
.Y(n_1480)
);

BUFx2_ASAP7_75t_R g1481 ( 
.A(n_1331),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1216),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1273),
.B(n_1247),
.Y(n_1483)
);

OR2x6_ASAP7_75t_L g1484 ( 
.A(n_1302),
.B(n_1067),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1374),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1397),
.A2(n_1432),
.B(n_1421),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1374),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1404),
.B(n_1405),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1383),
.B(n_1413),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1412),
.A2(n_1409),
.B(n_1428),
.Y(n_1490)
);

BUFx2_ASAP7_75t_R g1491 ( 
.A(n_1423),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1363),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1412),
.A2(n_1409),
.B(n_1421),
.Y(n_1493)
);

AO21x1_ASAP7_75t_SL g1494 ( 
.A1(n_1367),
.A2(n_1370),
.B(n_1371),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1360),
.B(n_1414),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1480),
.B(n_1388),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1404),
.B(n_1405),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1368),
.B(n_1392),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1410),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1394),
.B(n_1395),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1383),
.B(n_1413),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1361),
.B(n_1368),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1392),
.B(n_1437),
.Y(n_1503)
);

CKINVDCx11_ASAP7_75t_R g1504 ( 
.A(n_1387),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1479),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1371),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1389),
.Y(n_1507)
);

AO21x2_ASAP7_75t_L g1508 ( 
.A1(n_1453),
.A2(n_1384),
.B(n_1407),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1389),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1390),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1390),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1437),
.B(n_1424),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1393),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1393),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1420),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1426),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1469),
.A2(n_1358),
.B1(n_1484),
.B2(n_1375),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1456),
.Y(n_1518)
);

AO21x2_ASAP7_75t_L g1519 ( 
.A1(n_1453),
.A2(n_1384),
.B(n_1428),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_SL g1520 ( 
.A(n_1366),
.B(n_1369),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1416),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1479),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1450),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1484),
.B(n_1414),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1399),
.B(n_1379),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1401),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1365),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1372),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1396),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1377),
.Y(n_1530)
);

BUFx8_ASAP7_75t_L g1531 ( 
.A(n_1387),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1398),
.Y(n_1532)
);

CKINVDCx11_ASAP7_75t_R g1533 ( 
.A(n_1462),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1474),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1482),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1400),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1482),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1411),
.A2(n_1451),
.B(n_1455),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1478),
.B(n_1419),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1468),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1456),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1450),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1373),
.B(n_1470),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1471),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1380),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1450),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1481),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1475),
.B(n_1477),
.Y(n_1548)
);

INVxp67_ASAP7_75t_L g1549 ( 
.A(n_1402),
.Y(n_1549)
);

NOR2xp67_ASAP7_75t_SL g1550 ( 
.A(n_1443),
.B(n_1374),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1364),
.B(n_1362),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1364),
.B(n_1362),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1391),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1460),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1422),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1466),
.B(n_1463),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1403),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1408),
.B(n_1418),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1415),
.B(n_1378),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1439),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1406),
.B(n_1382),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1439),
.Y(n_1562)
);

AOI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1461),
.A2(n_1376),
.B(n_1385),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1441),
.Y(n_1564)
);

OR2x6_ASAP7_75t_L g1565 ( 
.A(n_1433),
.B(n_1473),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1460),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1436),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1447),
.A2(n_1452),
.B(n_1435),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1436),
.Y(n_1569)
);

AO21x2_ASAP7_75t_L g1570 ( 
.A1(n_1445),
.A2(n_1427),
.B(n_1425),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1467),
.B(n_1472),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1429),
.Y(n_1572)
);

INVxp33_ASAP7_75t_L g1573 ( 
.A(n_1438),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1381),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1448),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1414),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1465),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1423),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1476),
.A2(n_1473),
.B(n_1457),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1563),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1503),
.B(n_1415),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1563),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1503),
.B(n_1457),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1512),
.B(n_1457),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1505),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1505),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1522),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1488),
.B(n_1467),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1559),
.B(n_1454),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1559),
.B(n_1454),
.Y(n_1590)
);

AO31x2_ASAP7_75t_L g1591 ( 
.A1(n_1516),
.A2(n_1434),
.A3(n_1444),
.B(n_1430),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1498),
.B(n_1440),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1579),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1498),
.B(n_1440),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1486),
.B(n_1440),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1486),
.B(n_1519),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1570),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1522),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1533),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1535),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1504),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1488),
.B(n_1386),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1497),
.B(n_1386),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1486),
.B(n_1543),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1500),
.B(n_1374),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1497),
.B(n_1502),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1524),
.B(n_1360),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1539),
.B(n_1526),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1493),
.B(n_1538),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1535),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1493),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1538),
.B(n_1359),
.Y(n_1612)
);

OAI33xp33_ASAP7_75t_L g1613 ( 
.A1(n_1558),
.A2(n_1417),
.A3(n_1464),
.B1(n_1462),
.B2(n_1431),
.B3(n_1458),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1549),
.B(n_1442),
.Y(n_1614)
);

INVx4_ASAP7_75t_L g1615 ( 
.A(n_1538),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1521),
.B(n_1443),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1538),
.B(n_1359),
.Y(n_1617)
);

AND2x4_ASAP7_75t_SL g1618 ( 
.A(n_1565),
.B(n_1433),
.Y(n_1618)
);

NAND3xp33_ASAP7_75t_L g1619 ( 
.A(n_1517),
.B(n_1446),
.C(n_1449),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1490),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1548),
.B(n_1567),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1568),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_SL g1623 ( 
.A1(n_1547),
.A2(n_1433),
.B1(n_1360),
.B2(n_1483),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1537),
.B(n_1459),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1521),
.B(n_1553),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1581),
.B(n_1569),
.Y(n_1626)
);

AND2x2_ASAP7_75t_SL g1627 ( 
.A(n_1618),
.B(n_1524),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1606),
.B(n_1545),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_SL g1629 ( 
.A1(n_1609),
.A2(n_1571),
.B(n_1573),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1606),
.B(n_1530),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1606),
.B(n_1534),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1622),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1581),
.B(n_1542),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1608),
.B(n_1605),
.Y(n_1634)
);

NAND3xp33_ASAP7_75t_L g1635 ( 
.A(n_1596),
.B(n_1555),
.C(n_1577),
.Y(n_1635)
);

AOI211xp5_ASAP7_75t_L g1636 ( 
.A1(n_1609),
.A2(n_1556),
.B(n_1520),
.C(n_1572),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1619),
.A2(n_1525),
.B1(n_1515),
.B2(n_1499),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1589),
.B(n_1542),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1592),
.B(n_1499),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_L g1640 ( 
.A(n_1596),
.B(n_1510),
.C(n_1507),
.Y(n_1640)
);

NOR3xp33_ASAP7_75t_L g1641 ( 
.A(n_1615),
.B(n_1576),
.C(n_1575),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1608),
.B(n_1496),
.Y(n_1642)
);

OAI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1619),
.A2(n_1564),
.B1(n_1561),
.B2(n_1527),
.C(n_1529),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1589),
.B(n_1489),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1612),
.A2(n_1508),
.B(n_1617),
.Y(n_1645)
);

NAND4xp25_ASAP7_75t_L g1646 ( 
.A(n_1614),
.B(n_1576),
.C(n_1544),
.D(n_1540),
.Y(n_1646)
);

AND2x2_ASAP7_75t_SL g1647 ( 
.A(n_1618),
.B(n_1489),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1589),
.B(n_1489),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1621),
.B(n_1492),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1580),
.A2(n_1582),
.B(n_1620),
.Y(n_1650)
);

NAND2xp33_ASAP7_75t_SL g1651 ( 
.A(n_1599),
.B(n_1578),
.Y(n_1651)
);

OAI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1619),
.A2(n_1528),
.B1(n_1532),
.B2(n_1536),
.C(n_1560),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_SL g1653 ( 
.A1(n_1609),
.A2(n_1491),
.B(n_1551),
.Y(n_1653)
);

NAND2xp33_ASAP7_75t_L g1654 ( 
.A(n_1599),
.B(n_1578),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1621),
.B(n_1506),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_L g1656 ( 
.A(n_1596),
.B(n_1509),
.C(n_1514),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1589),
.B(n_1501),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1613),
.A2(n_1494),
.B1(n_1574),
.B2(n_1508),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1621),
.B(n_1506),
.Y(n_1659)
);

OA21x2_ASAP7_75t_L g1660 ( 
.A1(n_1597),
.A2(n_1560),
.B(n_1562),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1625),
.B(n_1507),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_L g1662 ( 
.A(n_1596),
.B(n_1511),
.C(n_1514),
.Y(n_1662)
);

AO221x1_ASAP7_75t_L g1663 ( 
.A1(n_1586),
.A2(n_1487),
.B1(n_1485),
.B2(n_1546),
.C(n_1523),
.Y(n_1663)
);

NAND3xp33_ASAP7_75t_L g1664 ( 
.A(n_1609),
.B(n_1509),
.C(n_1510),
.Y(n_1664)
);

OAI221xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1604),
.A2(n_1552),
.B1(n_1551),
.B2(n_1513),
.C(n_1511),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1625),
.B(n_1513),
.Y(n_1666)
);

NAND3xp33_ASAP7_75t_L g1667 ( 
.A(n_1615),
.B(n_1562),
.C(n_1566),
.Y(n_1667)
);

OAI21xp5_ASAP7_75t_SL g1668 ( 
.A1(n_1604),
.A2(n_1617),
.B(n_1612),
.Y(n_1668)
);

OAI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1615),
.A2(n_1557),
.B1(n_1554),
.B2(n_1442),
.C(n_1552),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1590),
.B(n_1508),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1590),
.B(n_1554),
.Y(n_1671)
);

NOR3xp33_ASAP7_75t_L g1672 ( 
.A(n_1615),
.B(n_1613),
.C(n_1611),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1590),
.B(n_1570),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1590),
.B(n_1501),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1612),
.B(n_1485),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1604),
.A2(n_1531),
.B(n_1501),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1588),
.B(n_1570),
.Y(n_1677)
);

NAND4xp25_ASAP7_75t_L g1678 ( 
.A(n_1614),
.B(n_1523),
.C(n_1546),
.D(n_1518),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1588),
.B(n_1541),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1617),
.A2(n_1531),
.B(n_1495),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1615),
.A2(n_1607),
.B(n_1595),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1628),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1663),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1675),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1660),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1660),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1644),
.B(n_1583),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1644),
.B(n_1583),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1677),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1660),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1648),
.B(n_1657),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1664),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1670),
.B(n_1587),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1634),
.B(n_1588),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1648),
.B(n_1583),
.Y(n_1695)
);

AND2x2_ASAP7_75t_SL g1696 ( 
.A(n_1627),
.B(n_1615),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1650),
.B(n_1593),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1673),
.B(n_1587),
.Y(n_1698)
);

INVx3_ASAP7_75t_L g1699 ( 
.A(n_1650),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1626),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1661),
.B(n_1598),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1626),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1640),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1656),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1632),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1666),
.B(n_1598),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1662),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1642),
.B(n_1600),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1633),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1633),
.Y(n_1710)
);

AND2x4_ASAP7_75t_SL g1711 ( 
.A(n_1657),
.B(n_1595),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1674),
.B(n_1593),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1636),
.B(n_1586),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1638),
.B(n_1584),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1678),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1655),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1638),
.B(n_1584),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1672),
.B(n_1600),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1668),
.B(n_1592),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1667),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1659),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1675),
.B(n_1592),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1671),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1649),
.Y(n_1724)
);

AND2x4_ASAP7_75t_SL g1725 ( 
.A(n_1639),
.B(n_1595),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1635),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1682),
.B(n_1637),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1692),
.B(n_1630),
.Y(n_1728)
);

OR2x6_ASAP7_75t_L g1729 ( 
.A(n_1720),
.B(n_1645),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1703),
.B(n_1601),
.Y(n_1730)
);

OAI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1726),
.A2(n_1643),
.B1(n_1629),
.B2(n_1658),
.C(n_1652),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1711),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1708),
.Y(n_1733)
);

NOR2xp67_ASAP7_75t_SL g1734 ( 
.A(n_1713),
.B(n_1601),
.Y(n_1734)
);

OAI211xp5_ASAP7_75t_L g1735 ( 
.A1(n_1703),
.A2(n_1646),
.B(n_1681),
.C(n_1651),
.Y(n_1735)
);

NOR2xp67_ASAP7_75t_L g1736 ( 
.A(n_1683),
.B(n_1653),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1718),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1682),
.B(n_1631),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1704),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1708),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1719),
.B(n_1592),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1690),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1719),
.B(n_1594),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1719),
.B(n_1594),
.Y(n_1744)
);

NOR3xp33_ASAP7_75t_L g1745 ( 
.A(n_1726),
.B(n_1669),
.C(n_1665),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1694),
.B(n_1586),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1724),
.Y(n_1747)
);

NAND2x1p5_ASAP7_75t_L g1748 ( 
.A(n_1696),
.B(n_1647),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1690),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1694),
.B(n_1591),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1707),
.B(n_1591),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1701),
.B(n_1602),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1718),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1700),
.B(n_1594),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1692),
.B(n_1610),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1700),
.B(n_1594),
.Y(n_1756)
);

OR2x6_ASAP7_75t_L g1757 ( 
.A(n_1720),
.B(n_1623),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1701),
.B(n_1602),
.Y(n_1758)
);

NOR2x1p5_ASAP7_75t_L g1759 ( 
.A(n_1726),
.B(n_1651),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1707),
.B(n_1591),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1700),
.B(n_1585),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1724),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1724),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1704),
.A2(n_1641),
.B(n_1654),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1692),
.B(n_1654),
.Y(n_1765)
);

INVx2_ASAP7_75t_SL g1766 ( 
.A(n_1711),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1706),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1728),
.B(n_1707),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1739),
.B(n_1720),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1728),
.B(n_1693),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1747),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1745),
.B(n_1720),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1762),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1732),
.B(n_1715),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1742),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1764),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1763),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1737),
.B(n_1716),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1751),
.B(n_1760),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1730),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1742),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1755),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1730),
.B(n_1531),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1755),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1767),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1749),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1732),
.B(n_1715),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1766),
.B(n_1741),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1753),
.B(n_1716),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1733),
.B(n_1693),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1766),
.B(n_1715),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1749),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1752),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1758),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1741),
.B(n_1702),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1765),
.B(n_1462),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1743),
.B(n_1702),
.Y(n_1797)
);

INVx2_ASAP7_75t_SL g1798 ( 
.A(n_1759),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1740),
.Y(n_1799)
);

AND2x2_ASAP7_75t_SL g1800 ( 
.A(n_1765),
.B(n_1696),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1738),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1734),
.B(n_1462),
.Y(n_1802)
);

OAI221xp5_ASAP7_75t_SL g1803 ( 
.A1(n_1729),
.A2(n_1686),
.B1(n_1685),
.B2(n_1690),
.C(n_1683),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1743),
.B(n_1702),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1754),
.Y(n_1805)
);

NOR2x1_ASAP7_75t_L g1806 ( 
.A(n_1735),
.B(n_1713),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1750),
.B(n_1727),
.Y(n_1807)
);

AND2x2_ASAP7_75t_SL g1808 ( 
.A(n_1761),
.B(n_1696),
.Y(n_1808)
);

INVx2_ASAP7_75t_SL g1809 ( 
.A(n_1761),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1754),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1771),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1771),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1782),
.Y(n_1813)
);

OR2x6_ASAP7_75t_L g1814 ( 
.A(n_1772),
.B(n_1729),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1773),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1773),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1800),
.B(n_1744),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1768),
.B(n_1698),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1800),
.B(n_1744),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1768),
.B(n_1698),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1776),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1780),
.B(n_1783),
.Y(n_1822)
);

CKINVDCx16_ASAP7_75t_R g1823 ( 
.A(n_1802),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1798),
.B(n_1729),
.Y(n_1824)
);

INVxp67_ASAP7_75t_L g1825 ( 
.A(n_1776),
.Y(n_1825)
);

INVxp67_ASAP7_75t_L g1826 ( 
.A(n_1796),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1775),
.Y(n_1827)
);

CKINVDCx16_ASAP7_75t_R g1828 ( 
.A(n_1806),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1777),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1782),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1808),
.B(n_1756),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1777),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1775),
.Y(n_1833)
);

AO21x2_ASAP7_75t_L g1834 ( 
.A1(n_1769),
.A2(n_1731),
.B(n_1686),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1803),
.A2(n_1729),
.B(n_1757),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1798),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1808),
.B(n_1795),
.Y(n_1837)
);

INVx1_ASAP7_75t_SL g1838 ( 
.A(n_1774),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1795),
.B(n_1756),
.Y(n_1839)
);

INVx1_ASAP7_75t_SL g1840 ( 
.A(n_1774),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1797),
.B(n_1748),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1770),
.B(n_1706),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1801),
.B(n_1746),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1781),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1807),
.A2(n_1736),
.B1(n_1748),
.B2(n_1757),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1784),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1837),
.B(n_1787),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1811),
.Y(n_1848)
);

AOI31xp33_ASAP7_75t_L g1849 ( 
.A1(n_1825),
.A2(n_1791),
.A3(n_1787),
.B(n_1809),
.Y(n_1849)
);

AOI21xp33_ASAP7_75t_SL g1850 ( 
.A1(n_1828),
.A2(n_1809),
.B(n_1791),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1834),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1839),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1834),
.A2(n_1757),
.B1(n_1807),
.B2(n_1801),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1834),
.A2(n_1757),
.B1(n_1793),
.B2(n_1794),
.Y(n_1854)
);

AOI322xp5_ASAP7_75t_L g1855 ( 
.A1(n_1821),
.A2(n_1685),
.A3(n_1686),
.B1(n_1690),
.B2(n_1784),
.C1(n_1786),
.C2(n_1792),
.Y(n_1855)
);

AOI221xp5_ASAP7_75t_L g1856 ( 
.A1(n_1835),
.A2(n_1779),
.B1(n_1786),
.B2(n_1685),
.C(n_1799),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1811),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1843),
.B(n_1838),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1812),
.Y(n_1859)
);

AOI21xp33_ASAP7_75t_L g1860 ( 
.A1(n_1814),
.A2(n_1846),
.B(n_1830),
.Y(n_1860)
);

NOR2xp67_ASAP7_75t_L g1861 ( 
.A(n_1845),
.B(n_1793),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1840),
.B(n_1794),
.Y(n_1862)
);

INVxp67_ASAP7_75t_SL g1863 ( 
.A(n_1836),
.Y(n_1863)
);

O2A1O1Ixp5_ASAP7_75t_L g1864 ( 
.A1(n_1846),
.A2(n_1785),
.B(n_1799),
.C(n_1778),
.Y(n_1864)
);

A2O1A1Ixp33_ASAP7_75t_L g1865 ( 
.A1(n_1837),
.A2(n_1831),
.B(n_1822),
.C(n_1819),
.Y(n_1865)
);

AOI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1814),
.A2(n_1824),
.B(n_1813),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1839),
.B(n_1785),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1827),
.Y(n_1868)
);

OAI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1814),
.A2(n_1789),
.B(n_1797),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1812),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1815),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1817),
.B(n_1819),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1831),
.A2(n_1683),
.B1(n_1804),
.B2(n_1805),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1848),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1863),
.B(n_1826),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1857),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1863),
.B(n_1817),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1859),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1864),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1852),
.B(n_1847),
.Y(n_1880)
);

INVx1_ASAP7_75t_SL g1881 ( 
.A(n_1858),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1854),
.A2(n_1814),
.B1(n_1824),
.B2(n_1823),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_1872),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1865),
.B(n_1841),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1865),
.B(n_1841),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1862),
.B(n_1804),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1867),
.B(n_1818),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1866),
.B(n_1818),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1861),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1849),
.B(n_1820),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1850),
.B(n_1820),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1869),
.B(n_1788),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1864),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1851),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_SL g1895 ( 
.A1(n_1879),
.A2(n_1824),
.B(n_1851),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1879),
.A2(n_1860),
.B(n_1853),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1883),
.B(n_1870),
.Y(n_1897)
);

OAI211xp5_ASAP7_75t_L g1898 ( 
.A1(n_1893),
.A2(n_1855),
.B(n_1856),
.C(n_1871),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1893),
.A2(n_1873),
.B(n_1816),
.Y(n_1899)
);

OAI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1889),
.A2(n_1779),
.B1(n_1868),
.B2(n_1770),
.Y(n_1900)
);

NAND3xp33_ASAP7_75t_L g1901 ( 
.A(n_1884),
.B(n_1868),
.C(n_1816),
.Y(n_1901)
);

NOR3xp33_ASAP7_75t_L g1902 ( 
.A(n_1875),
.B(n_1829),
.C(n_1815),
.Y(n_1902)
);

NAND3xp33_ASAP7_75t_L g1903 ( 
.A(n_1884),
.B(n_1832),
.C(n_1829),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1890),
.A2(n_1842),
.B1(n_1805),
.B2(n_1810),
.Y(n_1904)
);

OAI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1881),
.A2(n_1842),
.B1(n_1810),
.B2(n_1790),
.Y(n_1905)
);

NAND3xp33_ASAP7_75t_L g1906 ( 
.A(n_1885),
.B(n_1877),
.C(n_1882),
.Y(n_1906)
);

AOI222xp33_ASAP7_75t_L g1907 ( 
.A1(n_1885),
.A2(n_1844),
.B1(n_1833),
.B2(n_1827),
.C1(n_1832),
.C2(n_1792),
.Y(n_1907)
);

A2O1A1Ixp33_ASAP7_75t_L g1908 ( 
.A1(n_1888),
.A2(n_1891),
.B(n_1892),
.C(n_1887),
.Y(n_1908)
);

NAND3xp33_ASAP7_75t_SL g1909 ( 
.A(n_1898),
.B(n_1892),
.C(n_1886),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1908),
.B(n_1880),
.Y(n_1910)
);

NOR4xp25_ASAP7_75t_SL g1911 ( 
.A(n_1895),
.B(n_1874),
.C(n_1878),
.D(n_1876),
.Y(n_1911)
);

NAND4xp75_ASAP7_75t_L g1912 ( 
.A(n_1896),
.B(n_1894),
.C(n_1844),
.D(n_1833),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1900),
.B(n_1880),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1901),
.Y(n_1914)
);

NAND4xp25_ASAP7_75t_L g1915 ( 
.A(n_1899),
.B(n_1880),
.C(n_1894),
.D(n_1788),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1907),
.B(n_1790),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1906),
.B(n_1781),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1905),
.B(n_1696),
.Y(n_1918)
);

NOR3xp33_ASAP7_75t_L g1919 ( 
.A(n_1897),
.B(n_1699),
.C(n_1689),
.Y(n_1919)
);

OAI221xp5_ASAP7_75t_L g1920 ( 
.A1(n_1914),
.A2(n_1903),
.B1(n_1902),
.B2(n_1904),
.C(n_1699),
.Y(n_1920)
);

O2A1O1Ixp5_ASAP7_75t_L g1921 ( 
.A1(n_1913),
.A2(n_1699),
.B(n_1697),
.C(n_1723),
.Y(n_1921)
);

NAND4xp25_ASAP7_75t_L g1922 ( 
.A(n_1909),
.B(n_1699),
.C(n_1680),
.D(n_1697),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1911),
.A2(n_1699),
.B(n_1684),
.Y(n_1923)
);

INVxp67_ASAP7_75t_L g1924 ( 
.A(n_1910),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1916),
.B(n_1684),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1924),
.A2(n_1912),
.B1(n_1917),
.B2(n_1915),
.Y(n_1926)
);

AOI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1925),
.A2(n_1918),
.B1(n_1919),
.B2(n_1684),
.Y(n_1927)
);

OAI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1920),
.A2(n_1723),
.B1(n_1721),
.B2(n_1716),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1921),
.Y(n_1929)
);

NOR2x1_ASAP7_75t_L g1930 ( 
.A(n_1922),
.B(n_1697),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1923),
.A2(n_1697),
.B1(n_1689),
.B2(n_1711),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1924),
.B(n_1691),
.Y(n_1932)
);

NOR4xp25_ASAP7_75t_L g1933 ( 
.A(n_1929),
.B(n_1721),
.C(n_1723),
.D(n_1717),
.Y(n_1933)
);

OAI221xp5_ASAP7_75t_L g1934 ( 
.A1(n_1926),
.A2(n_1676),
.B1(n_1705),
.B2(n_1723),
.C(n_1597),
.Y(n_1934)
);

NOR2x1_ASAP7_75t_L g1935 ( 
.A(n_1932),
.B(n_1697),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1927),
.B(n_1721),
.Y(n_1936)
);

NOR3x2_ASAP7_75t_L g1937 ( 
.A(n_1928),
.B(n_1624),
.C(n_1603),
.Y(n_1937)
);

NOR4xp75_ASAP7_75t_SL g1938 ( 
.A(n_1931),
.B(n_1679),
.C(n_1616),
.D(n_1697),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1936),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1933),
.B(n_1930),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1935),
.B(n_1691),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1940),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1942),
.B(n_1940),
.Y(n_1943)
);

AOI221x1_ASAP7_75t_L g1944 ( 
.A1(n_1943),
.A2(n_1939),
.B1(n_1941),
.B2(n_1938),
.C(n_1934),
.Y(n_1944)
);

BUFx2_ASAP7_75t_L g1945 ( 
.A(n_1943),
.Y(n_1945)
);

OAI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1945),
.A2(n_1937),
.B1(n_1709),
.B2(n_1710),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1944),
.A2(n_1688),
.B(n_1687),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1947),
.A2(n_1946),
.B1(n_1688),
.B2(n_1695),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1947),
.A2(n_1688),
.B(n_1687),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1948),
.B(n_1705),
.Y(n_1950)
);

OAI211xp5_ASAP7_75t_L g1951 ( 
.A1(n_1950),
.A2(n_1949),
.B(n_1722),
.C(n_1717),
.Y(n_1951)
);

OAI221xp5_ASAP7_75t_R g1952 ( 
.A1(n_1951),
.A2(n_1717),
.B1(n_1714),
.B2(n_1712),
.C(n_1725),
.Y(n_1952)
);

AOI211xp5_ASAP7_75t_L g1953 ( 
.A1(n_1952),
.A2(n_1550),
.B(n_1623),
.C(n_1487),
.Y(n_1953)
);


endmodule