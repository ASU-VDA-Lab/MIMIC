module fake_jpeg_19016_n_144 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_16),
.B(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_77),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_72),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_50),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_1),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_58),
.B(n_60),
.C(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_66),
.Y(n_105)
);

INVx5_ASAP7_75t_SL g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_47),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_53),
.B1(n_70),
.B2(n_56),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_53),
.B1(n_70),
.B2(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_90),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_95),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_101),
.B1(n_54),
.B2(n_49),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_99),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_71),
.B1(n_51),
.B2(n_55),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_65),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_104),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_105),
.B(n_3),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_104),
.A2(n_63),
.B(n_57),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_117),
.B(n_4),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_116),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_67),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_119),
.C(n_13),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_19),
.Y(n_123)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_14),
.B(n_15),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_25),
.C(n_46),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_123),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_5),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_124),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_6),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_126),
.C(n_127),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_112),
.C(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_134),
.C(n_114),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_114),
.B(n_131),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_130),
.C(n_132),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_135),
.B1(n_32),
.B2(n_34),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_128),
.C(n_37),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_108),
.C(n_42),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_29),
.B(n_43),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_44),
.Y(n_144)
);


endmodule