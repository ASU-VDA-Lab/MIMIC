module fake_jpeg_3074_n_520 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_520);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_520;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_10),
.B(n_12),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_51),
.Y(n_157)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_54),
.Y(n_143)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_67),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_69),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_78),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_34),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_23),
.B(n_15),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_85),
.Y(n_131)
);

BUFx4f_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_15),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

BUFx16f_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_22),
.B(n_35),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_89),
.B(n_90),
.Y(n_154)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_47),
.B(n_16),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_94),
.Y(n_134)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_39),
.Y(n_132)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_14),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_21),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_97),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_28),
.B(n_14),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_99),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_48),
.B1(n_19),
.B2(n_28),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_107),
.A2(n_113),
.B1(n_117),
.B2(n_118),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_33),
.B1(n_46),
.B2(n_19),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_84),
.A2(n_33),
.B1(n_48),
.B2(n_36),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_55),
.A2(n_48),
.B1(n_40),
.B2(n_36),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_123),
.B(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_53),
.B(n_21),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_124),
.B(n_158),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_89),
.A2(n_36),
.B1(n_40),
.B2(n_32),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_127),
.A2(n_137),
.B1(n_93),
.B2(n_99),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_132),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_40),
.C(n_36),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_60),
.C(n_90),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_58),
.A2(n_40),
.B1(n_44),
.B2(n_24),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_136),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_75),
.A2(n_32),
.B1(n_30),
.B2(n_38),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_67),
.B(n_39),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_140),
.B(n_1),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_56),
.A2(n_44),
.B1(n_42),
.B2(n_41),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_142),
.A2(n_160),
.B1(n_2),
.B2(n_3),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_50),
.A2(n_30),
.B1(n_38),
.B2(n_39),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_144),
.A2(n_150),
.B1(n_86),
.B2(n_2),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_42),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_52),
.A2(n_38),
.B1(n_30),
.B2(n_37),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_69),
.B(n_37),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_151),
.B(n_63),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_53),
.B(n_41),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_76),
.A2(n_24),
.B1(n_18),
.B2(n_25),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_25),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_161),
.B(n_162),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_18),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_100),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_163),
.B(n_170),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_80),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_164),
.B(n_175),
.Y(n_246)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_165),
.Y(n_253)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_95),
.B(n_51),
.C(n_79),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_166),
.A2(n_112),
.B(n_157),
.C(n_101),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_168),
.B(n_195),
.Y(n_242)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_114),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_172),
.B(n_193),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_173),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_59),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_191),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_115),
.B(n_87),
.Y(n_175)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_176),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_177),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_103),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_178),
.B(n_182),
.Y(n_257)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_109),
.B1(n_97),
.B2(n_68),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g264 ( 
.A1(n_180),
.A2(n_183),
.B1(n_188),
.B2(n_196),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_108),
.B(n_87),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_70),
.B1(n_71),
.B2(n_129),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_184),
.B(n_11),
.Y(n_260)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_186),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_187),
.Y(n_270)
);

OA22x2_ASAP7_75t_SL g188 ( 
.A1(n_132),
.A2(n_90),
.B1(n_88),
.B2(n_54),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_154),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_54),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_192),
.B(n_198),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_149),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_128),
.B1(n_126),
.B2(n_138),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_127),
.B(n_1),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_199),
.A2(n_110),
.B1(n_143),
.B2(n_9),
.Y(n_241)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_200),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_120),
.B(n_13),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_120),
.B(n_3),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_203),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_122),
.B(n_3),
.Y(n_203)
);

OR2x2_ASAP7_75t_SL g204 ( 
.A(n_156),
.B(n_3),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_204),
.B(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_146),
.Y(n_205)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_205),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_4),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_206),
.B(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_122),
.B(n_4),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_208),
.B(n_217),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_5),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_130),
.B(n_5),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_211),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_119),
.B(n_6),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_125),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_141),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_213),
.A2(n_144),
.B1(n_117),
.B2(n_113),
.Y(n_225)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_119),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_102),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_112),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_133),
.B(n_7),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_110),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_137),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_219),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_162),
.A2(n_150),
.B(n_118),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_223),
.A2(n_230),
.B(n_252),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_245),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_219),
.A2(n_102),
.B1(n_126),
.B2(n_106),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_197),
.A2(n_152),
.B(n_121),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_166),
.A2(n_152),
.B(n_121),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_231),
.A2(n_169),
.B(n_185),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_234),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_167),
.A2(n_170),
.B1(n_188),
.B2(n_168),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_237),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_198),
.A2(n_138),
.B1(n_128),
.B2(n_133),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_238),
.A2(n_189),
.B1(n_176),
.B2(n_187),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_241),
.B(n_231),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_243),
.B(n_248),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_174),
.A2(n_157),
.B1(n_101),
.B2(n_9),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_186),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_188),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_195),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_184),
.B(n_11),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_268),
.C(n_165),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_191),
.B(n_13),
.C(n_192),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_195),
.A2(n_13),
.B1(n_190),
.B2(n_193),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_269),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_177),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_212),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_272),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_163),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_273),
.B(n_279),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_240),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_274),
.B(n_276),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_275),
.B(n_297),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_240),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_214),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_161),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_280),
.B(n_281),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_210),
.Y(n_281)
);

O2A1O1Ixp33_ASAP7_75t_SL g282 ( 
.A1(n_247),
.A2(n_223),
.B(n_252),
.C(n_264),
.Y(n_282)
);

OA21x2_ASAP7_75t_L g345 ( 
.A1(n_282),
.A2(n_301),
.B(n_307),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_242),
.A2(n_194),
.B1(n_209),
.B2(n_211),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_283),
.A2(n_268),
.B1(n_243),
.B2(n_264),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_171),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_284),
.B(n_285),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_206),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_220),
.B(n_171),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_286),
.B(n_267),
.C(n_297),
.Y(n_359)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_222),
.B(n_201),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_287),
.Y(n_357)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_288),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_204),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_295),
.Y(n_322)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_290),
.Y(n_333)
);

AOI22x1_ASAP7_75t_L g293 ( 
.A1(n_225),
.A2(n_201),
.B1(n_215),
.B2(n_216),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_293),
.A2(n_307),
.B1(n_310),
.B2(n_311),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_220),
.B(n_200),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_296),
.A2(n_301),
.B(n_313),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_257),
.B(n_207),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_300),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_224),
.B(n_205),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_230),
.B(n_242),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_303),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_228),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_304),
.B(n_306),
.Y(n_354)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_251),
.Y(n_305)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_255),
.B(n_179),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_221),
.B(n_271),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_308),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_222),
.B(n_181),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_309),
.B(n_312),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_247),
.A2(n_173),
.B1(n_187),
.B2(n_232),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_260),
.B(n_173),
.Y(n_312)
);

A2O1A1O1Ixp25_ASAP7_75t_L g313 ( 
.A1(n_249),
.A2(n_173),
.B(n_187),
.C(n_239),
.D(n_242),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_233),
.Y(n_314)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_234),
.A2(n_243),
.B(n_261),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_315),
.A2(n_318),
.B(n_313),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_235),
.Y(n_316)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_316),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_254),
.Y(n_317)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_229),
.B(n_249),
.Y(n_319)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_319),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_302),
.A2(n_245),
.B1(n_229),
.B2(n_264),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_320),
.A2(n_331),
.B(n_335),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_316),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_324),
.B(n_305),
.Y(n_391)
);

AO21x2_ASAP7_75t_L g325 ( 
.A1(n_294),
.A2(n_226),
.B(n_264),
.Y(n_325)
);

OA22x2_ASAP7_75t_L g366 ( 
.A1(n_325),
.A2(n_345),
.B1(n_350),
.B2(n_355),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_326),
.B(n_332),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_315),
.A2(n_266),
.B(n_241),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_302),
.A2(n_251),
.B1(n_244),
.B2(n_256),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_301),
.A2(n_258),
.B(n_254),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_294),
.A2(n_244),
.B1(n_256),
.B2(n_235),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_353),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_293),
.A2(n_248),
.B1(n_250),
.B2(n_228),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_343),
.A2(n_346),
.B1(n_298),
.B2(n_317),
.Y(n_392)
);

OAI22xp33_ASAP7_75t_L g346 ( 
.A1(n_282),
.A2(n_270),
.B1(n_267),
.B2(n_250),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_283),
.A2(n_309),
.B1(n_295),
.B2(n_319),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_282),
.A2(n_233),
.B1(n_236),
.B2(n_265),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_292),
.A2(n_236),
.B1(n_265),
.B2(n_270),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_277),
.Y(n_356)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_356),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_312),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_292),
.A2(n_267),
.B1(n_296),
.B2(n_281),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_298),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_361),
.A2(n_289),
.B(n_293),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_330),
.B(n_275),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_362),
.B(n_358),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_340),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_363),
.B(n_377),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_337),
.A2(n_318),
.B1(n_291),
.B2(n_274),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_365),
.A2(n_370),
.B(n_347),
.Y(n_400)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_323),
.Y(n_368)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_368),
.Y(n_405)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_369),
.Y(n_411)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_323),
.Y(n_371)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_371),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_376),
.C(n_387),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_321),
.B(n_286),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_373),
.Y(n_418)
);

XOR2x2_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_280),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_374),
.Y(n_415)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_327),
.Y(n_375)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_375),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_322),
.B(n_287),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_276),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_327),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_378),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_328),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_381),
.Y(n_399)
);

BUFx24_ASAP7_75t_SL g381 ( 
.A(n_339),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_338),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_382),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_384),
.Y(n_413)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_333),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_354),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_385),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_335),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_386),
.A2(n_388),
.B1(n_390),
.B2(n_392),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_322),
.B(n_287),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_304),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_285),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_389),
.B(n_391),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_329),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_278),
.C(n_288),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_342),
.C(n_303),
.Y(n_423)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_394),
.A2(n_395),
.B1(n_356),
.B2(n_334),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_351),
.B(n_290),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_367),
.A2(n_351),
.B1(n_325),
.B2(n_345),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_397),
.A2(n_398),
.B1(n_404),
.B2(n_408),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_383),
.A2(n_353),
.B1(n_341),
.B2(n_357),
.Y(n_398)
);

NAND3xp33_ASAP7_75t_SL g440 ( 
.A(n_400),
.B(n_422),
.C(n_413),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_367),
.A2(n_325),
.B1(n_345),
.B2(n_361),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_380),
.A2(n_357),
.B1(n_332),
.B2(n_347),
.Y(n_408)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_410),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_364),
.A2(n_325),
.B1(n_331),
.B2(n_346),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_412),
.A2(n_380),
.B1(n_366),
.B2(n_384),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_417),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_365),
.A2(n_325),
.B1(n_320),
.B2(n_326),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_416),
.A2(n_421),
.B1(n_397),
.B2(n_412),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_362),
.B(n_358),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_370),
.A2(n_350),
.B1(n_360),
.B2(n_334),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_364),
.A2(n_342),
.B(n_355),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_423),
.B(n_393),
.C(n_372),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_395),
.A2(n_336),
.B(n_338),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_424),
.B(n_375),
.Y(n_431)
);

NOR2x1_ASAP7_75t_L g426 ( 
.A(n_420),
.B(n_389),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_426),
.B(n_405),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_435),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_378),
.Y(n_429)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_429),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_431),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_407),
.B(n_374),
.Y(n_432)
);

NAND3xp33_ASAP7_75t_L g461 ( 
.A(n_432),
.B(n_439),
.C(n_441),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_376),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_436),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_387),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_366),
.Y(n_436)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_437),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_366),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_406),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_396),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_440),
.A2(n_419),
.B(n_411),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_403),
.B(n_348),
.Y(n_441)
);

NAND3xp33_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_394),
.C(n_371),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_418),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_368),
.Y(n_443)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_443),
.Y(n_463)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_420),
.Y(n_444)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_445),
.A2(n_449),
.B1(n_421),
.B2(n_416),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_404),
.A2(n_366),
.B1(n_382),
.B2(n_369),
.Y(n_446)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_446),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_336),
.C(n_314),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_406),
.C(n_419),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_401),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_448),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_408),
.A2(n_398),
.B1(n_422),
.B2(n_415),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_424),
.B(n_402),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_450),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_465),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_453),
.A2(n_430),
.B1(n_447),
.B2(n_448),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_449),
.A2(n_400),
.B(n_405),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_458),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_457),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_443),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_462),
.B(n_469),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_450),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_470),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_466),
.B(n_427),
.C(n_434),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_474),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_435),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_473),
.B(n_479),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_436),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_480),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_460),
.B(n_433),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_458),
.B(n_433),
.C(n_438),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_454),
.B(n_426),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_481),
.B(n_483),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_411),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_428),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_484),
.B(n_485),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_459),
.B(n_445),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_468),
.A2(n_429),
.B1(n_446),
.B2(n_437),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_486),
.A2(n_462),
.B1(n_463),
.B2(n_469),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_476),
.A2(n_464),
.B1(n_455),
.B2(n_468),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_488),
.B(n_494),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_471),
.B(n_455),
.C(n_465),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_491),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_475),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_456),
.C(n_451),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_496),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_482),
.A2(n_464),
.B1(n_467),
.B2(n_463),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_470),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_498),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_497),
.A2(n_478),
.B1(n_452),
.B2(n_472),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_502),
.B1(n_493),
.B2(n_495),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_492),
.B(n_477),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_501),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_491),
.A2(n_480),
.B(n_479),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_490),
.B(n_452),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_487),
.Y(n_507)
);

CKINVDCx14_ASAP7_75t_R g512 ( 
.A(n_507),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_L g508 ( 
.A(n_499),
.B(n_489),
.Y(n_508)
);

AO21x1_ASAP7_75t_L g514 ( 
.A1(n_508),
.A2(n_509),
.B(n_511),
.Y(n_514)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_505),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_510),
.B(n_503),
.Y(n_513)
);

NAND3xp33_ASAP7_75t_SL g515 ( 
.A(n_513),
.B(n_504),
.C(n_501),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_514),
.A2(n_504),
.B(n_498),
.Y(n_516)
);

NAND3xp33_ASAP7_75t_L g517 ( 
.A(n_515),
.B(n_516),
.C(n_512),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_517),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_518),
.B(n_486),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_519),
.B(n_495),
.Y(n_520)
);


endmodule