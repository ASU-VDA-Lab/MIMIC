module fake_netlist_5_164_n_1704 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1704);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1704;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1644;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1495;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_86),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_97),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_152),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_106),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_58),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_49),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_88),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_109),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_155),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_35),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_153),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_1),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_67),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_5),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_62),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_135),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_57),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_90),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_49),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_44),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_111),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_70),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_115),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_83),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_38),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_124),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_64),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_126),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_27),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_23),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_99),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_101),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_102),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_77),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_50),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_30),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_79),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_31),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_40),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_53),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_46),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_6),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_65),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_7),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_134),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_39),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_33),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_114),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_5),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_131),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_23),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_137),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_93),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_9),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_132),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_30),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_19),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_54),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_6),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_112),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_128),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_14),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_91),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_47),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_156),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_148),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_34),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_2),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_4),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_41),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_129),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_110),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_75),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_130),
.Y(n_248)
);

CKINVDCx11_ASAP7_75t_R g249 ( 
.A(n_71),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_141),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_11),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_157),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_54),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_22),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_10),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_105),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_7),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_1),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_32),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_96),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_120),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_17),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_59),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_104),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_140),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_68),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_72),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_117),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_123),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_163),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_66),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_92),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_147),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_43),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_63),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_165),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_143),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_21),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_76),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_122),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_44),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_84),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_2),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_95),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_107),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_25),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_133),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_29),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_138),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_0),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_3),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_11),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_36),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_145),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_46),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_159),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_56),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_103),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_60),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_81),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_80),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_39),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_61),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_149),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_136),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_48),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_38),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_98),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_18),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_31),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_73),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_45),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_160),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_87),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_94),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_119),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_43),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_113),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_36),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_16),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_74),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_150),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_32),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_56),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_16),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_33),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_27),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_8),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_69),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_53),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_13),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_15),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_189),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_189),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_224),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_179),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_328),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_325),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_195),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_170),
.Y(n_340)
);

NOR2xp67_ASAP7_75t_L g341 ( 
.A(n_173),
.B(n_0),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_332),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_238),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_208),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_178),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_182),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_268),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_196),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_201),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_205),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_186),
.B(n_3),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_168),
.B(n_4),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_168),
.B(n_8),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_249),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_205),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_199),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_277),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_212),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_213),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_214),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_211),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_216),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_223),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_304),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_215),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_217),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_232),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_255),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_219),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_171),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_170),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_200),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_259),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_203),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_206),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_262),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_207),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_283),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_221),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_286),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_222),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_170),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_290),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_237),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_228),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_225),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_193),
.B(n_9),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g390 ( 
.A(n_243),
.B(n_10),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_292),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_178),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_237),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_230),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_309),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_330),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_172),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_181),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_229),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_246),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_194),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_231),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_233),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_197),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_237),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_248),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_236),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_287),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_256),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_204),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_260),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_193),
.B(n_12),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_210),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_242),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_244),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_251),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_218),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_226),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_397),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_374),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_340),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_340),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_336),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_398),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_404),
.Y(n_426)
);

NOR2x1_ASAP7_75t_L g427 ( 
.A(n_408),
.B(n_227),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_R g428 ( 
.A(n_356),
.B(n_263),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_339),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_376),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_377),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_340),
.Y(n_432)
);

NAND2xp33_ASAP7_75t_SL g433 ( 
.A(n_338),
.B(n_342),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_340),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_349),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_373),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_379),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_364),
.B(n_209),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_392),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_381),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_373),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_373),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_373),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_373),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_384),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_365),
.B(n_241),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_384),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_344),
.Y(n_448)
);

NOR2x1_ASAP7_75t_L g449 ( 
.A(n_408),
.B(n_234),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_R g450 ( 
.A(n_388),
.B(n_264),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_384),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_357),
.B(n_243),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_410),
.Y(n_453)
);

NAND2x1_ASAP7_75t_L g454 ( 
.A(n_384),
.B(n_279),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_R g456 ( 
.A(n_344),
.B(n_166),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_348),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_413),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_372),
.B(n_279),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_350),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_351),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_352),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_399),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_363),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_400),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_335),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_406),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_359),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_369),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_417),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_370),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_375),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_378),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_380),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_R g475 ( 
.A(n_409),
.B(n_265),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_411),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_352),
.B(n_253),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_358),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_366),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_391),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_R g483 ( 
.A(n_360),
.B(n_266),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_338),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_395),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_342),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_333),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_334),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_360),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_355),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_337),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_361),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_347),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_361),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_439),
.B(n_362),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_491),
.B(n_175),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_462),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_462),
.B(n_401),
.Y(n_499)
);

AND3x2_ASAP7_75t_L g500 ( 
.A(n_448),
.B(n_412),
.C(n_354),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_421),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_483),
.Y(n_502)
);

AND3x2_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_353),
.C(n_235),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_491),
.B(n_346),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_459),
.A2(n_389),
.B1(n_253),
.B2(n_310),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_452),
.B(n_418),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_468),
.Y(n_507)
);

BUFx8_ASAP7_75t_SL g508 ( 
.A(n_424),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_421),
.Y(n_509)
);

NAND3xp33_ASAP7_75t_L g510 ( 
.A(n_452),
.B(n_367),
.C(n_362),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_367),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_450),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_491),
.B(n_346),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_421),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_466),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_419),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_425),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_459),
.B(n_175),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_421),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_459),
.B(n_368),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_426),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_459),
.B(n_368),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_421),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_423),
.B(n_434),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_490),
.B(n_371),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_479),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_477),
.B(n_240),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_479),
.B(n_235),
.Y(n_530)
);

AND3x4_ASAP7_75t_L g531 ( 
.A(n_427),
.B(n_341),
.C(n_390),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_484),
.B(n_371),
.Y(n_532)
);

INVx4_ASAP7_75t_SL g533 ( 
.A(n_443),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_453),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_477),
.B(n_245),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_495),
.B(n_343),
.Y(n_537)
);

AND2x6_ASAP7_75t_L g538 ( 
.A(n_449),
.B(n_315),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_L g539 ( 
.A(n_458),
.B(n_416),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_494),
.B(n_383),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_488),
.B(n_383),
.Y(n_541)
);

INVx4_ASAP7_75t_SL g542 ( 
.A(n_443),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_485),
.B(n_315),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_488),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_471),
.A2(n_310),
.B1(n_239),
.B2(n_308),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_489),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_429),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_446),
.A2(n_306),
.B1(n_324),
.B2(n_297),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_494),
.B(n_345),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_SL g550 ( 
.A(n_456),
.B(n_387),
.Y(n_550)
);

INVx4_ASAP7_75t_SL g551 ( 
.A(n_443),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_489),
.Y(n_552)
);

BUFx4f_ASAP7_75t_L g553 ( 
.A(n_485),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_485),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_443),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_446),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_455),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_444),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_444),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_492),
.B(n_387),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_485),
.B(n_394),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_485),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_423),
.B(n_394),
.Y(n_563)
);

OAI22x1_ASAP7_75t_L g564 ( 
.A1(n_438),
.A2(n_320),
.B1(n_188),
.B2(n_302),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_470),
.B(n_402),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g566 ( 
.A(n_433),
.B(n_403),
.C(n_402),
.Y(n_566)
);

INVxp67_ASAP7_75t_SL g567 ( 
.A(n_423),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_471),
.B(n_170),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_438),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_435),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_444),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_471),
.B(n_170),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_434),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_454),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_L g575 ( 
.A(n_486),
.B(n_403),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_470),
.B(n_239),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_454),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_486),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_434),
.B(n_407),
.Y(n_579)
);

INVx6_ASAP7_75t_L g580 ( 
.A(n_444),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_457),
.B(n_239),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_460),
.A2(n_308),
.B1(n_294),
.B2(n_269),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_460),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_461),
.A2(n_416),
.B1(n_415),
.B2(n_414),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_444),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_442),
.B(n_407),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_461),
.A2(n_269),
.B1(n_239),
.B2(n_294),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_445),
.Y(n_588)
);

CKINVDCx6p67_ASAP7_75t_R g589 ( 
.A(n_480),
.Y(n_589)
);

CKINVDCx6p67_ASAP7_75t_R g590 ( 
.A(n_440),
.Y(n_590)
);

INVxp67_ASAP7_75t_SL g591 ( 
.A(n_447),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_445),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_447),
.B(n_415),
.Y(n_593)
);

INVxp33_ASAP7_75t_SL g594 ( 
.A(n_428),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_467),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_447),
.B(n_174),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_478),
.B(n_386),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_464),
.B(n_239),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_445),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_464),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_420),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_445),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_L g603 ( 
.A(n_469),
.B(n_269),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_472),
.B(n_269),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_445),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_472),
.Y(n_606)
);

OAI21xp33_ASAP7_75t_L g607 ( 
.A1(n_473),
.A2(n_220),
.B(n_202),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_473),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_474),
.B(n_269),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_420),
.Y(n_610)
);

INVxp33_ASAP7_75t_L g611 ( 
.A(n_474),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_481),
.B(n_393),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_L g613 ( 
.A(n_481),
.B(n_293),
.C(n_288),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_430),
.B(n_405),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_482),
.Y(n_615)
);

INVxp33_ASAP7_75t_L g616 ( 
.A(n_487),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_451),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_487),
.A2(n_294),
.B1(n_308),
.B2(n_247),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_451),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_478),
.B(n_250),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_422),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_430),
.B(n_252),
.Y(n_622)
);

INVx5_ASAP7_75t_L g623 ( 
.A(n_451),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_422),
.A2(n_308),
.B1(n_294),
.B2(n_261),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_432),
.B(n_166),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_432),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_436),
.B(n_267),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_431),
.B(n_281),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_431),
.A2(n_295),
.B1(n_287),
.B2(n_326),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_436),
.B(n_270),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_451),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_437),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_451),
.B(n_294),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_437),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_463),
.Y(n_635)
);

AND2x6_ASAP7_75t_L g636 ( 
.A(n_463),
.B(n_308),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_504),
.B(n_513),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_504),
.A2(n_284),
.B1(n_271),
.B2(n_272),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_574),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_635),
.B(n_282),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_506),
.B(n_298),
.Y(n_641)
);

O2A1O1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_519),
.A2(n_311),
.B(n_314),
.C(n_329),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_537),
.B(n_465),
.Y(n_643)
);

NOR2xp67_ASAP7_75t_L g644 ( 
.A(n_512),
.B(n_465),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_506),
.B(n_511),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_521),
.B(n_307),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_574),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_544),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_506),
.B(n_300),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_523),
.B(n_476),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_561),
.B(n_305),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_546),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_611),
.B(n_167),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_561),
.B(n_322),
.Y(n_654)
);

BUFx8_ASAP7_75t_L g655 ( 
.A(n_610),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_552),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_L g657 ( 
.A(n_510),
.B(n_560),
.C(n_541),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_597),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_499),
.B(n_277),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_550),
.A2(n_276),
.B1(n_273),
.B2(n_275),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_565),
.A2(n_280),
.B1(n_285),
.B2(n_289),
.Y(n_661)
);

BUFx10_ASAP7_75t_L g662 ( 
.A(n_526),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_548),
.B(n_476),
.C(n_278),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_628),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_507),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_608),
.Y(n_666)
);

NOR2xp67_ASAP7_75t_L g667 ( 
.A(n_502),
.B(n_169),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_608),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_616),
.B(n_277),
.Y(n_669)
);

NOR2x1p5_ASAP7_75t_L g670 ( 
.A(n_589),
.B(n_180),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_616),
.B(n_277),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_505),
.A2(n_277),
.B1(n_327),
.B2(n_326),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_583),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_541),
.B(n_169),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_497),
.A2(n_176),
.B(n_177),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_600),
.B(n_176),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g677 ( 
.A(n_629),
.B(n_274),
.C(n_258),
.Y(n_677)
);

INVxp67_ASAP7_75t_SL g678 ( 
.A(n_514),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_553),
.A2(n_296),
.B(n_183),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_606),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_R g681 ( 
.A(n_601),
.B(n_183),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_508),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_540),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_615),
.B(n_184),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_565),
.B(n_184),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_560),
.B(n_277),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_516),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_SL g688 ( 
.A(n_594),
.B(n_517),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_625),
.B(n_185),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_518),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_505),
.A2(n_331),
.B1(n_327),
.B2(n_323),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_522),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_498),
.B(n_185),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_498),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_496),
.B(n_187),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_577),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_526),
.B(n_187),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_625),
.B(n_190),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_567),
.B(n_190),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_591),
.B(n_191),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_612),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_547),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_532),
.B(n_254),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_635),
.B(n_287),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_534),
.B(n_528),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_612),
.A2(n_303),
.B1(n_191),
.B2(n_321),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_528),
.A2(n_303),
.B1(n_192),
.B2(n_321),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_618),
.A2(n_331),
.B1(n_323),
.B2(n_320),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_515),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_528),
.B(n_301),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_530),
.B(n_301),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_530),
.B(n_299),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_536),
.B(n_299),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_549),
.B(n_578),
.Y(n_714)
);

O2A1O1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_497),
.A2(n_192),
.B(n_318),
.C(n_198),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_536),
.B(n_198),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_582),
.A2(n_319),
.B(n_180),
.C(n_317),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_536),
.B(n_318),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_584),
.B(n_296),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_577),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_620),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_620),
.Y(n_722)
);

NOR2xp67_ASAP7_75t_SL g723 ( 
.A(n_582),
.B(n_313),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_620),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_596),
.B(n_313),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_539),
.B(n_257),
.C(n_316),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_621),
.B(n_316),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_549),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_545),
.B(n_319),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_549),
.B(n_317),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_626),
.B(n_312),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_535),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_627),
.B(n_312),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_535),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_545),
.B(n_302),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_557),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_630),
.B(n_188),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_556),
.B(n_12),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_563),
.A2(n_164),
.B1(n_144),
.B2(n_142),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_579),
.A2(n_139),
.B1(n_127),
.B2(n_125),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_586),
.B(n_13),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_557),
.Y(n_742)
);

NAND3xp33_ASAP7_75t_L g743 ( 
.A(n_613),
.B(n_14),
.C(n_15),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_587),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_744)
);

AOI221xp5_ASAP7_75t_L g745 ( 
.A1(n_564),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.C(n_24),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_593),
.B(n_20),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_554),
.B(n_116),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_566),
.B(n_24),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_580),
.Y(n_749)
);

O2A1O1Ixp5_ASAP7_75t_L g750 ( 
.A1(n_568),
.A2(n_108),
.B(n_89),
.C(n_85),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_580),
.Y(n_751)
);

AOI22x1_ASAP7_75t_L g752 ( 
.A1(n_558),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_618),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_553),
.B(n_82),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_573),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_562),
.B(n_78),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_587),
.A2(n_34),
.B(n_35),
.C(n_37),
.Y(n_757)
);

NOR2x1p5_ASAP7_75t_L g758 ( 
.A(n_590),
.B(n_37),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_573),
.B(n_55),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_580),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_501),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_525),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_503),
.Y(n_763)
);

AND2x2_ASAP7_75t_SL g764 ( 
.A(n_624),
.B(n_41),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_558),
.B(n_42),
.Y(n_765)
);

AOI221xp5_ASAP7_75t_L g766 ( 
.A1(n_607),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.C(n_48),
.Y(n_766)
);

NOR3xp33_ASAP7_75t_L g767 ( 
.A(n_575),
.B(n_50),
.C(n_51),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_624),
.B(n_51),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_531),
.A2(n_52),
.B1(n_55),
.B2(n_538),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_571),
.B(n_585),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_531),
.A2(n_538),
.B1(n_636),
.B2(n_572),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_572),
.Y(n_772)
);

O2A1O1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_598),
.A2(n_609),
.B(n_543),
.C(n_576),
.Y(n_773)
);

AND2x2_ASAP7_75t_SL g774 ( 
.A(n_614),
.B(n_634),
.Y(n_774)
);

AND2x6_ASAP7_75t_L g775 ( 
.A(n_585),
.B(n_619),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_592),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_701),
.B(n_500),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_721),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_657),
.B(n_527),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_664),
.B(n_632),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_764),
.A2(n_538),
.B1(n_636),
.B2(n_633),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_637),
.A2(n_543),
.B(n_633),
.C(n_603),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_674),
.B(n_538),
.Y(n_783)
);

AO22x1_ASAP7_75t_L g784 ( 
.A1(n_748),
.A2(n_569),
.B1(n_538),
.B2(n_604),
.Y(n_784)
);

BUFx2_ASAP7_75t_SL g785 ( 
.A(n_644),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_674),
.B(n_527),
.Y(n_786)
);

OAI321xp33_ASAP7_75t_L g787 ( 
.A1(n_769),
.A2(n_622),
.A3(n_631),
.B1(n_619),
.B2(n_617),
.C(n_602),
.Y(n_787)
);

NAND2x1p5_ASAP7_75t_L g788 ( 
.A(n_639),
.B(n_524),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_744),
.A2(n_602),
.B(n_599),
.C(n_592),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_696),
.A2(n_622),
.B1(n_617),
.B2(n_555),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_714),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_683),
.B(n_622),
.Y(n_792)
);

AOI21x1_ASAP7_75t_L g793 ( 
.A1(n_770),
.A2(n_555),
.B(n_529),
.Y(n_793)
);

O2A1O1Ixp5_ASAP7_75t_L g794 ( 
.A1(n_686),
.A2(n_529),
.B(n_581),
.C(n_604),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_639),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_639),
.B(n_570),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_665),
.Y(n_797)
);

AOI33xp33_ASAP7_75t_L g798 ( 
.A1(n_691),
.A2(n_595),
.A3(n_604),
.B1(n_581),
.B2(n_533),
.B3(n_542),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_722),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_709),
.B(n_588),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_696),
.A2(n_720),
.B1(n_764),
.B2(n_771),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_639),
.B(n_588),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_646),
.B(n_514),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_724),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_646),
.B(n_520),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_658),
.A2(n_520),
.B1(n_588),
.B2(n_604),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_648),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_650),
.B(n_520),
.Y(n_808)
);

BUFx12f_ASAP7_75t_L g809 ( 
.A(n_655),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_647),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_685),
.B(n_653),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_665),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_647),
.B(n_551),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_659),
.A2(n_581),
.B1(n_604),
.B2(n_551),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_734),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_720),
.A2(n_771),
.B1(n_705),
.B2(n_641),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_703),
.B(n_542),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_647),
.B(n_662),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_678),
.A2(n_509),
.B(n_559),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_762),
.A2(n_559),
.B(n_605),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_689),
.B(n_581),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_698),
.B(n_581),
.Y(n_822)
);

AND2x2_ASAP7_75t_SL g823 ( 
.A(n_769),
.B(n_559),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_647),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_649),
.A2(n_654),
.B1(n_651),
.B2(n_753),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_652),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_662),
.B(n_605),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_774),
.B(n_623),
.Y(n_828)
);

BUFx8_ASAP7_75t_L g829 ( 
.A(n_702),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_711),
.A2(n_623),
.B(n_712),
.C(n_746),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_656),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_673),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_753),
.A2(n_766),
.B1(n_768),
.B2(n_748),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_738),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_680),
.B(n_741),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_741),
.B(n_746),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_734),
.Y(n_837)
);

NOR3xp33_ASAP7_75t_L g838 ( 
.A(n_719),
.B(n_697),
.C(n_663),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_772),
.A2(n_712),
.B1(n_711),
.B2(n_666),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_725),
.B(n_668),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_688),
.B(n_774),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_693),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_733),
.B(n_737),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_687),
.B(n_690),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_692),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_775),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_669),
.B(n_671),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_669),
.B(n_671),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_775),
.Y(n_849)
);

AOI21xp33_ASAP7_75t_L g850 ( 
.A1(n_719),
.A2(n_697),
.B(n_695),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_754),
.A2(n_756),
.B(n_747),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_730),
.B(n_695),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_699),
.B(n_700),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_776),
.A2(n_773),
.B(n_761),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_694),
.B(n_638),
.Y(n_855)
);

BUFx8_ASAP7_75t_L g856 ( 
.A(n_763),
.Y(n_856)
);

AO22x1_ASAP7_75t_L g857 ( 
.A1(n_677),
.A2(n_767),
.B1(n_728),
.B2(n_693),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_710),
.A2(n_716),
.B1(n_718),
.B2(n_713),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_736),
.Y(n_859)
);

AOI21x1_ASAP7_75t_L g860 ( 
.A1(n_736),
.A2(n_742),
.B(n_732),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_676),
.B(n_684),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_675),
.B(n_661),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_643),
.B(n_706),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_759),
.A2(n_731),
.B(n_750),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_727),
.B(n_723),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_744),
.A2(n_757),
.B(n_768),
.C(n_717),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_640),
.A2(n_726),
.B1(n_707),
.B2(n_660),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_694),
.B(n_667),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_749),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_751),
.Y(n_870)
);

INVxp67_ASAP7_75t_L g871 ( 
.A(n_640),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_765),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_760),
.A2(n_642),
.B(n_715),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_717),
.A2(n_729),
.B(n_735),
.Y(n_874)
);

BUFx12f_ASAP7_75t_L g875 ( 
.A(n_655),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_729),
.B(n_735),
.Y(n_876)
);

NAND3xp33_ASAP7_75t_L g877 ( 
.A(n_691),
.B(n_672),
.C(n_708),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_679),
.B(n_672),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_640),
.B(n_775),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_775),
.A2(n_704),
.B1(n_743),
.B2(n_740),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_704),
.B(n_708),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_775),
.A2(n_704),
.B1(n_739),
.B2(n_745),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_757),
.A2(n_752),
.B(n_681),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_670),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_758),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_681),
.B(n_682),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_664),
.Y(n_887)
);

OAI21xp33_ASAP7_75t_L g888 ( 
.A1(n_674),
.A2(n_691),
.B(n_646),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_665),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_645),
.A2(n_637),
.B(n_659),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_674),
.A2(n_711),
.B(n_712),
.C(n_645),
.Y(n_891)
);

AND2x2_ASAP7_75t_SL g892 ( 
.A(n_764),
.B(n_769),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_701),
.B(n_664),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_755),
.A2(n_645),
.B(n_553),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_637),
.A2(n_645),
.B1(n_657),
.B2(n_674),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_653),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_645),
.B(n_637),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_721),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_694),
.B(n_498),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_714),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_755),
.A2(n_645),
.B(n_553),
.Y(n_901)
);

AOI21xp33_ASAP7_75t_L g902 ( 
.A1(n_674),
.A2(n_657),
.B(n_646),
.Y(n_902)
);

NAND2xp33_ASAP7_75t_L g903 ( 
.A(n_639),
.B(n_647),
.Y(n_903)
);

NOR3xp33_ASAP7_75t_L g904 ( 
.A(n_657),
.B(n_674),
.C(n_719),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_674),
.A2(n_711),
.B(n_712),
.C(n_645),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_664),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_755),
.A2(n_645),
.B(n_553),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_701),
.B(n_664),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_645),
.B(n_637),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_694),
.B(n_498),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_674),
.B(n_712),
.C(n_711),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_665),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_764),
.A2(n_769),
.B1(n_753),
.B2(n_766),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_645),
.B(n_637),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_645),
.B(n_637),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_645),
.A2(n_637),
.B(n_659),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_721),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_645),
.A2(n_657),
.B1(n_637),
.B2(n_674),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_755),
.A2(n_645),
.B(n_553),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_645),
.B(n_637),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_755),
.A2(n_645),
.B(n_553),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_755),
.A2(n_645),
.B(n_553),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_764),
.A2(n_769),
.B1(n_753),
.B2(n_766),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_755),
.A2(n_645),
.B(n_553),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_645),
.B(n_637),
.Y(n_925)
);

OAI21xp33_ASAP7_75t_L g926 ( 
.A1(n_674),
.A2(n_691),
.B(n_646),
.Y(n_926)
);

BUFx8_ASAP7_75t_L g927 ( 
.A(n_702),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_755),
.A2(n_645),
.B(n_553),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_637),
.A2(n_645),
.B(n_757),
.C(n_744),
.Y(n_929)
);

BUFx4f_ASAP7_75t_L g930 ( 
.A(n_714),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_702),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_755),
.A2(n_645),
.B(n_553),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_755),
.A2(n_645),
.B(n_553),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_755),
.A2(n_645),
.B(n_553),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_755),
.A2(n_645),
.B(n_553),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_721),
.Y(n_936)
);

OAI221xp5_ASAP7_75t_L g937 ( 
.A1(n_657),
.A2(n_674),
.B1(n_646),
.B2(n_672),
.C(n_769),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_911),
.A2(n_905),
.B(n_891),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_795),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_811),
.B(n_896),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_899),
.B(n_910),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_896),
.B(n_843),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_807),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_846),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_826),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_793),
.A2(n_860),
.B(n_854),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_899),
.B(n_910),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_900),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_791),
.B(n_887),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_795),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_913),
.A2(n_923),
.B1(n_937),
.B2(n_892),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_930),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_836),
.B(n_888),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_897),
.A2(n_914),
.B(n_909),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_892),
.A2(n_913),
.B1(n_923),
.B2(n_877),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_834),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_930),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_926),
.B(n_835),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_795),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_797),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_823),
.B(n_895),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_887),
.Y(n_962)
);

AO21x1_ASAP7_75t_L g963 ( 
.A1(n_902),
.A2(n_904),
.B(n_918),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_894),
.A2(n_907),
.B(n_901),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_861),
.B(n_904),
.Y(n_965)
);

AOI21x1_ASAP7_75t_L g966 ( 
.A1(n_919),
.A2(n_922),
.B(n_921),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_852),
.B(n_908),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_915),
.A2(n_925),
.B(n_920),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_853),
.B(n_786),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_890),
.A2(n_916),
.B(n_851),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_833),
.A2(n_862),
.B1(n_801),
.B2(n_823),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_924),
.A2(n_932),
.B(n_935),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_786),
.B(n_840),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_831),
.Y(n_974)
);

AO31x2_ASAP7_75t_L g975 ( 
.A1(n_830),
.A2(n_825),
.A3(n_816),
.B(n_839),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_928),
.A2(n_933),
.B(n_934),
.Y(n_976)
);

INVxp67_ASAP7_75t_SL g977 ( 
.A(n_903),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_833),
.A2(n_850),
.B(n_881),
.C(n_866),
.Y(n_978)
);

AOI21x1_ASAP7_75t_SL g979 ( 
.A1(n_783),
.A2(n_878),
.B(n_822),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_812),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_832),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_795),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_908),
.B(n_893),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_858),
.B(n_808),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_881),
.B(n_863),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_780),
.B(n_863),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_842),
.B(n_871),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_845),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_R g989 ( 
.A(n_886),
.B(n_829),
.Y(n_989)
);

AOI21x1_ASAP7_75t_L g990 ( 
.A1(n_803),
.A2(n_805),
.B(n_821),
.Y(n_990)
);

AOI21x1_ASAP7_75t_L g991 ( 
.A1(n_865),
.A2(n_802),
.B(n_873),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_866),
.A2(n_787),
.B(n_929),
.C(n_838),
.Y(n_992)
);

OA21x2_ASAP7_75t_L g993 ( 
.A1(n_864),
.A2(n_874),
.B(n_883),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_871),
.B(n_936),
.Y(n_994)
);

AOI221xp5_ASAP7_75t_L g995 ( 
.A1(n_838),
.A2(n_929),
.B1(n_777),
.B2(n_844),
.C(n_841),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_815),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_847),
.A2(n_848),
.B(n_876),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_782),
.A2(n_855),
.B(n_872),
.Y(n_998)
);

OAI21x1_ASAP7_75t_SL g999 ( 
.A1(n_879),
.A2(n_789),
.B(n_868),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_837),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_794),
.A2(n_788),
.B(n_819),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_882),
.A2(n_781),
.B1(n_880),
.B2(n_867),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_906),
.B(n_931),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_782),
.A2(n_808),
.B(n_781),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_906),
.B(n_796),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_846),
.B(n_849),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_859),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_889),
.A2(n_912),
.B(n_778),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_885),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_817),
.A2(n_790),
.B(n_779),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_820),
.A2(n_813),
.B(n_824),
.Y(n_1011)
);

OA21x2_ASAP7_75t_L g1012 ( 
.A1(n_799),
.A2(n_917),
.B(n_898),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_804),
.B(n_800),
.Y(n_1013)
);

NAND2xp33_ASAP7_75t_L g1014 ( 
.A(n_846),
.B(n_849),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_814),
.A2(n_798),
.B(n_828),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_810),
.A2(n_824),
.B(n_869),
.Y(n_1016)
);

AO31x2_ASAP7_75t_L g1017 ( 
.A1(n_777),
.A2(n_792),
.A3(n_870),
.B(n_884),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_810),
.B(n_784),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_857),
.A2(n_818),
.B(n_806),
.Y(n_1019)
);

OA21x2_ASAP7_75t_L g1020 ( 
.A1(n_827),
.A2(n_792),
.B(n_846),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_849),
.A2(n_785),
.B(n_829),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_849),
.A2(n_856),
.B(n_927),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_927),
.A2(n_856),
.B(n_809),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_875),
.B(n_811),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_L g1025 ( 
.A(n_888),
.B(n_926),
.C(n_911),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_888),
.B(n_926),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_829),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_797),
.Y(n_1028)
);

AOI21x1_ASAP7_75t_SL g1029 ( 
.A1(n_783),
.A2(n_878),
.B(n_836),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_811),
.B(n_896),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_811),
.B(n_896),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_846),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_852),
.B(n_664),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_897),
.A2(n_914),
.B(n_909),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_897),
.A2(n_914),
.B(n_909),
.Y(n_1035)
);

AO21x1_ASAP7_75t_L g1036 ( 
.A1(n_836),
.A2(n_902),
.B(n_904),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_811),
.B(n_896),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_911),
.A2(n_905),
.B(n_891),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_888),
.B(n_926),
.Y(n_1039)
);

AND2x6_ASAP7_75t_L g1040 ( 
.A(n_846),
.B(n_849),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_811),
.B(n_896),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_899),
.B(n_910),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_913),
.A2(n_923),
.B(n_926),
.C(n_888),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_793),
.A2(n_860),
.B(n_854),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_897),
.A2(n_914),
.B(n_909),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_852),
.B(n_664),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_807),
.Y(n_1047)
);

NAND2x1_ASAP7_75t_L g1048 ( 
.A(n_795),
.B(n_775),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_897),
.A2(n_914),
.B(n_909),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_811),
.B(n_896),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_811),
.B(n_896),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_897),
.A2(n_914),
.B(n_909),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_897),
.A2(n_914),
.B(n_909),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_911),
.A2(n_905),
.B(n_891),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_913),
.A2(n_923),
.B(n_926),
.C(n_888),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_811),
.B(n_896),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_911),
.A2(n_905),
.B(n_891),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_911),
.A2(n_905),
.B(n_891),
.Y(n_1058)
);

OA22x2_ASAP7_75t_L g1059 ( 
.A1(n_888),
.A2(n_926),
.B1(n_548),
.B2(n_664),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_811),
.B(n_896),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_797),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_897),
.A2(n_914),
.B(n_909),
.Y(n_1062)
);

OAI22x1_ASAP7_75t_L g1063 ( 
.A1(n_877),
.A2(n_881),
.B1(n_863),
.B2(n_786),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_897),
.A2(n_914),
.B(n_909),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_931),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_911),
.A2(n_905),
.B(n_891),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_811),
.B(n_896),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_897),
.A2(n_914),
.B(n_909),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_900),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_897),
.A2(n_914),
.B(n_909),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_811),
.B(n_896),
.Y(n_1071)
);

OAI22x1_ASAP7_75t_L g1072 ( 
.A1(n_877),
.A2(n_881),
.B1(n_863),
.B2(n_786),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_941),
.B(n_947),
.Y(n_1073)
);

INVx5_ASAP7_75t_L g1074 ( 
.A(n_1040),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_965),
.B(n_942),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_969),
.B(n_986),
.Y(n_1076)
);

BUFx4f_ASAP7_75t_SL g1077 ( 
.A(n_1027),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_941),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_985),
.A2(n_955),
.B1(n_973),
.B2(n_951),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_985),
.B(n_983),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_947),
.B(n_1042),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_995),
.A2(n_1072),
.B1(n_1063),
.B2(n_1002),
.Y(n_1082)
);

AND2x6_ASAP7_75t_L g1083 ( 
.A(n_944),
.B(n_1032),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_949),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_967),
.B(n_1033),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1046),
.B(n_1059),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_943),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_945),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1059),
.B(n_940),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_1065),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1030),
.B(n_1031),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_974),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_1003),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_944),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_955),
.A2(n_978),
.B1(n_1055),
.B2(n_1043),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_948),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_1042),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1037),
.B(n_1041),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_995),
.A2(n_1039),
.B1(n_1026),
.B2(n_1024),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_954),
.A2(n_1034),
.B(n_1062),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_SL g1101 ( 
.A(n_1069),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_989),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_944),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_954),
.A2(n_1034),
.B(n_1035),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_SL g1105 ( 
.A(n_1036),
.B(n_963),
.C(n_978),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1050),
.B(n_1051),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_L g1107 ( 
.A(n_1025),
.B(n_1055),
.C(n_1043),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_989),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_968),
.A2(n_1068),
.B(n_1035),
.Y(n_1109)
);

INVx5_ASAP7_75t_L g1110 ( 
.A(n_1040),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_962),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_956),
.Y(n_1112)
);

AOI21xp33_ASAP7_75t_SL g1113 ( 
.A1(n_1005),
.A2(n_957),
.B(n_952),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1045),
.A2(n_1053),
.B(n_1049),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_994),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_SL g1116 ( 
.A(n_1022),
.B(n_1009),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_994),
.B(n_987),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1056),
.B(n_1060),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_1032),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1032),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_987),
.B(n_1021),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1067),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_981),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1045),
.A2(n_1068),
.B(n_1064),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_982),
.B(n_1032),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_988),
.Y(n_1126)
);

AND2x6_ASAP7_75t_L g1127 ( 
.A(n_1026),
.B(n_1039),
.Y(n_1127)
);

CKINVDCx16_ASAP7_75t_R g1128 ( 
.A(n_982),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_1071),
.Y(n_1129)
);

NAND2x1p5_ASAP7_75t_L g1130 ( 
.A(n_939),
.B(n_950),
.Y(n_1130)
);

OR2x6_ASAP7_75t_L g1131 ( 
.A(n_1023),
.B(n_1019),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1047),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_953),
.B(n_1049),
.Y(n_1133)
);

AND2x6_ASAP7_75t_L g1134 ( 
.A(n_939),
.B(n_950),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1040),
.Y(n_1135)
);

OR2x6_ASAP7_75t_L g1136 ( 
.A(n_1019),
.B(n_1010),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1017),
.B(n_1013),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_960),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_980),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_996),
.Y(n_1140)
);

NAND2x1p5_ASAP7_75t_L g1141 ( 
.A(n_959),
.B(n_1048),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_1040),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_992),
.A2(n_971),
.B1(n_961),
.B2(n_984),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1017),
.B(n_938),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_958),
.B(n_961),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1000),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1007),
.Y(n_1147)
);

NOR2x1_ASAP7_75t_L g1148 ( 
.A(n_959),
.B(n_1006),
.Y(n_1148)
);

NOR2x1_ASAP7_75t_L g1149 ( 
.A(n_1006),
.B(n_1014),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1028),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_1017),
.B(n_997),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1052),
.B(n_1070),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1052),
.B(n_1070),
.Y(n_1153)
);

AND2x6_ASAP7_75t_L g1154 ( 
.A(n_1018),
.B(n_1061),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_992),
.A2(n_1054),
.B1(n_1066),
.B2(n_1038),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_1020),
.Y(n_1156)
);

OAI221xp5_ASAP7_75t_L g1157 ( 
.A1(n_1057),
.A2(n_1058),
.B1(n_998),
.B2(n_1015),
.C(n_1010),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_1020),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1016),
.Y(n_1159)
);

CKINVDCx11_ASAP7_75t_R g1160 ( 
.A(n_1017),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_1008),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_993),
.B(n_1004),
.Y(n_1162)
);

OAI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_1004),
.A2(n_990),
.B(n_991),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_975),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1011),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_993),
.A2(n_976),
.B1(n_972),
.B2(n_964),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_999),
.B(n_972),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1001),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_1029),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_975),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_975),
.B(n_946),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1044),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_975),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_966),
.Y(n_1174)
);

AND2x2_ASAP7_75t_SL g1175 ( 
.A(n_1029),
.B(n_979),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_944),
.Y(n_1176)
);

AND2x2_ASAP7_75t_SL g1177 ( 
.A(n_955),
.B(n_892),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_941),
.B(n_947),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1065),
.Y(n_1179)
);

INVx8_ASAP7_75t_L g1180 ( 
.A(n_941),
.Y(n_1180)
);

NAND2x1p5_ASAP7_75t_L g1181 ( 
.A(n_1065),
.B(n_941),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_956),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_986),
.B(n_967),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_969),
.B(n_942),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_969),
.B(n_942),
.Y(n_1185)
);

NOR2xp67_ASAP7_75t_L g1186 ( 
.A(n_952),
.B(n_512),
.Y(n_1186)
);

AND2x6_ASAP7_75t_L g1187 ( 
.A(n_944),
.B(n_1032),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1012),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_986),
.B(n_967),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_986),
.B(n_969),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_985),
.A2(n_888),
.B1(n_926),
.B2(n_904),
.Y(n_1191)
);

AOI21xp33_ASAP7_75t_SL g1192 ( 
.A1(n_1059),
.A2(n_438),
.B(n_548),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_992),
.A2(n_977),
.B(n_1002),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_1027),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_969),
.B(n_942),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_SL g1196 ( 
.A1(n_1026),
.A2(n_786),
.B(n_777),
.C(n_674),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1012),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1012),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_986),
.B(n_967),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_949),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1012),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_949),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_985),
.A2(n_926),
.B(n_888),
.C(n_911),
.Y(n_1203)
);

OR2x6_ASAP7_75t_L g1204 ( 
.A(n_1065),
.B(n_952),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_970),
.A2(n_755),
.B(n_851),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_986),
.B(n_969),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1012),
.Y(n_1207)
);

BUFx12f_ASAP7_75t_L g1208 ( 
.A(n_1112),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1126),
.Y(n_1209)
);

OAI22x1_ASAP7_75t_SL g1210 ( 
.A1(n_1102),
.A2(n_1108),
.B1(n_1194),
.B2(n_1122),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1080),
.A2(n_1129),
.B1(n_1206),
.B2(n_1190),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1177),
.A2(n_1079),
.B1(n_1155),
.B2(n_1127),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1090),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1179),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_1093),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1099),
.A2(n_1185),
.B1(n_1184),
.B2(n_1195),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1203),
.A2(n_1191),
.B(n_1143),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1197),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1200),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1082),
.A2(n_1193),
.B(n_1157),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_1100),
.A2(n_1109),
.B(n_1104),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1089),
.B(n_1107),
.Y(n_1222)
);

NAND2x1p5_ASAP7_75t_L g1223 ( 
.A(n_1074),
.B(n_1110),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1076),
.A2(n_1075),
.B1(n_1118),
.B2(n_1098),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1088),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1106),
.B(n_1183),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1127),
.A2(n_1095),
.B1(n_1105),
.B2(n_1145),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1077),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1127),
.A2(n_1189),
.B1(n_1199),
.B2(n_1086),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1114),
.A2(n_1124),
.B(n_1205),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1091),
.B(n_1085),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1147),
.A2(n_1084),
.B1(n_1161),
.B2(n_1115),
.Y(n_1232)
);

CKINVDCx6p67_ASAP7_75t_R g1233 ( 
.A(n_1101),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1132),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1087),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1202),
.A2(n_1123),
.B1(n_1113),
.B2(n_1182),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1092),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1110),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1111),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_1180),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1133),
.A2(n_1196),
.B(n_1127),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1168),
.A2(n_1152),
.B(n_1153),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1136),
.A2(n_1163),
.B(n_1175),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1188),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1188),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1110),
.Y(n_1246)
);

CKINVDCx11_ASAP7_75t_R g1247 ( 
.A(n_1204),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1181),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1138),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1139),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1146),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1121),
.B(n_1131),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1150),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1136),
.A2(n_1137),
.B1(n_1170),
.B2(n_1144),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1140),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1128),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1167),
.A2(n_1166),
.B(n_1162),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1198),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1173),
.A2(n_1131),
.B1(n_1164),
.B2(n_1154),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1096),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1117),
.B(n_1192),
.Y(n_1261)
);

CKINVDCx11_ASAP7_75t_R g1262 ( 
.A(n_1204),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1164),
.A2(n_1154),
.B1(n_1121),
.B2(n_1160),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1151),
.B(n_1158),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1186),
.A2(n_1149),
.B1(n_1101),
.B2(n_1167),
.Y(n_1265)
);

BUFx2_ASAP7_75t_SL g1266 ( 
.A(n_1073),
.Y(n_1266)
);

BUFx8_ASAP7_75t_L g1267 ( 
.A(n_1078),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1201),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1078),
.A2(n_1097),
.B1(n_1081),
.B2(n_1178),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1078),
.A2(n_1097),
.B1(n_1081),
.B2(n_1178),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1207),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1116),
.A2(n_1154),
.B1(n_1180),
.B2(n_1097),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1154),
.A2(n_1171),
.B1(n_1073),
.B2(n_1207),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1094),
.Y(n_1274)
);

AO21x1_ASAP7_75t_L g1275 ( 
.A1(n_1172),
.A2(n_1159),
.B(n_1141),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1103),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1148),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1103),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1130),
.Y(n_1279)
);

BUFx8_ASAP7_75t_L g1280 ( 
.A(n_1142),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1103),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1169),
.A2(n_1174),
.B(n_1156),
.Y(n_1282)
);

CKINVDCx11_ASAP7_75t_R g1283 ( 
.A(n_1119),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_SL g1284 ( 
.A(n_1119),
.Y(n_1284)
);

INVx6_ASAP7_75t_L g1285 ( 
.A(n_1119),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1169),
.A2(n_1135),
.B1(n_1125),
.B2(n_1176),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1120),
.Y(n_1287)
);

INVx6_ASAP7_75t_L g1288 ( 
.A(n_1120),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1120),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1083),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1165),
.A2(n_1083),
.B(n_1187),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1134),
.A2(n_1165),
.B1(n_1187),
.B2(n_1083),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1134),
.A2(n_913),
.B1(n_923),
.B2(n_892),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_1187),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1187),
.Y(n_1295)
);

CKINVDCx11_ASAP7_75t_R g1296 ( 
.A(n_1194),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1075),
.B(n_1200),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1074),
.B(n_1110),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1200),
.Y(n_1299)
);

BUFx2_ASAP7_75t_SL g1300 ( 
.A(n_1101),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1080),
.A2(n_892),
.B1(n_985),
.B2(n_786),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1112),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1180),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1080),
.A2(n_892),
.B1(n_985),
.B2(n_786),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1080),
.B(n_1190),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1080),
.A2(n_888),
.B1(n_926),
.B2(n_985),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1180),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1193),
.A2(n_1104),
.B(n_1100),
.Y(n_1308)
);

AOI21xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1122),
.A2(n_601),
.B(n_430),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1075),
.B(n_1200),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1074),
.B(n_1110),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1126),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1100),
.A2(n_1109),
.B(n_1104),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1296),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1308),
.A2(n_1220),
.B(n_1257),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1222),
.B(n_1264),
.Y(n_1316)
);

BUFx8_ASAP7_75t_SL g1317 ( 
.A(n_1228),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1291),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1296),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1217),
.A2(n_1212),
.B1(n_1301),
.B2(n_1304),
.Y(n_1320)
);

AO21x2_ASAP7_75t_L g1321 ( 
.A1(n_1241),
.A2(n_1243),
.B(n_1230),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1244),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1245),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1211),
.B(n_1305),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1258),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1297),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1222),
.B(n_1264),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1291),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_1228),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1252),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1268),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1252),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1254),
.B(n_1271),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1254),
.B(n_1227),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1227),
.B(n_1209),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1242),
.A2(n_1273),
.B(n_1259),
.Y(n_1336)
);

INVxp67_ASAP7_75t_R g1337 ( 
.A(n_1210),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1282),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1273),
.A2(n_1259),
.B(n_1275),
.Y(n_1339)
);

AOI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1265),
.A2(n_1216),
.B(n_1313),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1280),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1310),
.B(n_1218),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1280),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1224),
.B(n_1231),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1221),
.Y(n_1345)
);

INVx11_ASAP7_75t_L g1346 ( 
.A(n_1280),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1299),
.B(n_1226),
.Y(n_1347)
);

OA21x2_ASAP7_75t_L g1348 ( 
.A1(n_1263),
.A2(n_1306),
.B(n_1312),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1249),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1293),
.A2(n_1277),
.B(n_1237),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1235),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1263),
.B(n_1229),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1250),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1219),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1229),
.B(n_1225),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1251),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1253),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_1223),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1234),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1255),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1292),
.A2(n_1311),
.B(n_1223),
.Y(n_1361)
);

INVx6_ASAP7_75t_L g1362 ( 
.A(n_1267),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1232),
.B(n_1215),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1306),
.B(n_1274),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1290),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1295),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1236),
.B(n_1261),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1272),
.A2(n_1286),
.B(n_1311),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1289),
.A2(n_1279),
.B(n_1294),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1267),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1238),
.B(n_1246),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1331),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1333),
.B(n_1336),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1336),
.B(n_1287),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1333),
.B(n_1214),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1345),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1344),
.B(n_1238),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1344),
.B(n_1246),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1336),
.B(n_1246),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1336),
.B(n_1281),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1315),
.B(n_1321),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1318),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1335),
.B(n_1214),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1314),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1315),
.B(n_1276),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1335),
.B(n_1349),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1324),
.A2(n_1320),
.B1(n_1334),
.B2(n_1367),
.Y(n_1387)
);

OR2x6_ASAP7_75t_L g1388 ( 
.A(n_1361),
.B(n_1298),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1328),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1322),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1325),
.Y(n_1391)
);

INVxp67_ASAP7_75t_L g1392 ( 
.A(n_1369),
.Y(n_1392)
);

INVx4_ASAP7_75t_R g1393 ( 
.A(n_1341),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1367),
.B(n_1239),
.Y(n_1394)
);

INVxp33_ASAP7_75t_L g1395 ( 
.A(n_1347),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1316),
.B(n_1266),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1338),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1334),
.B(n_1354),
.C(n_1309),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1316),
.B(n_1285),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1369),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1327),
.B(n_1285),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1340),
.A2(n_1269),
.B(n_1270),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1327),
.B(n_1288),
.Y(n_1403)
);

OAI21xp33_ASAP7_75t_L g1404 ( 
.A1(n_1352),
.A2(n_1302),
.B(n_1248),
.Y(n_1404)
);

AOI31xp33_ASAP7_75t_L g1405 ( 
.A1(n_1368),
.A2(n_1303),
.A3(n_1240),
.B(n_1307),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1338),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1323),
.B(n_1285),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1338),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1394),
.B(n_1326),
.Y(n_1409)
);

NAND3xp33_ASAP7_75t_L g1410 ( 
.A(n_1387),
.B(n_1354),
.C(n_1366),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1395),
.B(n_1326),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1395),
.B(n_1377),
.Y(n_1412)
);

OAI21xp33_ASAP7_75t_L g1413 ( 
.A1(n_1387),
.A2(n_1352),
.B(n_1355),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1398),
.A2(n_1368),
.B1(n_1348),
.B2(n_1381),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1405),
.A2(n_1363),
.B(n_1364),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_R g1416 ( 
.A(n_1384),
.B(n_1329),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1398),
.B(n_1319),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1378),
.B(n_1342),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1378),
.B(n_1394),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_L g1420 ( 
.A(n_1381),
.B(n_1404),
.C(n_1405),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1383),
.B(n_1342),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1374),
.B(n_1339),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1374),
.B(n_1339),
.Y(n_1423)
);

NAND3xp33_ASAP7_75t_L g1424 ( 
.A(n_1381),
.B(n_1366),
.C(n_1365),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1383),
.B(n_1356),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1375),
.B(n_1356),
.Y(n_1426)
);

AND2x2_ASAP7_75t_SL g1427 ( 
.A(n_1373),
.B(n_1339),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1372),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1404),
.B(n_1358),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1386),
.B(n_1356),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1386),
.B(n_1357),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1373),
.A2(n_1363),
.B1(n_1348),
.B2(n_1362),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1376),
.Y(n_1433)
);

NOR3xp33_ASAP7_75t_L g1434 ( 
.A(n_1402),
.B(n_1340),
.C(n_1371),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1407),
.B(n_1357),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_R g1436 ( 
.A(n_1384),
.B(n_1256),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1399),
.A2(n_1355),
.B1(n_1364),
.B2(n_1348),
.Y(n_1437)
);

NOR3xp33_ASAP7_75t_SL g1438 ( 
.A(n_1402),
.B(n_1371),
.C(n_1365),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1380),
.B(n_1350),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1407),
.B(n_1357),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1372),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1407),
.B(n_1351),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_L g1443 ( 
.A(n_1392),
.B(n_1359),
.C(n_1360),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1390),
.B(n_1350),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1379),
.B(n_1350),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1385),
.B(n_1350),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1399),
.B(n_1351),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1399),
.B(n_1353),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1401),
.B(n_1403),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1401),
.B(n_1353),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1396),
.A2(n_1330),
.B1(n_1332),
.B2(n_1348),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1419),
.B(n_1390),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1433),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1412),
.B(n_1391),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1428),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1430),
.B(n_1431),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1428),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1441),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1441),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1422),
.B(n_1373),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1427),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1426),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1444),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1422),
.B(n_1423),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1444),
.Y(n_1465)
);

AND2x4_ASAP7_75t_SL g1466 ( 
.A(n_1438),
.B(n_1388),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1446),
.B(n_1400),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1427),
.B(n_1397),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1427),
.B(n_1406),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_SL g1470 ( 
.A(n_1410),
.B(n_1384),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1424),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1442),
.Y(n_1472)
);

INVxp67_ASAP7_75t_SL g1473 ( 
.A(n_1443),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1443),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1435),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1439),
.B(n_1445),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1439),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1446),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1432),
.B(n_1408),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1440),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1424),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1455),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1455),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1458),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1452),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1457),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1471),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1461),
.B(n_1389),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1458),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1467),
.B(n_1411),
.Y(n_1490)
);

NAND2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1461),
.B(n_1389),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1467),
.B(n_1418),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1457),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1461),
.B(n_1389),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1457),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1476),
.B(n_1389),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1452),
.B(n_1409),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1457),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1462),
.B(n_1447),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1459),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1476),
.B(n_1389),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1462),
.B(n_1448),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1459),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1459),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1475),
.B(n_1450),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1476),
.B(n_1389),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1453),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1475),
.B(n_1421),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1469),
.B(n_1389),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1453),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1480),
.B(n_1425),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1460),
.B(n_1432),
.Y(n_1512)
);

CKINVDCx8_ASAP7_75t_R g1513 ( 
.A(n_1470),
.Y(n_1513)
);

NOR2xp67_ASAP7_75t_L g1514 ( 
.A(n_1471),
.B(n_1420),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1453),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1469),
.B(n_1382),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1469),
.B(n_1389),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1480),
.B(n_1449),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1453),
.Y(n_1519)
);

INVxp67_ASAP7_75t_SL g1520 ( 
.A(n_1473),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1482),
.Y(n_1521)
);

NAND2x1p5_ASAP7_75t_L g1522 ( 
.A(n_1514),
.B(n_1481),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1487),
.B(n_1472),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1520),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1497),
.B(n_1485),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1499),
.B(n_1502),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1509),
.B(n_1464),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1505),
.B(n_1472),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1486),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1513),
.A2(n_1420),
.B1(n_1414),
.B2(n_1415),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1482),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1488),
.B(n_1473),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1484),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1486),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1484),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1489),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1511),
.B(n_1474),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1508),
.B(n_1474),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1509),
.B(n_1464),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1488),
.B(n_1468),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1483),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1493),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1517),
.B(n_1464),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1517),
.B(n_1477),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1491),
.A2(n_1470),
.B(n_1417),
.Y(n_1545)
);

CKINVDCx16_ASAP7_75t_R g1546 ( 
.A(n_1494),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1513),
.B(n_1384),
.Y(n_1547)
);

O2A1O1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1491),
.A2(n_1481),
.B(n_1415),
.C(n_1434),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1518),
.B(n_1456),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1490),
.B(n_1492),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1490),
.B(n_1456),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1493),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1492),
.B(n_1481),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1496),
.B(n_1477),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1491),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1512),
.B(n_1460),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1489),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1512),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1495),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1494),
.B(n_1454),
.Y(n_1560)
);

NAND4xp25_ASAP7_75t_L g1561 ( 
.A(n_1496),
.B(n_1410),
.C(n_1413),
.D(n_1437),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1503),
.B(n_1460),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1495),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1521),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1547),
.B(n_1317),
.Y(n_1565)
);

INVx3_ASAP7_75t_SL g1566 ( 
.A(n_1546),
.Y(n_1566)
);

AND3x1_ASAP7_75t_L g1567 ( 
.A(n_1545),
.B(n_1548),
.C(n_1525),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1521),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1527),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1522),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1531),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1527),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1540),
.B(n_1516),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1522),
.B(n_1362),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1546),
.B(n_1516),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1522),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1524),
.B(n_1538),
.Y(n_1577)
);

INVxp67_ASAP7_75t_SL g1578 ( 
.A(n_1558),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1553),
.B(n_1463),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1532),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1539),
.B(n_1516),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1531),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1553),
.B(n_1463),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1540),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1533),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1530),
.A2(n_1413),
.B(n_1337),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1533),
.Y(n_1587)
);

AO21x2_ASAP7_75t_L g1588 ( 
.A1(n_1563),
.A2(n_1500),
.B(n_1498),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1537),
.B(n_1501),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1539),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1561),
.A2(n_1466),
.B1(n_1479),
.B2(n_1468),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1535),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1535),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1532),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1550),
.B(n_1465),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1526),
.B(n_1501),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1536),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1532),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1536),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1578),
.B(n_1532),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1566),
.B(n_1549),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1566),
.B(n_1551),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1567),
.A2(n_1540),
.B1(n_1466),
.B2(n_1523),
.Y(n_1603)
);

NOR2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1577),
.B(n_1208),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1584),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1596),
.B(n_1560),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1586),
.A2(n_1591),
.B1(n_1574),
.B2(n_1575),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1584),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1580),
.Y(n_1609)
);

AOI322xp5_ASAP7_75t_L g1610 ( 
.A1(n_1570),
.A2(n_1576),
.A3(n_1575),
.B1(n_1590),
.B2(n_1569),
.C1(n_1572),
.C2(n_1598),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1584),
.B(n_1540),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1571),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1588),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1581),
.B(n_1543),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1565),
.B(n_1594),
.Y(n_1615)
);

NAND2x1_ASAP7_75t_L g1616 ( 
.A(n_1574),
.B(n_1555),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1574),
.A2(n_1556),
.B1(n_1437),
.B2(n_1466),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1571),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1581),
.B(n_1543),
.Y(n_1619)
);

OAI321xp33_ASAP7_75t_L g1620 ( 
.A1(n_1574),
.A2(n_1556),
.A3(n_1557),
.B1(n_1528),
.B2(n_1429),
.C(n_1544),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1569),
.A2(n_1466),
.B1(n_1436),
.B2(n_1541),
.Y(n_1621)
);

NAND2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1573),
.B(n_1370),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1573),
.A2(n_1555),
.B1(n_1477),
.B2(n_1478),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1582),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1573),
.B(n_1544),
.Y(n_1625)
);

NOR2x1_ASAP7_75t_L g1626 ( 
.A(n_1605),
.B(n_1582),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1611),
.B(n_1572),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1609),
.B(n_1590),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1612),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1618),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1624),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1605),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1610),
.B(n_1602),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1601),
.B(n_1589),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1600),
.B(n_1564),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1608),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1608),
.B(n_1606),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1611),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1622),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1614),
.B(n_1568),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1614),
.B(n_1585),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1625),
.B(n_1595),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1625),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1622),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1613),
.Y(n_1645)
);

NOR3xp33_ASAP7_75t_L g1646 ( 
.A(n_1633),
.B(n_1615),
.C(n_1607),
.Y(n_1646)
);

AOI322xp5_ASAP7_75t_L g1647 ( 
.A1(n_1626),
.A2(n_1615),
.A3(n_1603),
.B1(n_1621),
.B2(n_1619),
.C1(n_1613),
.C2(n_1616),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_SL g1648 ( 
.A(n_1639),
.B(n_1621),
.C(n_1617),
.Y(n_1648)
);

NOR4xp25_ASAP7_75t_SL g1649 ( 
.A(n_1638),
.B(n_1620),
.C(n_1593),
.D(n_1599),
.Y(n_1649)
);

AOI311xp33_ASAP7_75t_L g1650 ( 
.A1(n_1632),
.A2(n_1623),
.A3(n_1587),
.B(n_1599),
.C(n_1593),
.Y(n_1650)
);

O2A1O1Ixp5_ASAP7_75t_L g1651 ( 
.A1(n_1643),
.A2(n_1587),
.B(n_1597),
.C(n_1592),
.Y(n_1651)
);

AOI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1635),
.A2(n_1643),
.B1(n_1640),
.B2(n_1641),
.C(n_1634),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_SL g1653 ( 
.A1(n_1644),
.A2(n_1628),
.B(n_1642),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1629),
.A2(n_1595),
.B1(n_1557),
.B2(n_1555),
.C(n_1583),
.Y(n_1654)
);

AOI222xp33_ASAP7_75t_L g1655 ( 
.A1(n_1630),
.A2(n_1604),
.B1(n_1479),
.B2(n_1468),
.C1(n_1554),
.C2(n_1563),
.Y(n_1655)
);

OAI211xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1628),
.A2(n_1260),
.B(n_1262),
.C(n_1247),
.Y(n_1656)
);

NOR3xp33_ASAP7_75t_L g1657 ( 
.A(n_1636),
.B(n_1262),
.C(n_1247),
.Y(n_1657)
);

NOR3xp33_ASAP7_75t_L g1658 ( 
.A(n_1646),
.B(n_1637),
.C(n_1631),
.Y(n_1658)
);

NOR3xp33_ASAP7_75t_L g1659 ( 
.A(n_1653),
.B(n_1637),
.C(n_1645),
.Y(n_1659)
);

AOI211xp5_ASAP7_75t_L g1660 ( 
.A1(n_1648),
.A2(n_1642),
.B(n_1627),
.C(n_1645),
.Y(n_1660)
);

AO22x1_ASAP7_75t_L g1661 ( 
.A1(n_1657),
.A2(n_1627),
.B1(n_1213),
.B2(n_1370),
.Y(n_1661)
);

OAI322xp33_ASAP7_75t_L g1662 ( 
.A1(n_1649),
.A2(n_1583),
.A3(n_1579),
.B1(n_1627),
.B2(n_1562),
.C1(n_1534),
.C2(n_1552),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1656),
.A2(n_1554),
.B1(n_1337),
.B2(n_1579),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1651),
.Y(n_1664)
);

NOR3xp33_ASAP7_75t_L g1665 ( 
.A(n_1652),
.B(n_1654),
.C(n_1647),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1655),
.B(n_1208),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1650),
.B(n_1233),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1653),
.B(n_1506),
.Y(n_1668)
);

NAND3x1_ASAP7_75t_SL g1669 ( 
.A(n_1662),
.B(n_1233),
.C(n_1300),
.Y(n_1669)
);

OAI211xp5_ASAP7_75t_L g1670 ( 
.A1(n_1665),
.A2(n_1416),
.B(n_1283),
.C(n_1256),
.Y(n_1670)
);

NAND4xp75_ASAP7_75t_L g1671 ( 
.A(n_1664),
.B(n_1479),
.C(n_1506),
.D(n_1534),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1667),
.B(n_1213),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1660),
.B(n_1529),
.Y(n_1673)
);

NOR3xp33_ASAP7_75t_L g1674 ( 
.A(n_1658),
.B(n_1283),
.C(n_1240),
.Y(n_1674)
);

NAND4xp25_ASAP7_75t_L g1675 ( 
.A(n_1666),
.B(n_1370),
.C(n_1343),
.D(n_1341),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1673),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1671),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1675),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1670),
.B(n_1659),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1672),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1674),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1669),
.B(n_1668),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1670),
.B(n_1661),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1677),
.A2(n_1663),
.B1(n_1529),
.B2(n_1542),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1676),
.B(n_1679),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1678),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1680),
.B(n_1562),
.Y(n_1687)
);

OR5x1_ASAP7_75t_L g1688 ( 
.A(n_1682),
.B(n_1588),
.C(n_1542),
.D(n_1552),
.E(n_1559),
.Y(n_1688)
);

NAND4xp25_ASAP7_75t_L g1689 ( 
.A(n_1683),
.B(n_1341),
.C(n_1343),
.D(n_1451),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1687),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1686),
.B(n_1681),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1688),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1690),
.Y(n_1693)
);

NOR3xp33_ASAP7_75t_L g1694 ( 
.A(n_1693),
.B(n_1691),
.C(n_1685),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1694),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1694),
.A2(n_1682),
.B1(n_1684),
.B2(n_1689),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1696),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1695),
.B(n_1692),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1698),
.A2(n_1588),
.B(n_1559),
.Y(n_1699)
);

AOI21x1_ASAP7_75t_L g1700 ( 
.A1(n_1697),
.A2(n_1510),
.B(n_1507),
.Y(n_1700)
);

AOI222xp33_ASAP7_75t_L g1701 ( 
.A1(n_1699),
.A2(n_1519),
.B1(n_1515),
.B2(n_1507),
.C1(n_1510),
.C2(n_1498),
.Y(n_1701)
);

OAI33xp33_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1700),
.A3(n_1519),
.B1(n_1515),
.B2(n_1500),
.B3(n_1504),
.Y(n_1702)
);

OAI221xp5_ASAP7_75t_R g1703 ( 
.A1(n_1702),
.A2(n_1278),
.B1(n_1346),
.B2(n_1393),
.C(n_1284),
.Y(n_1703)
);

AOI211xp5_ASAP7_75t_L g1704 ( 
.A1(n_1703),
.A2(n_1343),
.B(n_1303),
.C(n_1307),
.Y(n_1704)
);


endmodule