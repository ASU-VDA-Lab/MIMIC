module fake_jpeg_2112_n_365 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_365);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_365;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_48),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_20),
.B(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_56),
.Y(n_104)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_28),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_67),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_12),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_69),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_74),
.B1(n_75),
.B2(n_78),
.Y(n_90)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_15),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_76),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_79),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_15),
.B(n_31),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_21),
.B1(n_40),
.B2(n_18),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_84),
.A2(n_96),
.B1(n_100),
.B2(n_102),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_28),
.B1(n_33),
.B2(n_19),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_92),
.A2(n_99),
.B1(n_103),
.B2(n_110),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_29),
.B1(n_37),
.B2(n_35),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_42),
.A2(n_28),
.B1(n_15),
.B2(n_31),
.Y(n_97)
);

AO22x1_ASAP7_75t_L g161 ( 
.A1(n_97),
.A2(n_91),
.B1(n_93),
.B2(n_101),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_27),
.B(n_29),
.C(n_35),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_105),
.B(n_82),
.C(n_88),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_43),
.A2(n_28),
.B1(n_33),
.B2(n_24),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_45),
.A2(n_40),
.B1(n_21),
.B2(n_31),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_40),
.B1(n_21),
.B2(n_31),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_48),
.A2(n_33),
.B1(n_19),
.B2(n_24),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_60),
.A2(n_27),
.B(n_37),
.C(n_22),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_53),
.B1(n_58),
.B2(n_46),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_78),
.B1(n_6),
.B2(n_7),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_24),
.B1(n_19),
.B2(n_38),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_62),
.A2(n_39),
.B1(n_22),
.B2(n_15),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_113),
.B1(n_123),
.B2(n_124),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_72),
.A2(n_39),
.B1(n_40),
.B2(n_21),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_100),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_32),
.B1(n_13),
.B2(n_10),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_54),
.B(n_0),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_91),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_63),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_75),
.A2(n_13),
.B1(n_32),
.B2(n_4),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_117),
.B1(n_102),
.B2(n_126),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_44),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_61),
.A2(n_55),
.B1(n_70),
.B2(n_5),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_55),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_91),
.B1(n_86),
.B2(n_87),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_69),
.B1(n_65),
.B2(n_68),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_131),
.A2(n_142),
.B1(n_160),
.B2(n_161),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_132),
.B(n_135),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_13),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_133),
.B(n_154),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_4),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_69),
.B(n_74),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_137),
.A2(n_155),
.B(n_157),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_104),
.B(n_6),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_141),
.B(n_143),
.Y(n_213)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_146),
.A2(n_153),
.B1(n_156),
.B2(n_174),
.Y(n_212)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_147),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_109),
.B(n_94),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_151),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_84),
.A2(n_109),
.B1(n_108),
.B2(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_83),
.B(n_86),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_95),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_156),
.B(n_159),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_98),
.A2(n_105),
.B(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_87),
.B(n_120),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_162),
.Y(n_177)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_106),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_167),
.Y(n_178)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_97),
.A2(n_93),
.B1(n_101),
.B2(n_115),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_131),
.B(n_161),
.C(n_142),
.Y(n_181)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_115),
.B(n_101),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_89),
.B(n_97),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_169),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_89),
.B(n_127),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_97),
.B(n_121),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_172),
.C(n_137),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_128),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_118),
.A2(n_64),
.B1(n_28),
.B2(n_33),
.Y(n_173)
);

AO21x1_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_176),
.B(n_146),
.Y(n_192)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_90),
.B(n_114),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_153),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_114),
.A2(n_122),
.B1(n_94),
.B2(n_117),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_175),
.A2(n_171),
.B1(n_168),
.B2(n_161),
.Y(n_180)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_180),
.B(n_181),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_167),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_190),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_189),
.B(n_201),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_157),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_197),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_192),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_SL g195 ( 
.A(n_151),
.B(n_143),
.C(n_160),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_195),
.B(n_138),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_166),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_176),
.A2(n_134),
.B1(n_145),
.B2(n_151),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_152),
.A2(n_140),
.B1(n_165),
.B2(n_135),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_202),
.A2(n_212),
.B1(n_147),
.B2(n_149),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_136),
.B(n_163),
.C(n_139),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_199),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_141),
.B(n_152),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_206),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_144),
.B(n_159),
.Y(n_206)
);

AND2x6_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_164),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_147),
.Y(n_225)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_138),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_221),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_241),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_170),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_210),
.B(n_150),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_223),
.B(n_229),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_226),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_164),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_228),
.A2(n_234),
.B1(n_238),
.B2(n_239),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_213),
.B(n_149),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_230),
.Y(n_255)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_177),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_233),
.B(n_242),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_180),
.A2(n_196),
.B1(n_204),
.B2(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_237),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_211),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_196),
.A2(n_181),
.B1(n_192),
.B2(n_208),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_181),
.A2(n_188),
.B1(n_193),
.B2(n_191),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_211),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_245),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_178),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_188),
.A2(n_211),
.B(n_184),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_243),
.A2(n_198),
.B(n_214),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_184),
.B1(n_182),
.B2(n_179),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_246),
.Y(n_263)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_203),
.B(n_200),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_223),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_200),
.B(n_209),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_250),
.A2(n_258),
.B(n_271),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_244),
.Y(n_252)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_252),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_216),
.A2(n_215),
.B1(n_185),
.B2(n_198),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_264),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_185),
.B1(n_214),
.B2(n_207),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_247),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_216),
.A2(n_207),
.B1(n_228),
.B2(n_220),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_267),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_221),
.A2(n_236),
.B1(n_231),
.B2(n_226),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_231),
.A2(n_224),
.B1(n_219),
.B2(n_222),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_235),
.A2(n_237),
.B(n_240),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_235),
.A2(n_239),
.B(n_234),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_275),
.B(n_258),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_235),
.A2(n_229),
.B1(n_227),
.B2(n_230),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_248),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g275 ( 
.A1(n_245),
.A2(n_246),
.B(n_232),
.Y(n_275)
);

NAND5xp2_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_217),
.C(n_241),
.D(n_264),
.E(n_259),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_276),
.A2(n_270),
.B1(n_286),
.B2(n_289),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_259),
.Y(n_277)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_265),
.C(n_267),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_285),
.C(n_263),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_250),
.B(n_273),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_282),
.A2(n_289),
.B(n_290),
.Y(n_309)
);

BUFx12_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_286),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_265),
.C(n_261),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_268),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_249),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_261),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_291),
.A2(n_295),
.B(n_256),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_251),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_292),
.A2(n_256),
.B1(n_270),
.B2(n_287),
.Y(n_311)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_297),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_260),
.B(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_255),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_288),
.B(n_274),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_313),
.C(n_284),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_253),
.B1(n_266),
.B2(n_252),
.Y(n_301)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_301),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_278),
.B(n_249),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_304),
.C(n_307),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_277),
.B(n_253),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_305),
.B(n_291),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_279),
.A2(n_263),
.B(n_257),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_310),
.B(n_308),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_284),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_312),
.A2(n_292),
.B1(n_293),
.B2(n_297),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_296),
.C(n_280),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_283),
.A2(n_280),
.B1(n_282),
.B2(n_276),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_279),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_281),
.A2(n_283),
.B1(n_295),
.B2(n_294),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_317),
.A2(n_315),
.B1(n_306),
.B2(n_314),
.Y(n_338)
);

BUFx12_ASAP7_75t_L g318 ( 
.A(n_298),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_326),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_290),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_320),
.B(n_323),
.Y(n_333)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_300),
.Y(n_321)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_321),
.Y(n_335)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_303),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_324),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_313),
.B(n_292),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_294),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_328),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_307),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_336),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_299),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_337),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_325),
.A2(n_312),
.B1(n_309),
.B2(n_310),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_340),
.A2(n_341),
.B1(n_324),
.B2(n_319),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_319),
.A2(n_309),
.B1(n_298),
.B2(n_311),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_332),
.B(n_321),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_348),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_343),
.Y(n_355)
);

AO21x2_ASAP7_75t_L g344 ( 
.A1(n_341),
.A2(n_316),
.B(n_328),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_346),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_339),
.A2(n_327),
.B(n_324),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_329),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_331),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_337),
.A2(n_329),
.B(n_318),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_349),
.B(n_340),
.Y(n_352)
);

OAI211xp5_ASAP7_75t_L g351 ( 
.A1(n_348),
.A2(n_335),
.B(n_334),
.C(n_338),
.Y(n_351)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_351),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_352),
.B(n_302),
.C(n_336),
.Y(n_356)
);

NOR2x1_ASAP7_75t_L g359 ( 
.A(n_354),
.B(n_344),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_356),
.B(n_358),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_355),
.B(n_345),
.C(n_334),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_359),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_357),
.C(n_353),
.Y(n_362)
);

BUFx24_ASAP7_75t_SL g363 ( 
.A(n_362),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_363),
.B(n_360),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_350),
.Y(n_365)
);


endmodule