module fake_jpeg_31563_n_421 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_421);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_421;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_52),
.Y(n_133)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_53),
.Y(n_118)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_13),
.C(n_20),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_56),
.B(n_48),
.C(n_45),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_65),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_66),
.B(n_40),
.Y(n_135)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_43),
.A2(n_12),
.B1(n_19),
.B2(n_18),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_69),
.A2(n_48),
.B1(n_31),
.B2(n_45),
.Y(n_120)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_83),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_87),
.Y(n_119)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_86),
.Y(n_96)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_89),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_93),
.B(n_109),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_111),
.B1(n_120),
.B2(n_131),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_80),
.A2(n_46),
.B1(n_47),
.B2(n_22),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_50),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_114),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_50),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_58),
.B(n_31),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_116),
.B(n_129),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_32),
.C(n_22),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_79),
.B(n_24),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_69),
.A2(n_47),
.B1(n_46),
.B2(n_32),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_23),
.Y(n_162)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_140),
.Y(n_182)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_62),
.B1(n_60),
.B2(n_51),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_142),
.A2(n_148),
.B1(n_105),
.B2(n_108),
.Y(n_189)
);

BUFx8_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

BUFx4f_ASAP7_75t_SL g195 ( 
.A(n_143),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_76),
.B1(n_81),
.B2(n_84),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_154),
.B1(n_166),
.B2(n_127),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_89),
.B1(n_87),
.B2(n_83),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_145),
.A2(n_107),
.B1(n_113),
.B2(n_156),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_96),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_150),
.Y(n_179)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_134),
.A2(n_52),
.B1(n_41),
.B2(n_26),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_23),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_82),
.B1(n_70),
.B2(n_71),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_161),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_99),
.A2(n_68),
.B(n_61),
.C(n_59),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_106),
.B(n_100),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_91),
.B(n_34),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_95),
.C(n_24),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_160),
.Y(n_172)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_164),
.Y(n_180)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_97),
.A2(n_57),
.B1(n_34),
.B2(n_26),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_103),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_170),
.Y(n_176)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

BUFx12_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_128),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_183),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_119),
.C(n_108),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_193),
.B1(n_139),
.B2(n_161),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_160),
.B1(n_169),
.B2(n_168),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_138),
.A2(n_110),
.B1(n_107),
.B2(n_127),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_190),
.A2(n_149),
.B1(n_170),
.B2(n_141),
.Y(n_205)
);

NAND2xp33_ASAP7_75t_SL g191 ( 
.A(n_159),
.B(n_133),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_197),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_105),
.C(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_200),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_162),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_202),
.Y(n_235)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_204),
.A2(n_172),
.B1(n_188),
.B2(n_101),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_207),
.B1(n_179),
.B2(n_180),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_153),
.B1(n_158),
.B2(n_136),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_165),
.B1(n_125),
.B2(n_147),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_179),
.B1(n_172),
.B2(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_150),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_213),
.Y(n_220)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_212),
.Y(n_240)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_176),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_170),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_214),
.B(n_216),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_215),
.A2(n_182),
.B(n_124),
.Y(n_224)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_218),
.B(n_196),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_219),
.A2(n_227),
.B1(n_204),
.B2(n_209),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_176),
.B(n_174),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_223),
.A2(n_238),
.B1(n_216),
.B2(n_212),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_200),
.B(n_181),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_231),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_208),
.B1(n_206),
.B2(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_232),
.Y(n_250)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_205),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_230),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_201),
.B(n_197),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_195),
.B(n_157),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_237),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_182),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_199),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_207),
.A2(n_118),
.B(n_124),
.Y(n_237)
);

INVx3_ASAP7_75t_SL g239 ( 
.A(n_211),
.Y(n_239)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_228),
.B(n_203),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_242),
.B(n_245),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_251),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_203),
.C(n_202),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_263),
.Y(n_284)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_252),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_259),
.B1(n_227),
.B2(n_223),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_171),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_254),
.B(n_256),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_192),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_225),
.B(n_234),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_219),
.A2(n_215),
.B1(n_218),
.B2(n_188),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_262),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_261),
.A2(n_239),
.B1(n_222),
.B2(n_188),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_217),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_192),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_250),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_278),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_251),
.B(n_226),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_274),
.B(n_281),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_L g275 ( 
.A1(n_241),
.A2(n_220),
.B(n_225),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_275),
.A2(n_178),
.B(n_143),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_276),
.A2(n_288),
.B1(n_264),
.B2(n_244),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_220),
.Y(n_277)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_243),
.B(n_221),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_243),
.A2(n_233),
.B(n_234),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_290),
.B(n_244),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_234),
.B(n_224),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_285),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g281 ( 
.A(n_263),
.B(n_238),
.CI(n_237),
.CON(n_281),
.SN(n_281)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_262),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_230),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_195),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_287),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_253),
.B1(n_265),
.B2(n_264),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_239),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_278),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_255),
.A2(n_239),
.B(n_195),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_309),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_255),
.C(n_261),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_297),
.C(n_302),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_296),
.A2(n_171),
.B(n_186),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_246),
.C(n_247),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_299),
.A2(n_310),
.B1(n_290),
.B2(n_281),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_269),
.A2(n_252),
.B1(n_260),
.B2(n_175),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_300),
.A2(n_271),
.B1(n_270),
.B2(n_268),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_301),
.B(n_303),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_173),
.C(n_163),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_282),
.B(n_195),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_314),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_164),
.C(n_155),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_186),
.C(n_171),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_283),
.Y(n_308)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_282),
.B(n_178),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_288),
.A2(n_175),
.B1(n_118),
.B2(n_132),
.Y(n_310)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_283),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_313),
.A2(n_304),
.B1(n_307),
.B2(n_299),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_178),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_178),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_186),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_186),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_280),
.Y(n_322)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_319),
.Y(n_348)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_321),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_322),
.B(n_329),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_306),
.A2(n_268),
.B1(n_270),
.B2(n_281),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_333),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_324),
.A2(n_315),
.B1(n_297),
.B2(n_314),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_294),
.B(n_267),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_339),
.Y(n_354)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_303),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_327),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_293),
.A2(n_140),
.B(n_151),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_328),
.A2(n_171),
.B(n_109),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_312),
.B(n_143),
.Y(n_329)
);

NAND2x1p5_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_175),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_330),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_306),
.A2(n_14),
.B1(n_21),
.B2(n_18),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_41),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_335),
.A2(n_41),
.B(n_109),
.Y(n_347)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_338),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_335),
.A2(n_304),
.B(n_316),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_340),
.A2(n_346),
.B(n_325),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_352),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_317),
.A2(n_310),
.B1(n_305),
.B2(n_301),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_342),
.A2(n_318),
.B1(n_339),
.B2(n_337),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_291),
.C(n_302),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_332),
.C(n_326),
.Y(n_358)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_345),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_331),
.B(n_291),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_334),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_324),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_353),
.A2(n_322),
.B1(n_330),
.B2(n_329),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_360),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_366),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_364),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_325),
.C(n_337),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_371),
.C(n_357),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_341),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_354),
.A2(n_12),
.B(n_21),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_367),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_12),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_369),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_356),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_355),
.A2(n_41),
.B1(n_10),
.B2(n_13),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_370),
.B(n_371),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_10),
.C(n_17),
.Y(n_371)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_372),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_368),
.Y(n_373)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_373),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_358),
.B(n_349),
.Y(n_378)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_378),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_351),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_380),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_361),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_383),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_9),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_363),
.A2(n_355),
.B1(n_348),
.B2(n_350),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_375),
.A2(n_343),
.B1(n_340),
.B2(n_347),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_395),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_361),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

OAI322xp33_ASAP7_75t_L g387 ( 
.A1(n_377),
.A2(n_343),
.A3(n_365),
.B1(n_359),
.B2(n_352),
.C1(n_345),
.C2(n_7),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_387),
.A2(n_10),
.B(n_16),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_379),
.A2(n_376),
.B1(n_382),
.B2(n_374),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_390),
.A2(n_4),
.B1(n_15),
.B2(n_14),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_376),
.B(n_9),
.C(n_16),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_391),
.B(n_392),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_379),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_396),
.B(n_399),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_7),
.C(n_16),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_401),
.B(n_391),
.C(n_389),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_394),
.A2(n_13),
.B(n_15),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_402),
.A2(n_404),
.B(n_2),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_21),
.Y(n_403)
);

AOI21x1_ASAP7_75t_L g408 ( 
.A1(n_403),
.A2(n_0),
.B(n_1),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_392),
.A2(n_0),
.B(n_1),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_405),
.B(n_406),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_397),
.A2(n_388),
.B(n_386),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_398),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_407),
.B(n_400),
.C(n_2),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_408),
.B(n_410),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_409),
.B(n_400),
.C(n_390),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_412),
.B(n_414),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_413),
.A2(n_2),
.B(n_3),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_411),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_417),
.Y(n_418)
);

AOI31xp33_ASAP7_75t_L g419 ( 
.A1(n_418),
.A2(n_415),
.A3(n_2),
.B(n_3),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_419),
.B(n_3),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_3),
.Y(n_421)
);


endmodule