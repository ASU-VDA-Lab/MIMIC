module fake_netlist_6_3940_n_1501 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_364, n_295, n_190, n_262, n_187, n_60, n_361, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1501);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_364;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1501;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_474;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_482;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_1485;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1109;
wire n_712;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_359),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_157),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_47),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_336),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_45),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_280),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_25),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_22),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_321),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_169),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_155),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_46),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_273),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_367),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_43),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_112),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_156),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_101),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_140),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_147),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_26),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_84),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_44),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_72),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_115),
.Y(n_400)
);

BUFx10_ASAP7_75t_L g401 ( 
.A(n_259),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_341),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_22),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_122),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_364),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_286),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_355),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_10),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_258),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_288),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_357),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_97),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_141),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_236),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_76),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_89),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_130),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_348),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_354),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_209),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_195),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_14),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_271),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_325),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_228),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_216),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_87),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_92),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_289),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_137),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_340),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_302),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_366),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_106),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_60),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_349),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_48),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_90),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_215),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_210),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_23),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_265),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_117),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_368),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_345),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_212),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_12),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_230),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_243),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_170),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_172),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_34),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_16),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_65),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_320),
.Y(n_455)
);

BUFx2_ASAP7_75t_SL g456 ( 
.A(n_295),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_214),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_298),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_343),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_213),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_77),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_177),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_337),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_200),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_6),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_282),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_217),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_370),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_105),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_208),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_143),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_38),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_103),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_218),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_191),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_316),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_352),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_347),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_31),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_221),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_306),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_31),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_241),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_127),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_26),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_91),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_138),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_344),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_300),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_121),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_81),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_176),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_88),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_240),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_123),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_168),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_330),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_196),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_279),
.Y(n_499)
);

BUFx10_ASAP7_75t_L g500 ( 
.A(n_175),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_296),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_292),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_171),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_272),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_183),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_267),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_75),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_128),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_33),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_119),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_95),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_59),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_247),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_53),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_185),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_23),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_64),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_192),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_249),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_275),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_244),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_318),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_80),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_238),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_24),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_41),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_67),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_255),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_308),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_219),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_7),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_62),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_118),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_231),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_113),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_69),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_201),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_339),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_233),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_199),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_52),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_73),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_229),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_148),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_299),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_328),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_159),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_124),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_125),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_180),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_309),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_203),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_224),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_40),
.Y(n_554)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_74),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_290),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_338),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_361),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_20),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_17),
.Y(n_560)
);

BUFx10_ASAP7_75t_L g561 ( 
.A(n_285),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_114),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_7),
.Y(n_563)
);

NOR2xp67_ASAP7_75t_L g564 ( 
.A(n_144),
.B(n_274),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_79),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_346),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_401),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_381),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_381),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_381),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_401),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_381),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_405),
.B(n_0),
.Y(n_573)
);

BUFx12f_ASAP7_75t_L g574 ( 
.A(n_500),
.Y(n_574)
);

OA22x2_ASAP7_75t_L g575 ( 
.A1(n_396),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_575)
);

BUFx12f_ASAP7_75t_L g576 ( 
.A(n_500),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_403),
.Y(n_577)
);

BUFx8_ASAP7_75t_SL g578 ( 
.A(n_422),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_479),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_519),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_379),
.Y(n_581)
);

BUFx8_ASAP7_75t_SL g582 ( 
.A(n_527),
.Y(n_582)
);

BUFx12f_ASAP7_75t_L g583 ( 
.A(n_519),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_501),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_465),
.Y(n_585)
);

BUFx8_ASAP7_75t_SL g586 ( 
.A(n_388),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_560),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_528),
.B(n_1),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_472),
.Y(n_589)
);

BUFx12f_ASAP7_75t_L g590 ( 
.A(n_561),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_525),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_559),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_561),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_501),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_409),
.B(n_2),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_409),
.B(n_3),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_432),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_542),
.B(n_3),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_394),
.B(n_4),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_432),
.B(n_4),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_501),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_533),
.B(n_5),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_533),
.B(n_5),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_382),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_501),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_394),
.B(n_6),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_413),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_413),
.B(n_8),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_376),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_434),
.B(n_9),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_434),
.B(n_11),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_450),
.A2(n_49),
.B(n_42),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_408),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_436),
.B(n_11),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_378),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_436),
.B(n_12),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_442),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_383),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_386),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_442),
.B(n_13),
.Y(n_620)
);

BUFx8_ASAP7_75t_SL g621 ( 
.A(n_466),
.Y(n_621)
);

INVx6_ASAP7_75t_L g622 ( 
.A(n_392),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_441),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_395),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_447),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_513),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_398),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_406),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_452),
.Y(n_629)
);

BUFx8_ASAP7_75t_L g630 ( 
.A(n_513),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_549),
.B(n_13),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_486),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_375),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_549),
.B(n_14),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_453),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_412),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_414),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_482),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_377),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_417),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_471),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_489),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_418),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_421),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_485),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_380),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_509),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_384),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_427),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_438),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_440),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_423),
.B(n_555),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_443),
.Y(n_653)
);

BUFx12f_ASAP7_75t_L g654 ( 
.A(n_516),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_446),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_451),
.Y(n_656)
);

BUFx8_ASAP7_75t_L g657 ( 
.A(n_454),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_526),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_531),
.Y(n_659)
);

BUFx12f_ASAP7_75t_L g660 ( 
.A(n_554),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_457),
.B(n_15),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_463),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_563),
.B(n_18),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_469),
.A2(n_51),
.B(n_50),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_473),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_480),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_487),
.B(n_18),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_568),
.Y(n_668)
);

BUFx10_ASAP7_75t_L g669 ( 
.A(n_622),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_581),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_586),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_569),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_570),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_621),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_572),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_639),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_646),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_578),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_607),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_632),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_582),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_633),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_607),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_607),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_626),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_648),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_567),
.Y(n_687)
);

BUFx10_ASAP7_75t_L g688 ( 
.A(n_622),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_626),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_626),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_615),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_574),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_576),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_583),
.Y(n_694)
);

AOI21x1_ASAP7_75t_L g695 ( 
.A1(n_617),
.A2(n_511),
.B(n_494),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_590),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_654),
.Y(n_697)
);

INVxp33_ASAP7_75t_SL g698 ( 
.A(n_625),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_R g699 ( 
.A(n_613),
.B(n_496),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_584),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_660),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_604),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_645),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_584),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_618),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_584),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_601),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_587),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_571),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_652),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_580),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_593),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_635),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_624),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_647),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_627),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_R g717 ( 
.A(n_613),
.B(n_529),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_SL g718 ( 
.A1(n_573),
.A2(n_598),
.B1(n_588),
.B2(n_609),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_601),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_657),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_663),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_637),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_657),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_601),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_623),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_623),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_605),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_643),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_R g729 ( 
.A(n_629),
.B(n_385),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_629),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_630),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_575),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_638),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_638),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_605),
.Y(n_735)
);

NOR2xp67_ASAP7_75t_L g736 ( 
.A(n_659),
.B(n_514),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_659),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_630),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_595),
.B(n_505),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_597),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_665),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_619),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_SL g743 ( 
.A1(n_658),
.A2(n_538),
.B1(n_565),
.B2(n_545),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_661),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_641),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_605),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_628),
.B(n_506),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_641),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_641),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_642),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_642),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_642),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_606),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_699),
.B(n_596),
.Y(n_754)
);

OAI21xp33_ASAP7_75t_L g755 ( 
.A1(n_739),
.A2(n_631),
.B(n_599),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_739),
.B(n_594),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_717),
.B(n_596),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_750),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_679),
.B(n_594),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_725),
.B(n_667),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_700),
.Y(n_761)
);

OA21x2_ASAP7_75t_L g762 ( 
.A1(n_695),
.A2(n_664),
.B(n_612),
.Y(n_762)
);

NAND2xp33_ASAP7_75t_L g763 ( 
.A(n_726),
.B(n_730),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_733),
.B(n_600),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_734),
.B(n_600),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_704),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_683),
.B(n_684),
.Y(n_767)
);

BUFx6f_ASAP7_75t_SL g768 ( 
.A(n_669),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_685),
.B(n_689),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_737),
.B(n_602),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_690),
.B(n_736),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_713),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_707),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_719),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_742),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_698),
.B(n_602),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_753),
.B(n_594),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_724),
.Y(n_778)
);

OR2x2_ASAP7_75t_SL g779 ( 
.A(n_713),
.B(n_611),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_727),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_753),
.B(n_603),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_735),
.B(n_603),
.Y(n_782)
);

AO221x1_ASAP7_75t_L g783 ( 
.A1(n_743),
.A2(n_522),
.B1(n_535),
.B2(n_524),
.C(n_521),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_751),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_715),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_746),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_751),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_745),
.B(n_606),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_721),
.B(n_636),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_702),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_721),
.B(n_614),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_751),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_749),
.B(n_640),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_751),
.Y(n_794)
);

AO221x1_ASAP7_75t_L g795 ( 
.A1(n_718),
.A2(n_543),
.B1(n_556),
.B2(n_548),
.C(n_541),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_748),
.Y(n_796)
);

AND2x6_ASAP7_75t_SL g797 ( 
.A(n_708),
.B(n_620),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_752),
.B(n_740),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_747),
.B(n_608),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_706),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_676),
.B(n_634),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_672),
.B(n_640),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_677),
.B(n_608),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_709),
.B(n_610),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_706),
.B(n_644),
.Y(n_805)
);

INVx3_ASAP7_75t_R g806 ( 
.A(n_687),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_706),
.B(n_644),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_691),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_711),
.B(n_610),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_706),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_L g811 ( 
.A(n_732),
.B(n_550),
.C(n_577),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_L g812 ( 
.A(n_732),
.B(n_387),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_705),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_686),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_714),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_712),
.B(n_649),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_703),
.B(n_649),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_668),
.B(n_650),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_716),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_L g820 ( 
.A(n_729),
.B(n_616),
.C(n_592),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_744),
.B(n_616),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_673),
.B(n_650),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_669),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_L g824 ( 
.A(n_722),
.B(n_653),
.C(n_651),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_710),
.B(n_651),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_682),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_675),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_728),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_688),
.B(n_738),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_741),
.B(n_653),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_688),
.Y(n_831)
);

NOR2xp67_ASAP7_75t_L g832 ( 
.A(n_697),
.B(n_617),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_701),
.B(n_389),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_692),
.B(n_655),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_693),
.B(n_655),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_694),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_696),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_720),
.B(n_656),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_723),
.B(n_656),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_670),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_731),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_L g842 ( 
.A(n_671),
.B(n_579),
.C(n_662),
.Y(n_842)
);

NOR2xp67_ASAP7_75t_L g843 ( 
.A(n_674),
.B(n_390),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_680),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_755),
.A2(n_564),
.B1(n_558),
.B2(n_562),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_791),
.A2(n_393),
.B1(n_397),
.B2(n_391),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_816),
.B(n_591),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_760),
.B(n_801),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_828),
.Y(n_849)
);

BUFx12f_ASAP7_75t_L g850 ( 
.A(n_823),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_765),
.B(n_662),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_770),
.B(n_662),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_796),
.B(n_585),
.Y(n_853)
);

NOR2x2_ASAP7_75t_L g854 ( 
.A(n_797),
.B(n_678),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_840),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_776),
.B(n_681),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_775),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_808),
.Y(n_858)
);

OAI22xp33_ASAP7_75t_L g859 ( 
.A1(n_820),
.A2(n_400),
.B1(n_402),
.B2(n_399),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_813),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_827),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_814),
.Y(n_862)
);

BUFx6f_ASAP7_75t_SL g863 ( 
.A(n_826),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_756),
.B(n_666),
.Y(n_864)
);

BUFx4f_ASAP7_75t_L g865 ( 
.A(n_814),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_825),
.B(n_404),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_819),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_758),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_755),
.A2(n_812),
.B1(n_757),
.B2(n_754),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_761),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_768),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_805),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_817),
.B(n_407),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_766),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_807),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_789),
.A2(n_411),
.B(n_415),
.C(n_410),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_772),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_803),
.B(n_416),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_782),
.A2(n_420),
.B(n_419),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_799),
.A2(n_425),
.B1(n_426),
.B2(n_424),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_781),
.B(n_666),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_768),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_815),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_767),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_773),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_774),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_769),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_793),
.B(n_666),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_777),
.B(n_428),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_821),
.B(n_589),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_788),
.A2(n_430),
.B(n_429),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_795),
.A2(n_456),
.B1(n_433),
.B2(n_435),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_798),
.B(n_431),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_SL g894 ( 
.A(n_811),
.B(n_439),
.C(n_437),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_778),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_780),
.Y(n_896)
);

BUFx8_ASAP7_75t_SL g897 ( 
.A(n_814),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_844),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_764),
.A2(n_445),
.B1(n_448),
.B2(n_444),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_784),
.Y(n_900)
);

BUFx12f_ASAP7_75t_SL g901 ( 
.A(n_806),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_804),
.A2(n_455),
.B1(n_458),
.B2(n_449),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_838),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_784),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_784),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_787),
.B(n_459),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_792),
.B(n_460),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_790),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_786),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_800),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_809),
.A2(n_462),
.B1(n_464),
.B2(n_461),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_783),
.A2(n_468),
.B1(n_470),
.B2(n_467),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_810),
.B(n_474),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_830),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_771),
.B(n_475),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_794),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_839),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_794),
.B(n_476),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_802),
.Y(n_919)
);

AND2x6_ASAP7_75t_L g920 ( 
.A(n_831),
.B(n_585),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_794),
.B(n_477),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_818),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_832),
.B(n_478),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_779),
.A2(n_483),
.B1(n_484),
.B2(n_481),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_785),
.B(n_589),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_832),
.B(n_488),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_762),
.A2(n_491),
.B1(n_492),
.B2(n_490),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_834),
.B(n_493),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_822),
.Y(n_929)
);

AND3x1_ASAP7_75t_L g930 ( 
.A(n_835),
.B(n_19),
.C(n_20),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_797),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_763),
.B(n_495),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_833),
.B(n_497),
.Y(n_933)
);

NAND2x2_ASAP7_75t_L g934 ( 
.A(n_836),
.B(n_19),
.Y(n_934)
);

OAI21xp33_ASAP7_75t_L g935 ( 
.A1(n_842),
.A2(n_499),
.B(n_498),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_L g936 ( 
.A(n_759),
.B(n_502),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_837),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_843),
.Y(n_938)
);

NAND3xp33_ASAP7_75t_L g939 ( 
.A(n_843),
.B(n_504),
.C(n_503),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_841),
.B(n_21),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_762),
.B(n_507),
.Y(n_941)
);

OR2x2_ASAP7_75t_SL g942 ( 
.A(n_824),
.B(n_21),
.Y(n_942)
);

AND2x6_ASAP7_75t_SL g943 ( 
.A(n_829),
.B(n_24),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_865),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_941),
.A2(n_824),
.B(n_510),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_897),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_848),
.B(n_508),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_876),
.A2(n_515),
.B(n_517),
.C(n_512),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_853),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_865),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_869),
.A2(n_520),
.B(n_523),
.C(n_518),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_853),
.Y(n_952)
);

BUFx8_ASAP7_75t_L g953 ( 
.A(n_863),
.Y(n_953)
);

O2A1O1Ixp5_ASAP7_75t_L g954 ( 
.A1(n_864),
.A2(n_532),
.B(n_534),
.C(n_530),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_881),
.A2(n_875),
.B(n_872),
.Y(n_955)
);

CKINVDCx14_ASAP7_75t_R g956 ( 
.A(n_901),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_877),
.Y(n_957)
);

AOI33xp33_ASAP7_75t_L g958 ( 
.A1(n_845),
.A2(n_25),
.A3(n_27),
.B1(n_28),
.B2(n_29),
.B3(n_30),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_866),
.A2(n_537),
.B1(n_539),
.B2(n_536),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_862),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_SL g961 ( 
.A1(n_845),
.A2(n_544),
.B(n_546),
.C(n_540),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_862),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_919),
.A2(n_551),
.B(n_547),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_857),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_910),
.A2(n_55),
.B(n_54),
.Y(n_965)
);

NAND2xp33_ASAP7_75t_R g966 ( 
.A(n_937),
.B(n_552),
.Y(n_966)
);

AOI21x1_ASAP7_75t_L g967 ( 
.A1(n_906),
.A2(n_557),
.B(n_553),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_900),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_858),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_903),
.B(n_566),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_917),
.B(n_27),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_868),
.Y(n_972)
);

O2A1O1Ixp5_ASAP7_75t_L g973 ( 
.A1(n_873),
.A2(n_223),
.B(n_373),
.C(n_372),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_893),
.B(n_28),
.Y(n_974)
);

OA22x2_ASAP7_75t_L g975 ( 
.A1(n_931),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_870),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_SL g977 ( 
.A(n_908),
.B(n_56),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_SL g978 ( 
.A1(n_892),
.A2(n_933),
.B(n_922),
.C(n_929),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_856),
.B(n_32),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_913),
.A2(n_888),
.B(n_914),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_884),
.B(n_33),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_883),
.B(n_34),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_907),
.A2(n_58),
.B(n_57),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_926),
.B(n_61),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_887),
.A2(n_860),
.B1(n_847),
.B2(n_867),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_927),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_859),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_925),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_R g989 ( 
.A(n_855),
.B(n_63),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_918),
.A2(n_68),
.B(n_66),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_863),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_912),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_909),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_921),
.A2(n_71),
.B(n_70),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_851),
.B(n_78),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_SL g996 ( 
.A1(n_849),
.A2(n_245),
.B(n_371),
.C(n_82),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_898),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_852),
.A2(n_39),
.B(n_41),
.C(n_83),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_938),
.A2(n_85),
.B1(n_86),
.B2(n_93),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_SL g1000 ( 
.A(n_899),
.B(n_94),
.C(n_96),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_896),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_846),
.B(n_98),
.Y(n_1002)
);

NOR2x1_ASAP7_75t_SL g1003 ( 
.A(n_904),
.B(n_99),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_890),
.B(n_100),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_889),
.A2(n_102),
.B(n_104),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_915),
.B(n_107),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_861),
.B(n_108),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_923),
.A2(n_109),
.B(n_110),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_932),
.A2(n_111),
.B1(n_116),
.B2(n_120),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_924),
.B(n_126),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_885),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_SL g1012 ( 
.A(n_871),
.B(n_129),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_895),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_910),
.A2(n_131),
.B(n_132),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_940),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_879),
.A2(n_133),
.B(n_134),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_L g1017 ( 
.A(n_894),
.B(n_135),
.C(n_136),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_874),
.B(n_139),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_SL g1019 ( 
.A(n_882),
.B(n_142),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_SL g1020 ( 
.A(n_979),
.B(n_850),
.Y(n_1020)
);

INVx6_ASAP7_75t_SL g1021 ( 
.A(n_956),
.Y(n_1021)
);

BUFx8_ASAP7_75t_L g1022 ( 
.A(n_946),
.Y(n_1022)
);

BUFx5_ASAP7_75t_L g1023 ( 
.A(n_964),
.Y(n_1023)
);

BUFx2_ASAP7_75t_SL g1024 ( 
.A(n_944),
.Y(n_1024)
);

INVx6_ASAP7_75t_L g1025 ( 
.A(n_944),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_962),
.Y(n_1026)
);

AO21x2_ASAP7_75t_L g1027 ( 
.A1(n_945),
.A2(n_928),
.B(n_878),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_953),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_953),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_944),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_969),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_972),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_993),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1001),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_965),
.A2(n_916),
.B(n_905),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_950),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_SL g1037 ( 
.A1(n_1003),
.A2(n_891),
.B(n_902),
.Y(n_1037)
);

INVx8_ASAP7_75t_L g1038 ( 
.A(n_950),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_950),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_955),
.A2(n_939),
.B(n_880),
.Y(n_1040)
);

BUFx12f_ASAP7_75t_L g1041 ( 
.A(n_991),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_997),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1011),
.Y(n_1043)
);

AO21x2_ASAP7_75t_L g1044 ( 
.A1(n_980),
.A2(n_935),
.B(n_936),
.Y(n_1044)
);

INVx5_ASAP7_75t_L g1045 ( 
.A(n_962),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_962),
.B(n_874),
.Y(n_1046)
);

AO21x2_ASAP7_75t_L g1047 ( 
.A1(n_1016),
.A2(n_911),
.B(n_920),
.Y(n_1047)
);

AO21x2_ASAP7_75t_L g1048 ( 
.A1(n_951),
.A2(n_920),
.B(n_886),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_960),
.B(n_886),
.Y(n_1049)
);

OR2x6_ASAP7_75t_L g1050 ( 
.A(n_957),
.B(n_854),
.Y(n_1050)
);

AOI22x1_ASAP7_75t_L g1051 ( 
.A1(n_1004),
.A2(n_920),
.B1(n_934),
.B2(n_942),
.Y(n_1051)
);

INVx8_ASAP7_75t_L g1052 ( 
.A(n_968),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_976),
.Y(n_1053)
);

OA21x2_ASAP7_75t_L g1054 ( 
.A1(n_1014),
.A2(n_973),
.B(n_954),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_947),
.B(n_920),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1013),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_968),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_968),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_988),
.Y(n_1059)
);

AO21x2_ASAP7_75t_L g1060 ( 
.A1(n_1006),
.A2(n_930),
.B(n_145),
.Y(n_1060)
);

AOI22x1_ASAP7_75t_L g1061 ( 
.A1(n_1005),
.A2(n_943),
.B1(n_149),
.B2(n_150),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_949),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_952),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_1018),
.A2(n_146),
.B(n_151),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_1007),
.A2(n_152),
.B(n_153),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_989),
.Y(n_1066)
);

BUFx12f_ASAP7_75t_L g1067 ( 
.A(n_1012),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_985),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_967),
.A2(n_154),
.B(n_158),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_981),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_982),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_1015),
.B(n_984),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_1010),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_958),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_975),
.Y(n_1075)
);

NAND2x1_ASAP7_75t_L g1076 ( 
.A(n_983),
.B(n_160),
.Y(n_1076)
);

INVxp67_ASAP7_75t_SL g1077 ( 
.A(n_971),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_970),
.B(n_161),
.Y(n_1078)
);

AO21x2_ASAP7_75t_L g1079 ( 
.A1(n_978),
.A2(n_995),
.B(n_974),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_977),
.Y(n_1080)
);

BUFx12f_ASAP7_75t_L g1081 ( 
.A(n_1019),
.Y(n_1081)
);

INVx4_ASAP7_75t_L g1082 ( 
.A(n_966),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_1042),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1031),
.Y(n_1084)
);

AOI21x1_ASAP7_75t_L g1085 ( 
.A1(n_1055),
.A2(n_994),
.B(n_990),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_1045),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1033),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1034),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_1059),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1043),
.Y(n_1090)
);

NAND2x1p5_ASAP7_75t_L g1091 ( 
.A(n_1045),
.B(n_1002),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_1022),
.Y(n_1092)
);

OA21x2_ASAP7_75t_L g1093 ( 
.A1(n_1035),
.A2(n_986),
.B(n_998),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_1059),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1032),
.Y(n_1095)
);

OR2x6_ASAP7_75t_L g1096 ( 
.A(n_1038),
.B(n_987),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1056),
.Y(n_1097)
);

BUFx2_ASAP7_75t_R g1098 ( 
.A(n_1028),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1053),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1073),
.A2(n_992),
.B1(n_1017),
.B2(n_1000),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_1045),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1064),
.A2(n_1008),
.B(n_948),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1071),
.B(n_963),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1068),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_SL g1105 ( 
.A1(n_1073),
.A2(n_999),
.B1(n_1009),
.B2(n_959),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1021),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_1022),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1023),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1061),
.A2(n_961),
.B1(n_996),
.B2(n_164),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1080),
.A2(n_1082),
.B1(n_1072),
.B2(n_1066),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_1041),
.Y(n_1111)
);

AO21x1_ASAP7_75t_SL g1112 ( 
.A1(n_1055),
.A2(n_162),
.B(n_163),
.Y(n_1112)
);

AOI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1054),
.A2(n_165),
.B(n_166),
.Y(n_1113)
);

OAI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_1020),
.A2(n_1077),
.B1(n_1080),
.B2(n_1082),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1063),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1072),
.A2(n_1066),
.B1(n_1078),
.B2(n_1081),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1023),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1023),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1077),
.B(n_167),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1075),
.B(n_173),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1023),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1023),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1062),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1045),
.Y(n_1124)
);

BUFx8_ASAP7_75t_L g1125 ( 
.A(n_1029),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1074),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1038),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1070),
.Y(n_1128)
);

INVxp67_ASAP7_75t_SL g1129 ( 
.A(n_1057),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_1038),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_SL g1131 ( 
.A1(n_1067),
.A2(n_174),
.B1(n_178),
.B2(n_179),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1070),
.Y(n_1132)
);

AO21x1_ASAP7_75t_L g1133 ( 
.A1(n_1040),
.A2(n_1076),
.B(n_1069),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1058),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_1021),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_1030),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_SL g1137 ( 
.A1(n_1050),
.A2(n_181),
.B1(n_182),
.B2(n_184),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1030),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1036),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1075),
.B(n_186),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1058),
.Y(n_1141)
);

BUFx12f_ASAP7_75t_L g1142 ( 
.A(n_1050),
.Y(n_1142)
);

CKINVDCx11_ASAP7_75t_R g1143 ( 
.A(n_1050),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1057),
.Y(n_1144)
);

NAND2xp33_ASAP7_75t_R g1145 ( 
.A(n_1106),
.B(n_1054),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1110),
.B(n_1036),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_L g1147 ( 
.A(n_1100),
.B(n_1020),
.C(n_1051),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1106),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1100),
.A2(n_1060),
.B1(n_1047),
.B2(n_1079),
.Y(n_1149)
);

NOR2x1_ASAP7_75t_SL g1150 ( 
.A(n_1112),
.B(n_1048),
.Y(n_1150)
);

AND2x2_ASAP7_75t_SL g1151 ( 
.A(n_1119),
.B(n_1026),
.Y(n_1151)
);

NAND2xp33_ASAP7_75t_R g1152 ( 
.A(n_1135),
.B(n_1040),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1084),
.Y(n_1153)
);

INVxp67_ASAP7_75t_L g1154 ( 
.A(n_1094),
.Y(n_1154)
);

CKINVDCx16_ASAP7_75t_R g1155 ( 
.A(n_1092),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1104),
.Y(n_1156)
);

AND2x2_ASAP7_75t_SL g1157 ( 
.A(n_1119),
.B(n_1026),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1125),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1105),
.A2(n_1065),
.B(n_1024),
.C(n_1039),
.Y(n_1159)
);

OAI222xp33_ASAP7_75t_L g1160 ( 
.A1(n_1131),
.A2(n_1046),
.B1(n_1049),
.B2(n_1060),
.C1(n_1047),
.C2(n_1079),
.Y(n_1160)
);

BUFx4f_ASAP7_75t_SL g1161 ( 
.A(n_1125),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1090),
.Y(n_1162)
);

NAND2xp33_ASAP7_75t_SL g1163 ( 
.A(n_1130),
.B(n_1136),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1087),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1098),
.Y(n_1165)
);

OR2x6_ASAP7_75t_L g1166 ( 
.A(n_1130),
.B(n_1052),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1103),
.B(n_1025),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1127),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1127),
.B(n_1027),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1136),
.B(n_1027),
.Y(n_1170)
);

CKINVDCx16_ASAP7_75t_R g1171 ( 
.A(n_1107),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1089),
.B(n_1025),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1089),
.B(n_1128),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1088),
.Y(n_1174)
);

NAND2xp33_ASAP7_75t_R g1175 ( 
.A(n_1083),
.B(n_1025),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_1133),
.A2(n_1048),
.A3(n_1044),
.B(n_1037),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1098),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1086),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_SL g1179 ( 
.A1(n_1140),
.A2(n_1052),
.B(n_1046),
.C(n_1049),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_SL g1180 ( 
.A(n_1116),
.B(n_1052),
.C(n_1044),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1132),
.B(n_187),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_1094),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1138),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1120),
.B(n_188),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_SL g1185 ( 
.A1(n_1140),
.A2(n_189),
.B(n_190),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1095),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1136),
.Y(n_1187)
);

OR2x6_ASAP7_75t_L g1188 ( 
.A(n_1096),
.B(n_193),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_1123),
.B(n_194),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1139),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1144),
.B(n_197),
.Y(n_1191)
);

NAND2xp33_ASAP7_75t_SL g1192 ( 
.A(n_1139),
.B(n_198),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1099),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1139),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1097),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1115),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1111),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1126),
.B(n_374),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1142),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_R g1200 ( 
.A(n_1086),
.B(n_202),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_R g1201 ( 
.A(n_1143),
.B(n_204),
.Y(n_1201)
);

CKINVDCx16_ASAP7_75t_R g1202 ( 
.A(n_1137),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1134),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1143),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1108),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1105),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1114),
.B(n_369),
.Y(n_1207)
);

CKINVDCx16_ASAP7_75t_R g1208 ( 
.A(n_1096),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1114),
.B(n_211),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1096),
.A2(n_220),
.B1(n_222),
.B2(n_225),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1131),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1141),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1124),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1129),
.B(n_226),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1129),
.B(n_227),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1117),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1173),
.B(n_1091),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1211),
.A2(n_1091),
.B1(n_1109),
.B2(n_1118),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1167),
.B(n_1101),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1182),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1169),
.B(n_1121),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1156),
.Y(n_1222)
);

INVxp67_ASAP7_75t_SL g1223 ( 
.A(n_1154),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1164),
.B(n_1122),
.Y(n_1224)
);

NOR2x1p5_ASAP7_75t_L g1225 ( 
.A(n_1147),
.B(n_1113),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1183),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1156),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1195),
.Y(n_1228)
);

AOI211xp5_ASAP7_75t_L g1229 ( 
.A1(n_1207),
.A2(n_1209),
.B(n_1201),
.C(n_1160),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1164),
.Y(n_1230)
);

BUFx12f_ASAP7_75t_L g1231 ( 
.A(n_1158),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1194),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1174),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1169),
.B(n_1101),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1196),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1170),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1174),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1205),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1205),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1170),
.B(n_1153),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1151),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1162),
.B(n_1093),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1206),
.A2(n_1109),
.B1(n_1093),
.B2(n_1102),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1203),
.B(n_1085),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1190),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1202),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1216),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1212),
.B(n_365),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1190),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1193),
.B(n_237),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1186),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1176),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1146),
.B(n_363),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1176),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1208),
.B(n_239),
.Y(n_1255)
);

INVx4_ASAP7_75t_L g1256 ( 
.A(n_1188),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_1172),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1149),
.B(n_362),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1157),
.B(n_242),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1213),
.Y(n_1260)
);

OAI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1188),
.A2(n_246),
.B1(n_248),
.B2(n_250),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1176),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1150),
.B(n_251),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1215),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1150),
.Y(n_1265)
);

BUFx12f_ASAP7_75t_L g1266 ( 
.A(n_1204),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1187),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1180),
.B(n_360),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1178),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1178),
.B(n_252),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1181),
.B(n_358),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1189),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1198),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1185),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1191),
.B(n_253),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1184),
.B(n_356),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1214),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1190),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1179),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1210),
.A2(n_1192),
.B1(n_1199),
.B2(n_1148),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1159),
.B(n_1168),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1168),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1229),
.B(n_1273),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1230),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1233),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1257),
.B(n_1155),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1226),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1267),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1236),
.B(n_1171),
.Y(n_1289)
);

OA21x2_ASAP7_75t_L g1290 ( 
.A1(n_1262),
.A2(n_1145),
.B(n_1152),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1222),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1222),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1268),
.B(n_1175),
.C(n_1163),
.Y(n_1293)
);

AND2x4_ASAP7_75t_SL g1294 ( 
.A(n_1256),
.B(n_1168),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1236),
.B(n_1197),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1227),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1249),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1280),
.A2(n_1200),
.B(n_1161),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1227),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1237),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1240),
.B(n_1165),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1237),
.B(n_1166),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1244),
.Y(n_1303)
);

AND2x4_ASAP7_75t_SL g1304 ( 
.A(n_1256),
.B(n_1234),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1238),
.Y(n_1305)
);

INVxp33_ASAP7_75t_L g1306 ( 
.A(n_1219),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1240),
.B(n_1177),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1238),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1239),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1241),
.B(n_1166),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1241),
.B(n_254),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1239),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1217),
.B(n_353),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1228),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1235),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1244),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1265),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1242),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1224),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1232),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1224),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1264),
.B(n_256),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1223),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1234),
.B(n_351),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1256),
.B(n_1277),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1234),
.B(n_257),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1277),
.B(n_1272),
.Y(n_1327)
);

NOR3xp33_ASAP7_75t_L g1328 ( 
.A(n_1261),
.B(n_260),
.C(n_261),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1273),
.B(n_262),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1251),
.B(n_1220),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1253),
.B(n_263),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1242),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1253),
.B(n_350),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1305),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1305),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1284),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1287),
.B(n_1255),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1303),
.B(n_1262),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1303),
.B(n_1265),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1288),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1316),
.B(n_1252),
.Y(n_1341)
);

AND2x2_ASAP7_75t_SL g1342 ( 
.A(n_1290),
.B(n_1281),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1285),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1308),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1291),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1318),
.B(n_1252),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1318),
.B(n_1254),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1316),
.B(n_1254),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1320),
.B(n_1255),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1317),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1314),
.B(n_1268),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1306),
.B(n_1323),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1317),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1308),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1306),
.B(n_1221),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1332),
.B(n_1221),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1295),
.B(n_1221),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1292),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1283),
.B(n_1293),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1315),
.B(n_1247),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1296),
.Y(n_1361)
);

NOR2x1_ASAP7_75t_SL g1362 ( 
.A(n_1283),
.B(n_1279),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1327),
.B(n_1260),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1309),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1289),
.B(n_1282),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1290),
.B(n_1319),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1309),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1352),
.B(n_1330),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1359),
.A2(n_1328),
.B1(n_1298),
.B2(n_1258),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1336),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1343),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1350),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1345),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1355),
.B(n_1288),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1339),
.B(n_1321),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1358),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1361),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1366),
.B(n_1299),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1350),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1338),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1349),
.B(n_1304),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1366),
.B(n_1286),
.Y(n_1382)
);

NAND2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1340),
.B(n_1290),
.Y(n_1383)
);

AOI322xp5_ASAP7_75t_L g1384 ( 
.A1(n_1359),
.A2(n_1328),
.A3(n_1258),
.B1(n_1259),
.B2(n_1281),
.C1(n_1218),
.C2(n_1311),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1353),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1353),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1334),
.Y(n_1387)
);

O2A1O1Ixp5_ASAP7_75t_R g1388 ( 
.A1(n_1360),
.A2(n_1329),
.B(n_1275),
.C(n_1325),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1334),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_SL g1390 ( 
.A1(n_1388),
.A2(n_1362),
.B(n_1363),
.C(n_1351),
.Y(n_1390)
);

INVxp67_ASAP7_75t_L g1391 ( 
.A(n_1368),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1369),
.A2(n_1342),
.B1(n_1274),
.B2(n_1259),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1373),
.Y(n_1393)
);

OAI22x1_ASAP7_75t_L g1394 ( 
.A1(n_1383),
.A2(n_1337),
.B1(n_1365),
.B2(n_1325),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1382),
.B(n_1342),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1376),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1369),
.A2(n_1274),
.B1(n_1326),
.B2(n_1304),
.Y(n_1397)
);

INVx2_ASAP7_75t_SL g1398 ( 
.A(n_1374),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1377),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1381),
.A2(n_1326),
.B1(n_1310),
.B2(n_1302),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1380),
.A2(n_1326),
.B1(n_1371),
.B2(n_1370),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1379),
.A2(n_1302),
.B1(n_1263),
.B2(n_1246),
.Y(n_1402)
);

XOR2x2_ASAP7_75t_L g1403 ( 
.A(n_1384),
.B(n_1301),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1393),
.Y(n_1404)
);

AOI222xp33_ASAP7_75t_L g1405 ( 
.A1(n_1403),
.A2(n_1384),
.B1(n_1322),
.B2(n_1378),
.C1(n_1385),
.C2(n_1386),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1391),
.B(n_1378),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1392),
.A2(n_1375),
.B1(n_1294),
.B2(n_1302),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1397),
.A2(n_1331),
.B1(n_1333),
.B2(n_1225),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1396),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1399),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1402),
.A2(n_1294),
.B1(n_1372),
.B2(n_1357),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1390),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1394),
.A2(n_1324),
.B1(n_1307),
.B2(n_1313),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1395),
.A2(n_1263),
.B1(n_1276),
.B2(n_1356),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1401),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1398),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1400),
.B(n_1387),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1393),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1404),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1412),
.B(n_1231),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1416),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1405),
.B(n_1413),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1415),
.B(n_1389),
.Y(n_1423)
);

OAI221xp5_ASAP7_75t_L g1424 ( 
.A1(n_1413),
.A2(n_1407),
.B1(n_1411),
.B2(n_1408),
.C(n_1414),
.Y(n_1424)
);

NAND3xp33_ASAP7_75t_SL g1425 ( 
.A(n_1417),
.B(n_1243),
.C(n_1271),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1410),
.B(n_1356),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1406),
.B(n_1266),
.Y(n_1427)
);

AOI211xp5_ASAP7_75t_L g1428 ( 
.A1(n_1422),
.A2(n_1424),
.B(n_1425),
.C(n_1420),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1427),
.A2(n_1418),
.B(n_1409),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1419),
.Y(n_1430)
);

NOR2x1_ASAP7_75t_L g1431 ( 
.A(n_1421),
.B(n_1278),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1423),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1426),
.B(n_1338),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1429),
.A2(n_1276),
.B(n_1271),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1428),
.B(n_1266),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1430),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_L g1437 ( 
.A(n_1432),
.B(n_1269),
.C(n_1250),
.Y(n_1437)
);

AOI211x1_ASAP7_75t_SL g1438 ( 
.A1(n_1433),
.A2(n_1297),
.B(n_1367),
.C(n_1354),
.Y(n_1438)
);

OAI222xp33_ASAP7_75t_L g1439 ( 
.A1(n_1431),
.A2(n_1367),
.B1(n_1364),
.B2(n_1354),
.C1(n_1335),
.C2(n_1344),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1436),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_SL g1441 ( 
.A(n_1435),
.B(n_1231),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1434),
.B(n_1335),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1437),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1438),
.B(n_1344),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1439),
.Y(n_1445)
);

NOR2xp67_ASAP7_75t_L g1446 ( 
.A(n_1435),
.B(n_1245),
.Y(n_1446)
);

NOR2x1_ASAP7_75t_L g1447 ( 
.A(n_1435),
.B(n_1270),
.Y(n_1447)
);

NOR2x1_ASAP7_75t_L g1448 ( 
.A(n_1440),
.B(n_1270),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1443),
.Y(n_1449)
);

OAI22x1_ASAP7_75t_L g1450 ( 
.A1(n_1447),
.A2(n_1445),
.B1(n_1441),
.B2(n_1446),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1442),
.B(n_1364),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_L g1452 ( 
.A(n_1444),
.B(n_1270),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1443),
.B(n_1245),
.Y(n_1453)
);

NOR2x1_ASAP7_75t_L g1454 ( 
.A(n_1440),
.B(n_1250),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1449),
.Y(n_1455)
);

AOI221xp5_ASAP7_75t_L g1456 ( 
.A1(n_1450),
.A2(n_1297),
.B1(n_1249),
.B2(n_1248),
.C(n_1312),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1453),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1448),
.Y(n_1458)
);

AOI222xp33_ASAP7_75t_L g1459 ( 
.A1(n_1452),
.A2(n_1454),
.B1(n_1451),
.B2(n_1248),
.C1(n_1297),
.C2(n_1249),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1449),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1449),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1458),
.Y(n_1462)
);

CKINVDCx20_ASAP7_75t_R g1463 ( 
.A(n_1461),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1457),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1460),
.B(n_1455),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1457),
.A2(n_1249),
.B1(n_1297),
.B2(n_1247),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1456),
.A2(n_1348),
.B1(n_1347),
.B2(n_1346),
.Y(n_1467)
);

XNOR2x1_ASAP7_75t_L g1468 ( 
.A(n_1459),
.B(n_264),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1458),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1458),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1461),
.A2(n_1341),
.B1(n_1300),
.B2(n_1348),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1469),
.A2(n_1346),
.B1(n_1347),
.B2(n_269),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1463),
.Y(n_1473)
);

OAI31xp33_ASAP7_75t_L g1474 ( 
.A1(n_1462),
.A2(n_266),
.A3(n_268),
.B(n_270),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1470),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1464),
.Y(n_1476)
);

AOI31xp33_ASAP7_75t_L g1477 ( 
.A1(n_1465),
.A2(n_276),
.A3(n_277),
.B(n_278),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1468),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_1478)
);

AOI31xp33_ASAP7_75t_L g1479 ( 
.A1(n_1471),
.A2(n_1466),
.A3(n_1467),
.B(n_293),
.Y(n_1479)
);

OAI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1469),
.A2(n_287),
.B1(n_291),
.B2(n_294),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1463),
.A2(n_297),
.B1(n_301),
.B2(n_303),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1475),
.B(n_304),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_SL g1483 ( 
.A1(n_1473),
.A2(n_1478),
.B1(n_1476),
.B2(n_1472),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1479),
.A2(n_305),
.B1(n_307),
.B2(n_310),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_SL g1485 ( 
.A1(n_1481),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1477),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1480),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1474),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1473),
.Y(n_1489)
);

O2A1O1Ixp5_ASAP7_75t_SL g1490 ( 
.A1(n_1488),
.A2(n_314),
.B(n_315),
.C(n_317),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1489),
.A2(n_319),
.B1(n_322),
.B2(n_323),
.Y(n_1491)
);

XNOR2xp5_ASAP7_75t_L g1492 ( 
.A(n_1483),
.B(n_1484),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1482),
.Y(n_1493)
);

OAI211xp5_ASAP7_75t_L g1494 ( 
.A1(n_1487),
.A2(n_1486),
.B(n_1485),
.C(n_327),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1493),
.B(n_324),
.Y(n_1495)
);

XNOR2xp5_ASAP7_75t_L g1496 ( 
.A(n_1492),
.B(n_326),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1494),
.A2(n_329),
.B(n_331),
.Y(n_1497)
);

NOR2x1_ASAP7_75t_SL g1498 ( 
.A(n_1495),
.B(n_1490),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_R g1499 ( 
.A1(n_1496),
.A2(n_1491),
.B1(n_332),
.B2(n_333),
.Y(n_1499)
);

OR2x6_ASAP7_75t_L g1500 ( 
.A(n_1499),
.B(n_1497),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1500),
.A2(n_1498),
.B1(n_334),
.B2(n_335),
.Y(n_1501)
);


endmodule