module fake_aes_2149_n_625 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_625);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_625;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_31), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_21), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_10), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_14), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_9), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_33), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_36), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_52), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_34), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_57), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_75), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_53), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_37), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_46), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_4), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_14), .Y(n_92) );
INVx1_ASAP7_75t_SL g93 ( .A(n_27), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_28), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_55), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_67), .Y(n_96) );
HB1xp67_ASAP7_75t_L g97 ( .A(n_66), .Y(n_97) );
BUFx6f_ASAP7_75t_L g98 ( .A(n_8), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_6), .Y(n_99) );
BUFx6f_ASAP7_75t_L g100 ( .A(n_49), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_54), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_65), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_62), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_24), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_44), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_20), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_71), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_35), .Y(n_108) );
INVx2_ASAP7_75t_SL g109 ( .A(n_12), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_73), .Y(n_110) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_19), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_6), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_58), .Y(n_113) );
INVxp33_ASAP7_75t_SL g114 ( .A(n_8), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_16), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_1), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_42), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_70), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_16), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_30), .Y(n_120) );
NOR2xp67_ASAP7_75t_L g121 ( .A(n_40), .B(n_63), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_60), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_4), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_9), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_83), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_97), .B(n_0), .Y(n_126) );
CKINVDCx16_ASAP7_75t_R g127 ( .A(n_111), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_77), .Y(n_128) );
CKINVDCx11_ASAP7_75t_R g129 ( .A(n_108), .Y(n_129) );
CKINVDCx16_ASAP7_75t_R g130 ( .A(n_107), .Y(n_130) );
BUFx3_ASAP7_75t_L g131 ( .A(n_95), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_109), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_77), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_100), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_109), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_114), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_100), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_79), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_79), .B(n_0), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_100), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_78), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_81), .B(n_91), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_78), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_114), .Y(n_145) );
AND2x6_ASAP7_75t_L g146 ( .A(n_95), .B(n_38), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_81), .B(n_1), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_84), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_82), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_91), .B(n_2), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_93), .Y(n_151) );
NOR2xp33_ASAP7_75t_R g152 ( .A(n_101), .B(n_39), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_100), .Y(n_153) );
NAND2x1_ASAP7_75t_L g154 ( .A(n_92), .B(n_2), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_85), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_92), .B(n_3), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_89), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_100), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_115), .B(n_3), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_112), .B(n_5), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_85), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_87), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_115), .B(n_5), .Y(n_163) );
NAND2xp33_ASAP7_75t_SL g164 ( .A(n_116), .B(n_7), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_116), .B(n_7), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_124), .B(n_10), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_119), .B(n_11), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
AO22x2_ASAP7_75t_L g169 ( .A1(n_147), .A2(n_123), .B1(n_119), .B2(n_80), .Y(n_169) );
BUFx4f_ASAP7_75t_L g170 ( .A(n_147), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_147), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_156), .Y(n_175) );
NAND2x1p5_ASAP7_75t_L g176 ( .A(n_139), .B(n_123), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_156), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_128), .B(n_82), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
INVxp33_ASAP7_75t_L g180 ( .A(n_138), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_134), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_142), .B(n_99), .Y(n_182) );
INVx5_ASAP7_75t_L g183 ( .A(n_146), .Y(n_183) );
INVxp67_ASAP7_75t_L g184 ( .A(n_126), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_134), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_157), .B(n_118), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_140), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_156), .Y(n_188) );
AND2x4_ASAP7_75t_SL g189 ( .A(n_132), .B(n_98), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_134), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_159), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_146), .Y(n_192) );
INVxp67_ASAP7_75t_L g193 ( .A(n_142), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_127), .B(n_118), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_128), .B(n_120), .Y(n_195) );
NAND2x1p5_ASAP7_75t_L g196 ( .A(n_139), .B(n_122), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_159), .B(n_122), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_159), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_159), .Y(n_199) );
AND2x6_ASAP7_75t_L g200 ( .A(n_150), .B(n_88), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_131), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_150), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_131), .Y(n_203) );
INVxp67_ASAP7_75t_L g204 ( .A(n_163), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_133), .B(n_120), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_133), .A2(n_98), .B1(n_117), .B2(n_90), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_141), .B(n_88), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_163), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_127), .B(n_102), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_140), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_165), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_137), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_151), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_141), .B(n_94), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_130), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_165), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_143), .B(n_103), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_143), .B(n_105), .Y(n_218) );
AND2x2_ASAP7_75t_SL g219 ( .A(n_167), .B(n_90), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_149), .Y(n_220) );
INVxp67_ASAP7_75t_L g221 ( .A(n_167), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_144), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_144), .B(n_94), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_146), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_140), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_140), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_148), .B(n_104), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_148), .B(n_96), .Y(n_228) );
INVx1_ASAP7_75t_SL g229 ( .A(n_215), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_184), .B(n_162), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_193), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_204), .B(n_221), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_184), .B(n_162), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_176), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_222), .B(n_161), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_207), .B(n_161), .Y(n_237) );
INVxp67_ASAP7_75t_L g238 ( .A(n_213), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_174), .Y(n_239) );
INVx2_ASAP7_75t_SL g240 ( .A(n_196), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_204), .B(n_155), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_168), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_174), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_219), .A2(n_155), .B1(n_130), .B2(n_160), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_192), .Y(n_245) );
NOR2xp33_ASAP7_75t_R g246 ( .A(n_170), .B(n_125), .Y(n_246) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_180), .Y(n_247) );
INVx4_ASAP7_75t_L g248 ( .A(n_183), .Y(n_248) );
CKINVDCx8_ASAP7_75t_R g249 ( .A(n_200), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_194), .B(n_136), .Y(n_250) );
INVx8_ASAP7_75t_L g251 ( .A(n_200), .Y(n_251) );
NAND3xp33_ASAP7_75t_SL g252 ( .A(n_180), .B(n_145), .C(n_135), .Y(n_252) );
AND2x6_ASAP7_75t_L g253 ( .A(n_172), .B(n_96), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_176), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_189), .Y(n_255) );
CKINVDCx11_ASAP7_75t_R g256 ( .A(n_182), .Y(n_256) );
OR2x6_ASAP7_75t_L g257 ( .A(n_169), .B(n_154), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_189), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_221), .B(n_166), .Y(n_259) );
NAND3xp33_ASAP7_75t_SL g260 ( .A(n_209), .B(n_154), .C(n_164), .Y(n_260) );
AOI21xp33_ASAP7_75t_L g261 ( .A1(n_169), .A2(n_113), .B(n_106), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_207), .B(n_146), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_223), .B(n_146), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_201), .Y(n_264) );
BUFx3_ASAP7_75t_L g265 ( .A(n_220), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_192), .B(n_152), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_219), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_182), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_203), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_224), .B(n_110), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_196), .B(n_129), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_223), .Y(n_272) );
AOI21x1_ASAP7_75t_L g273 ( .A1(n_214), .A2(n_149), .B(n_87), .Y(n_273) );
AND2x6_ASAP7_75t_L g274 ( .A(n_175), .B(n_117), .Y(n_274) );
OR2x4_ASAP7_75t_L g275 ( .A(n_186), .B(n_98), .Y(n_275) );
INVx1_ASAP7_75t_SL g276 ( .A(n_200), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_228), .B(n_146), .Y(n_277) );
AND2x6_ASAP7_75t_L g278 ( .A(n_177), .B(n_101), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_228), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_170), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_200), .B(n_146), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_181), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_197), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_200), .B(n_86), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_224), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_169), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_202), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_197), .B(n_98), .Y(n_288) );
AND2x6_ASAP7_75t_L g289 ( .A(n_179), .B(n_98), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_188), .B(n_121), .Y(n_290) );
NOR3xp33_ASAP7_75t_SL g291 ( .A(n_186), .B(n_11), .C(n_12), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_191), .B(n_158), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_181), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_230), .B(n_211), .Y(n_294) );
OAI21xp33_ASAP7_75t_L g295 ( .A1(n_230), .A2(n_208), .B(n_216), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_247), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_282), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_262), .A2(n_183), .B(n_199), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_245), .Y(n_299) );
NOR2x1_ASAP7_75t_SL g300 ( .A(n_257), .B(n_183), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g301 ( .A1(n_261), .A2(n_198), .B(n_227), .C(n_205), .Y(n_301) );
CKINVDCx11_ASAP7_75t_R g302 ( .A(n_229), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_245), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_245), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_234), .B(n_227), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_240), .B(n_183), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_285), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_229), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_255), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_234), .B(n_218), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_262), .A2(n_195), .B(n_178), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_258), .Y(n_312) );
OAI21xp33_ASAP7_75t_L g313 ( .A1(n_250), .A2(n_206), .B(n_217), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_293), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_286), .A2(n_214), .B1(n_178), .B2(n_195), .Y(n_315) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_276), .B(n_205), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_235), .B(n_206), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_233), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_259), .B(n_13), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_239), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_285), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_239), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_243), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_243), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_251), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_285), .B(n_185), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_249), .A2(n_137), .B1(n_158), .B2(n_190), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_259), .B(n_13), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_241), .B(n_15), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_251), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_254), .B(n_15), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_236), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_251), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_233), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_242), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_268), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_256), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_275), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_246), .Y(n_339) );
NOR2xp67_ASAP7_75t_L g340 ( .A(n_260), .B(n_64), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_241), .B(n_17), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_244), .A2(n_137), .B1(n_158), .B2(n_212), .C(n_190), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_264), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_236), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_308), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_332), .Y(n_346) );
OAI22xp33_ASAP7_75t_L g347 ( .A1(n_308), .A2(n_244), .B1(n_267), .B2(n_257), .Y(n_347) );
AO21x2_ASAP7_75t_L g348 ( .A1(n_301), .A2(n_261), .B(n_291), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_310), .B(n_252), .Y(n_349) );
BUFx10_ASAP7_75t_L g350 ( .A(n_330), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_299), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_297), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_332), .B(n_237), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_344), .A2(n_237), .B1(n_275), .B2(n_276), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_297), .Y(n_355) );
CKINVDCx6p67_ASAP7_75t_R g356 ( .A(n_302), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_344), .B(n_231), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_341), .A2(n_257), .B1(n_232), .B2(n_283), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_341), .A2(n_287), .B1(n_272), .B2(n_279), .Y(n_359) );
INVx6_ASAP7_75t_L g360 ( .A(n_330), .Y(n_360) );
XNOR2xp5_ASAP7_75t_L g361 ( .A(n_337), .B(n_271), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_296), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_314), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_310), .B(n_283), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_296), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_294), .B(n_253), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_341), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_314), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_294), .B(n_280), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_299), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_317), .A2(n_253), .B1(n_274), .B2(n_284), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_325), .B(n_265), .Y(n_372) );
OAI21x1_ASAP7_75t_L g373 ( .A1(n_298), .A2(n_273), .B(n_281), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_318), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_305), .B(n_263), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_330), .Y(n_376) );
AOI222xp33_ASAP7_75t_L g377 ( .A1(n_347), .A2(n_319), .B1(n_295), .B2(n_334), .C1(n_328), .C2(n_331), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_346), .B(n_319), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_346), .B(n_375), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_350), .Y(n_380) );
AOI21xp33_ASAP7_75t_L g381 ( .A1(n_348), .A2(n_338), .B(n_329), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_352), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_359), .A2(n_313), .B1(n_317), .B2(n_274), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_352), .Y(n_384) );
NAND3xp33_ASAP7_75t_L g385 ( .A(n_354), .B(n_340), .C(n_342), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_359), .A2(n_338), .B1(n_339), .B2(n_300), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_349), .A2(n_253), .B1(n_274), .B2(n_317), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_367), .A2(n_316), .B1(n_290), .B2(n_288), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_353), .B(n_367), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_358), .A2(n_316), .B1(n_290), .B2(n_288), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_349), .A2(n_339), .B1(n_336), .B2(n_238), .Y(n_391) );
OA21x2_ASAP7_75t_L g392 ( .A1(n_373), .A2(n_311), .B(n_340), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_353), .B(n_335), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_366), .A2(n_316), .B1(n_277), .B2(n_263), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_368), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_375), .B(n_364), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_352), .Y(n_398) );
AOI33xp33_ASAP7_75t_L g399 ( .A1(n_369), .A2(n_315), .A3(n_320), .B1(n_322), .B2(n_185), .B3(n_212), .Y(n_399) );
OAI21x1_ASAP7_75t_L g400 ( .A1(n_373), .A2(n_281), .B(n_327), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_345), .A2(n_253), .B1(n_274), .B2(n_278), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_365), .B(n_312), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_355), .Y(n_403) );
AO21x2_ASAP7_75t_L g404 ( .A1(n_348), .A2(n_277), .B(n_292), .Y(n_404) );
OAI33xp33_ASAP7_75t_L g405 ( .A1(n_391), .A2(n_354), .A3(n_357), .B1(n_366), .B2(n_364), .B3(n_348), .Y(n_405) );
INVxp67_ASAP7_75t_L g406 ( .A(n_393), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_395), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_382), .Y(n_408) );
INVx5_ASAP7_75t_SL g409 ( .A(n_389), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_382), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_377), .A2(n_345), .B1(n_348), .B2(n_369), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_382), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_384), .Y(n_413) );
OA21x2_ASAP7_75t_L g414 ( .A1(n_381), .A2(n_373), .B(n_370), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_403), .B(n_355), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_395), .B(n_365), .Y(n_416) );
AO21x2_ASAP7_75t_L g417 ( .A1(n_381), .A2(n_370), .B(n_357), .Y(n_417) );
OAI21x1_ASAP7_75t_L g418 ( .A1(n_400), .A2(n_392), .B(n_390), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_384), .Y(n_419) );
BUFx4f_ASAP7_75t_SL g420 ( .A(n_380), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_397), .B(n_362), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_380), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_403), .B(n_355), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_398), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_377), .A2(n_369), .B1(n_362), .B2(n_356), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_402), .B(n_361), .Y(n_427) );
NOR2x2_ASAP7_75t_L g428 ( .A(n_398), .B(n_356), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_398), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_393), .Y(n_431) );
NAND4xp25_ASAP7_75t_L g432 ( .A(n_402), .B(n_369), .C(n_371), .D(n_292), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_380), .B(n_370), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_383), .A2(n_363), .B1(n_374), .B2(n_356), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_392), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_396), .A2(n_374), .B1(n_361), .B2(n_278), .Y(n_436) );
OAI31xp33_ASAP7_75t_SL g437 ( .A1(n_386), .A2(n_390), .A3(n_389), .B(n_388), .Y(n_437) );
AOI211xp5_ASAP7_75t_SL g438 ( .A1(n_383), .A2(n_376), .B(n_363), .C(n_372), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_420), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
AOI33xp33_ASAP7_75t_L g441 ( .A1(n_426), .A2(n_378), .A3(n_396), .B1(n_387), .B2(n_389), .B3(n_401), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_432), .A2(n_389), .B1(n_378), .B2(n_379), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_410), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_410), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_406), .B(n_379), .Y(n_445) );
INVx5_ASAP7_75t_L g446 ( .A(n_422), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_413), .B(n_404), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_406), .B(n_404), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_431), .B(n_17), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_431), .B(n_404), .Y(n_450) );
INVx4_ASAP7_75t_L g451 ( .A(n_420), .Y(n_451) );
OAI33xp33_ASAP7_75t_L g452 ( .A1(n_434), .A2(n_388), .A3(n_394), .B1(n_385), .B2(n_320), .B3(n_322), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_416), .B(n_404), .Y(n_453) );
INVx6_ASAP7_75t_L g454 ( .A(n_433), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_413), .B(n_363), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_407), .B(n_399), .Y(n_456) );
NOR2xp33_ASAP7_75t_SL g457 ( .A(n_432), .B(n_350), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_423), .B(n_421), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_423), .B(n_394), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_408), .Y(n_460) );
OAI21xp33_ASAP7_75t_L g461 ( .A1(n_437), .A2(n_385), .B(n_153), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_421), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_422), .B(n_400), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_427), .B(n_18), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_416), .B(n_18), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_408), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_415), .B(n_372), .Y(n_467) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_422), .B(n_376), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_415), .B(n_392), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_412), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_437), .B(n_351), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_436), .A2(n_372), .B1(n_351), .B2(n_360), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_409), .B(n_351), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_409), .B(n_309), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_405), .A2(n_372), .B1(n_153), .B2(n_324), .C(n_323), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_415), .B(n_376), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_424), .B(n_400), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_424), .B(n_376), .Y(n_478) );
NAND2x1p5_ASAP7_75t_L g479 ( .A(n_422), .B(n_330), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_412), .Y(n_480) );
OAI33xp33_ASAP7_75t_L g481 ( .A1(n_434), .A2(n_324), .A3(n_323), .B1(n_343), .B2(n_335), .B3(n_326), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_412), .B(n_300), .Y(n_482) );
NAND2xp33_ASAP7_75t_SL g483 ( .A(n_428), .B(n_330), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_419), .B(n_343), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_458), .B(n_409), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_481), .A2(n_438), .B(n_405), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_462), .B(n_411), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_443), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_442), .B(n_433), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_477), .B(n_417), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_477), .B(n_417), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_469), .B(n_417), .Y(n_492) );
OAI33xp33_ASAP7_75t_L g493 ( .A1(n_465), .A2(n_435), .A3(n_430), .B1(n_425), .B2(n_429), .B3(n_419), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_469), .B(n_417), .Y(n_494) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_443), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_483), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_457), .B(n_433), .Y(n_497) );
NAND5xp2_ASAP7_75t_SL g498 ( .A(n_464), .B(n_438), .C(n_409), .D(n_25), .E(n_26), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_470), .Y(n_499) );
BUFx2_ASAP7_75t_L g500 ( .A(n_483), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_440), .Y(n_501) );
NAND5xp2_ASAP7_75t_SL g502 ( .A(n_449), .B(n_409), .C(n_23), .D(n_29), .E(n_32), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_467), .B(n_409), .Y(n_503) );
HB1xp67_ASAP7_75t_SL g504 ( .A(n_439), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_445), .B(n_419), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_439), .Y(n_506) );
OR2x6_ASAP7_75t_L g507 ( .A(n_444), .B(n_418), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_463), .B(n_435), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_447), .B(n_430), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_455), .B(n_429), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_440), .Y(n_511) );
NAND4xp25_ASAP7_75t_SL g512 ( .A(n_441), .B(n_429), .C(n_425), .D(n_430), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_450), .B(n_418), .Y(n_513) );
CKINVDCx14_ASAP7_75t_R g514 ( .A(n_451), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_453), .B(n_425), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_456), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_461), .B(n_153), .C(n_414), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_476), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_478), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_460), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_441), .B(n_414), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_471), .A2(n_278), .B1(n_414), .B2(n_360), .Y(n_522) );
BUFx3_ASAP7_75t_L g523 ( .A(n_451), .Y(n_523) );
OAI221xp5_ASAP7_75t_L g524 ( .A1(n_471), .A2(n_414), .B1(n_360), .B2(n_153), .C(n_304), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_448), .B(n_480), .Y(n_525) );
OAI221xp5_ASAP7_75t_L g526 ( .A1(n_474), .A2(n_360), .B1(n_153), .B2(n_321), .C(n_304), .Y(n_526) );
NAND5xp2_ASAP7_75t_L g527 ( .A(n_475), .B(n_278), .C(n_350), .D(n_43), .E(n_45), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_466), .B(n_153), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_517), .A2(n_452), .B(n_482), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_489), .A2(n_472), .B1(n_454), .B2(n_482), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_488), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_506), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_516), .B(n_459), .Y(n_533) );
OAI21xp33_ASAP7_75t_L g534 ( .A1(n_512), .A2(n_463), .B(n_482), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_514), .A2(n_446), .B(n_468), .C(n_473), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_493), .A2(n_480), .B1(n_484), .B2(n_446), .C(n_225), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_500), .B(n_446), .Y(n_537) );
INVxp67_ASAP7_75t_L g538 ( .A(n_495), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_518), .B(n_446), .Y(n_539) );
AOI321xp33_ASAP7_75t_L g540 ( .A1(n_489), .A2(n_269), .A3(n_266), .B1(n_270), .B2(n_479), .C(n_306), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_505), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_499), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_519), .B(n_22), .Y(n_543) );
AOI222xp33_ASAP7_75t_SL g544 ( .A1(n_496), .A2(n_289), .B1(n_321), .B2(n_48), .C1(n_50), .C2(n_51), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_524), .A2(n_307), .B(n_299), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_498), .A2(n_333), .B(n_325), .C(n_306), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_487), .A2(n_350), .B1(n_289), .B2(n_303), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_499), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_509), .B(n_41), .Y(n_549) );
AOI321xp33_ASAP7_75t_L g550 ( .A1(n_521), .A2(n_306), .A3(n_56), .B1(n_59), .B2(n_61), .C(n_68), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_492), .B(n_47), .Y(n_551) );
NAND2x1_ASAP7_75t_L g552 ( .A(n_507), .B(n_289), .Y(n_552) );
INVx2_ASAP7_75t_SL g553 ( .A(n_506), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_525), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_492), .B(n_69), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g556 ( .A1(n_522), .A2(n_225), .B1(n_226), .B2(n_210), .C(n_171), .Y(n_556) );
NOR3xp33_ASAP7_75t_L g557 ( .A(n_526), .B(n_72), .C(n_74), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_523), .B(n_307), .Y(n_558) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_523), .A2(n_307), .B1(n_303), .B2(n_299), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_504), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_486), .A2(n_307), .B(n_303), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_510), .B(n_515), .Y(n_562) );
OAI221xp5_ASAP7_75t_L g563 ( .A1(n_507), .A2(n_226), .B1(n_171), .B2(n_173), .C(n_187), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_485), .B(n_76), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_494), .B(n_289), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_536), .B(n_497), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_533), .B(n_490), .Y(n_567) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_533), .A2(n_491), .B1(n_490), .B2(n_513), .C(n_502), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_558), .A2(n_497), .B(n_507), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_554), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_560), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_562), .B(n_491), .Y(n_572) );
NAND2xp33_ASAP7_75t_L g573 ( .A(n_535), .B(n_503), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_541), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_538), .B(n_508), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_532), .Y(n_576) );
NAND2xp33_ASAP7_75t_SL g577 ( .A(n_537), .B(n_508), .Y(n_577) );
XNOR2xp5_ASAP7_75t_L g578 ( .A(n_553), .B(n_513), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_531), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_531), .B(n_508), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_542), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_538), .B(n_527), .Y(n_582) );
XOR2x2_ASAP7_75t_L g583 ( .A(n_530), .B(n_528), .Y(n_583) );
AOI221xp5_ASAP7_75t_SL g584 ( .A1(n_534), .A2(n_520), .B1(n_511), .B2(n_501), .C(n_210), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_539), .B(n_520), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_548), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_529), .Y(n_587) );
OAI21xp5_ASAP7_75t_L g588 ( .A1(n_557), .A2(n_248), .B(n_303), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_577), .B(n_559), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_587), .A2(n_551), .B1(n_555), .B2(n_543), .C(n_561), .Y(n_590) );
XNOR2x1_ASAP7_75t_L g591 ( .A(n_571), .B(n_564), .Y(n_591) );
AOI222xp33_ASAP7_75t_L g592 ( .A1(n_587), .A2(n_549), .B1(n_565), .B2(n_563), .C1(n_556), .C2(n_547), .Y(n_592) );
OAI211xp5_ASAP7_75t_SL g593 ( .A1(n_576), .A2(n_550), .B(n_540), .C(n_547), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_578), .Y(n_594) );
INVxp67_ASAP7_75t_SL g595 ( .A(n_581), .Y(n_595) );
XNOR2xp5_ASAP7_75t_L g596 ( .A(n_583), .B(n_552), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_582), .A2(n_545), .B1(n_544), .B2(n_299), .Y(n_597) );
OAI21xp33_ASAP7_75t_L g598 ( .A1(n_567), .A2(n_546), .B(n_187), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_584), .A2(n_173), .B1(n_187), .B2(n_210), .C(n_225), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_579), .A2(n_173), .B1(n_187), .B2(n_210), .C(n_225), .Y(n_600) );
OAI221xp5_ASAP7_75t_L g601 ( .A1(n_582), .A2(n_173), .B1(n_226), .B2(n_568), .C(n_573), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_570), .B(n_226), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_566), .A2(n_580), .B1(n_585), .B2(n_575), .Y(n_603) );
XNOR2xp5_ASAP7_75t_L g604 ( .A(n_572), .B(n_574), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_598), .B(n_566), .C(n_588), .Y(n_605) );
AND2x2_ASAP7_75t_SL g606 ( .A(n_597), .B(n_575), .Y(n_606) );
NAND2xp33_ASAP7_75t_R g607 ( .A(n_594), .B(n_569), .Y(n_607) );
NAND2x1p5_ASAP7_75t_L g608 ( .A(n_589), .B(n_591), .Y(n_608) );
BUFx2_ASAP7_75t_L g609 ( .A(n_596), .Y(n_609) );
AOI211xp5_ASAP7_75t_L g610 ( .A1(n_593), .A2(n_586), .B(n_599), .C(n_590), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_602), .A2(n_587), .B1(n_601), .B2(n_604), .C(n_579), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_600), .A2(n_587), .B1(n_601), .B2(n_604), .C(n_579), .Y(n_612) );
AO22x1_ASAP7_75t_L g613 ( .A1(n_592), .A2(n_594), .B1(n_560), .B2(n_595), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_603), .A2(n_587), .B1(n_593), .B2(n_601), .Y(n_614) );
NOR3xp33_ASAP7_75t_SL g615 ( .A(n_607), .B(n_611), .C(n_612), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_609), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_613), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_616), .A2(n_608), .B(n_606), .Y(n_618) );
NOR3xp33_ASAP7_75t_L g619 ( .A(n_617), .B(n_605), .C(n_610), .Y(n_619) );
XNOR2xp5_ASAP7_75t_L g620 ( .A(n_615), .B(n_614), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_620), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_618), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_621), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_623), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_624), .A2(n_622), .B(n_619), .Y(n_625) );
endmodule