module fake_jpeg_7051_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_45),
.Y(n_53)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_47),
.B1(n_18),
.B2(n_24),
.Y(n_62)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_22),
.B1(n_27),
.B2(n_17),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_52),
.A2(n_61),
.B1(n_73),
.B2(n_23),
.Y(n_95)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_59),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_22),
.B1(n_27),
.B2(n_17),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_55),
.A2(n_65),
.B1(n_32),
.B2(n_40),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_56),
.B(n_68),
.Y(n_96)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_27),
.B1(n_21),
.B2(n_24),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_25),
.B1(n_21),
.B2(n_31),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_24),
.Y(n_68)
);

AND2x4_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_33),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_23),
.B(n_33),
.C(n_41),
.Y(n_89)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_34),
.B1(n_31),
.B2(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_81),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_80),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_85),
.Y(n_110)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_91),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_30),
.B(n_26),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_89),
.B(n_91),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_69),
.A2(n_34),
.B1(n_43),
.B2(n_32),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_97),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_52),
.B1(n_73),
.B2(n_56),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_108),
.Y(n_133)
);

AOI32xp33_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_69),
.A3(n_53),
.B1(n_55),
.B2(n_49),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_SL g139 ( 
.A(n_102),
.B(n_126),
.Y(n_139)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_107),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_98),
.A2(n_63),
.B1(n_70),
.B2(n_71),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_122),
.B1(n_83),
.B2(n_78),
.Y(n_131)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_53),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_61),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_112),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_128),
.B1(n_78),
.B2(n_76),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_20),
.B(n_33),
.Y(n_149)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_119),
.Y(n_156)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_85),
.A2(n_54),
.B1(n_50),
.B2(n_58),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_127),
.B(n_29),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_82),
.A2(n_72),
.B1(n_50),
.B2(n_40),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_57),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_33),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_89),
.B(n_57),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_59),
.B1(n_67),
.B2(n_14),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_82),
.A2(n_41),
.B1(n_40),
.B2(n_37),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_86),
.B1(n_83),
.B2(n_76),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_135),
.B1(n_136),
.B2(n_141),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_120),
.B1(n_125),
.B2(n_104),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_75),
.B1(n_79),
.B2(n_41),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_137),
.Y(n_172)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_101),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_140),
.B(n_142),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_126),
.B1(n_102),
.B2(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_75),
.B1(n_79),
.B2(n_37),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_144),
.B1(n_147),
.B2(n_122),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_37),
.B1(n_93),
.B2(n_67),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_67),
.B1(n_77),
.B2(n_33),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_107),
.B(n_0),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_151),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_153),
.B(n_30),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_125),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_111),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

AO22x1_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_30),
.B1(n_26),
.B2(n_20),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_26),
.B(n_100),
.C(n_29),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_108),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_159),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_117),
.B(n_112),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_160),
.A2(n_174),
.B(n_177),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_105),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_167),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_117),
.B1(n_114),
.B2(n_113),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_166),
.B1(n_178),
.B2(n_182),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_104),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_157),
.B1(n_142),
.B2(n_134),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_110),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_110),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_150),
.B(n_109),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_175),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_148),
.B(n_157),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_133),
.A2(n_118),
.B(n_20),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_29),
.C(n_19),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_185),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_135),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_153),
.B1(n_168),
.B2(n_170),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_131),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_140),
.A2(n_1),
.B(n_2),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_162),
.B(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_3),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_189),
.B(n_193),
.Y(n_233)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_194),
.B(n_196),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_151),
.C(n_164),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_199),
.B(n_201),
.Y(n_224)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_172),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_203),
.A2(n_187),
.B(n_194),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_163),
.A2(n_143),
.B1(n_144),
.B2(n_147),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_204),
.A2(n_211),
.B1(n_213),
.B2(n_169),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_207),
.B1(n_212),
.B2(n_171),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_184),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_208),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_176),
.A2(n_181),
.B1(n_163),
.B2(n_175),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_134),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_210),
.A2(n_179),
.B(n_146),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_130),
.B1(n_136),
.B2(n_132),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_174),
.A2(n_152),
.B1(n_156),
.B2(n_137),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_166),
.A2(n_156),
.B1(n_146),
.B2(n_138),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_162),
.A2(n_10),
.B(n_14),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_182),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_167),
.C(n_160),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_225),
.C(n_237),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_183),
.B(n_180),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_216),
.A2(n_236),
.B(n_12),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_241),
.B1(n_200),
.B2(n_208),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_232),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_159),
.C(n_179),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_178),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_231),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_234),
.B(n_203),
.Y(n_246)
);

INVx4_ASAP7_75t_SL g229 ( 
.A(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_184),
.Y(n_230)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_SL g231 ( 
.A(n_202),
.B(n_155),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_3),
.B(n_4),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_190),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_238),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_137),
.C(n_4),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_3),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_196),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_241)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_223),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_201),
.B(n_206),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_254),
.B1(n_256),
.B2(n_264),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_197),
.B(n_204),
.C(n_198),
.Y(n_249)
);

AO21x1_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_239),
.B(n_238),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_197),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_253),
.Y(n_269)
);

NOR3xp33_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_191),
.C(n_189),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_257),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_11),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_221),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_6),
.C(n_7),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_237),
.C(n_263),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_235),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_259),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_12),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_240),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_218),
.B(n_12),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_263),
.C(n_224),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_9),
.Y(n_264)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_220),
.B(n_230),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_245),
.B(n_232),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_270),
.C(n_271),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_250),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_216),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_249),
.B(n_242),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_274),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_275),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_279),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_277),
.B(n_278),
.Y(n_285)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_280),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_228),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_259),
.Y(n_298)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_236),
.C(n_222),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_246),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_218),
.C(n_233),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_269),
.C(n_271),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_287),
.C(n_279),
.Y(n_305)
);

XNOR2x1_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_242),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_267),
.B(n_265),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_288),
.A2(n_294),
.B(n_296),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_253),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_300),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_298),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_260),
.C(n_248),
.Y(n_299)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_258),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_268),
.B(n_248),
.Y(n_301)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_281),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_303),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_243),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_292),
.C(n_294),
.Y(n_319)
);

AO21x2_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_278),
.B(n_251),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_307),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_293),
.A2(n_244),
.B1(n_217),
.B2(n_283),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_309),
.B(n_296),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_243),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_311),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_254),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_256),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_6),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_286),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_297),
.Y(n_315)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_319),
.A2(n_322),
.B(n_302),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_289),
.Y(n_320)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_274),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_321),
.B(n_307),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_7),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_330),
.Y(n_336)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_326),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_318),
.A2(n_307),
.B1(n_304),
.B2(n_303),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_316),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_328),
.A2(n_332),
.B(n_319),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_317),
.B(n_313),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_333),
.B(n_337),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_335),
.A2(n_325),
.B(n_331),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_329),
.A2(n_324),
.B1(n_308),
.B2(n_9),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_338),
.A2(n_336),
.B(n_334),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_339),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_7),
.B(n_9),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_343),
.B(n_9),
.Y(n_344)
);


endmodule