module real_jpeg_30970_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_525;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_0),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_0),
.Y(n_172)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_0),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_541),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_1),
.B(n_542),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_2),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_2),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_2),
.B(n_140),
.Y(n_139)
);

NAND2x1_ASAP7_75t_L g162 ( 
.A(n_2),
.B(n_163),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g291 ( 
.A(n_2),
.B(n_171),
.C(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_2),
.B(n_297),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_2),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_2),
.B(n_292),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_SL g377 ( 
.A(n_2),
.B(n_171),
.C(n_292),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_2),
.B(n_434),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_3),
.Y(n_149)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_4),
.Y(n_91)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_5),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_5),
.Y(n_294)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_5),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_6),
.Y(n_131)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_6),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_6),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_7),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_7),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_7),
.B(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_7),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_SL g204 ( 
.A(n_7),
.B(n_205),
.Y(n_204)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_7),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_7),
.B(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_8),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_9),
.B(n_80),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g132 ( 
.A(n_9),
.B(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_9),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_9),
.B(n_49),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_9),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_9),
.B(n_467),
.Y(n_466)
);

BUFx2_ASAP7_75t_R g527 ( 
.A(n_9),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_10),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_10),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_12),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_13),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_13),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_13),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_13),
.B(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_13),
.B(n_253),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g281 ( 
.A(n_13),
.B(n_188),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_13),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_13),
.B(n_352),
.Y(n_351)
);

AOI22x1_ASAP7_75t_L g108 ( 
.A1(n_14),
.A2(n_15),
.B1(n_109),
.B2(n_112),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g122 ( 
.A(n_14),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_14),
.B(n_188),
.Y(n_187)
);

NAND2x1_ASAP7_75t_L g82 ( 
.A(n_15),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_15),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_15),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_15),
.B(n_250),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_15),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_15),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_15),
.B(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_16),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_16),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_16),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_16),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_17),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_17),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_17),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_17),
.B(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_17),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_17),
.B(n_129),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_496),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_487),
.Y(n_22)
);

NAND3xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_266),
.C(n_394),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_237),
.Y(n_24)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_25),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_195),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_26),
.B(n_195),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_116),
.B2(n_194),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_27),
.B(n_481),
.C(n_482),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

MAJx2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_75),
.C(n_93),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_29),
.B(n_197),
.Y(n_196)
);

AO21x1_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_57),
.B(n_74),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_42),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_42),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_31),
.B(n_42),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_32),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_32),
.Y(n_169)
);

OAI211xp5_ASAP7_75t_L g175 ( 
.A1(n_32),
.A2(n_170),
.B(n_173),
.C(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_32),
.B(n_170),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_32),
.B(n_171),
.C(n_174),
.Y(n_406)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_35),
.Y(n_126)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_35),
.Y(n_356)
);

XNOR2x1_ASAP7_75t_L g246 ( 
.A(n_36),
.B(n_169),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_37),
.B(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_37),
.B(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_41),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_41),
.Y(n_413)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_41),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.C(n_52),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_43),
.A2(n_46),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

CKINVDCx11_ASAP7_75t_R g245 ( 
.A(n_43),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_43),
.A2(n_245),
.B1(n_474),
.B2(n_475),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_43),
.A2(n_245),
.B1(n_526),
.B2(n_532),
.Y(n_525)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_45),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_45),
.Y(n_349)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_46),
.Y(n_244)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_50),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2x1_ASAP7_75t_SL g242 ( 
.A(n_52),
.B(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_55),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_57),
.B(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_71),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_59),
.B(n_69),
.C(n_71),
.Y(n_150)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_64),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_64),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_65),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_65),
.A2(n_69),
.B1(n_524),
.B2(n_525),
.Y(n_523)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_75),
.B(n_93),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_87),
.B2(n_92),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_79),
.B(n_82),
.C(n_88),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_79),
.B(n_204),
.Y(n_203)
);

XOR2x2_ASAP7_75t_L g287 ( 
.A(n_79),
.B(n_288),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_80),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_84),
.Y(n_477)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_89),
.Y(n_280)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_91),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_91),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_108),
.B2(n_115),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_153),
.C(n_154),
.Y(n_152)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_110),
.B(n_307),
.Y(n_306)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_115),
.A2(n_222),
.B(n_225),
.Y(n_221)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_116),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_165),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_117),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_151),
.Y(n_117)
);

INVxp33_ASAP7_75t_SL g436 ( 
.A(n_118),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_137),
.C(n_150),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_119),
.B(n_137),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_127),
.Y(n_119)
);

NOR2xp67_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_L g192 ( 
.A(n_121),
.B(n_123),
.C(n_136),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_121),
.A2(n_123),
.B(n_136),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_122),
.B(n_223),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_122),
.B(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_122),
.B(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_122),
.B(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_127)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_132),
.A2(n_136),
.B1(n_463),
.B2(n_465),
.Y(n_462)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_134),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_135),
.A2(n_192),
.B(n_193),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_136),
.B(n_463),
.C(n_466),
.Y(n_534)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_146),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_138),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_232)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_141),
.B(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_142),
.B(n_171),
.C(n_433),
.Y(n_453)
);

OR2x2_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_143),
.Y(n_298)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_144),
.Y(n_324)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_146),
.Y(n_231)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_148),
.Y(n_434)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_148),
.Y(n_531)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_150),
.Y(n_235)
);

XNOR2x1_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_152),
.Y(n_437)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_155),
.Y(n_438)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_164),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_157),
.Y(n_404)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_162),
.B(n_403),
.C(n_404),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_164),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_165),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_177),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_167),
.B(n_191),
.C(n_400),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_173),
.B(n_175),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2x2_ASAP7_75t_L g311 ( 
.A(n_171),
.B(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_171),
.B(n_433),
.Y(n_432)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_173),
.A2(n_174),
.B1(n_506),
.B2(n_511),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_191),
.Y(n_177)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_178),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_179),
.Y(n_420)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_190),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_184),
.Y(n_421)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g419 ( 
.A(n_190),
.B(n_420),
.C(n_421),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.C(n_233),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_196),
.B(n_265),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_199),
.B(n_234),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_221),
.C(n_229),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.C(n_214),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_202),
.A2(n_203),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_204),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_204),
.B(n_428),
.C(n_471),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_204),
.A2(n_288),
.B1(n_476),
.B2(n_478),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_204),
.B(n_245),
.C(n_478),
.Y(n_535)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_208),
.A2(n_209),
.B1(n_215),
.B2(n_216),
.Y(n_380)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_213),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_230),
.Y(n_240)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

INVxp33_ASAP7_75t_SL g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_264),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_238),
.B(n_264),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.C(n_261),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_239),
.B(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_241),
.A2(n_262),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_241),
.Y(n_389)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.C(n_247),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_242),
.B(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_246),
.A2(n_247),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_246),
.Y(n_373)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_247),
.Y(n_372)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.C(n_256),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_249),
.B1(n_256),
.B2(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_262),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_384),
.B(n_393),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_367),
.B(n_383),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_313),
.B(n_366),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_299),
.C(n_300),
.Y(n_270)
);

AOI21xp33_ASAP7_75t_SL g366 ( 
.A1(n_271),
.A2(n_299),
.B(n_300),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_285),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp33_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_286),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_274),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_276),
.B(n_285),
.C(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_281),
.C(n_282),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_277),
.A2(n_278),
.B1(n_281),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_281),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_283),
.B(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_287),
.B(n_295),
.C(n_377),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_R g392 ( 
.A(n_287),
.B(n_295),
.C(n_377),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_288),
.B(n_423),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_295),
.B2(n_296),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_304),
.C(n_311),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_301),
.B(n_330),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_304),
.A2(n_305),
.B1(n_311),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_308),
.B1(n_309),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_332),
.B(n_365),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_329),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_329),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.C(n_325),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_316),
.A2(n_317),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_320),
.B(n_325),
.Y(n_361)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_327),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_359),
.B(n_364),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_344),
.B(n_358),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_350),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_350),
.Y(n_358)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_353),
.B1(n_354),
.B2(n_357),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_351),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_357),
.Y(n_363)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_360),
.B(n_363),
.Y(n_364)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_361),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_381),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_381),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_370),
.B1(n_374),
.B2(n_375),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_391),
.C(n_392),
.Y(n_390)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_378),
.Y(n_391)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_390),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_386),
.B(n_390),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_394),
.A2(n_488),
.B(n_492),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_440),
.B1(n_479),
.B2(n_483),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_396),
.B(n_441),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_396),
.B(n_441),
.Y(n_495)
);

OAI22x1_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_416),
.B1(n_435),
.B2(n_439),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_398),
.B(n_417),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_401),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_399),
.B(n_456),
.C(n_457),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_405),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_402),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_405),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_SL g447 ( 
.A1(n_406),
.A2(n_412),
.B(n_414),
.C(n_448),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_412),
.B1(n_414),
.B2(n_415),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_408),
.B(n_415),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_409),
.B(n_410),
.Y(n_414)
);

NOR2x1_ASAP7_75t_R g512 ( 
.A(n_409),
.B(n_513),
.Y(n_512)
);

INVx5_ASAP7_75t_SL g410 ( 
.A(n_411),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_412),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_412),
.A2(n_415),
.B1(n_451),
.B2(n_452),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_413),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_415),
.B(n_452),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_415),
.B(n_452),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_435),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_417),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_431),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_422),
.Y(n_418)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_419),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g444 ( 
.A(n_422),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_428),
.Y(n_423)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_424),
.Y(n_471)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_444),
.C(n_445),
.Y(n_443)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_435),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.C(n_438),
.Y(n_435)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_454),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_442),
.B(n_537),
.C(n_538),
.Y(n_536)
);

XOR2x1_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_446),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_443),
.B(n_447),
.C(n_449),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_449),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_453),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g517 ( 
.A1(n_453),
.A2(n_518),
.B(n_519),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_458),
.Y(n_454)
);

INVxp33_ASAP7_75t_SL g537 ( 
.A(n_455),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_458),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_472),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_461),
.B1(n_469),
.B2(n_470),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_461),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_461),
.B(n_469),
.C(n_473),
.Y(n_521)
);

XOR2x2_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_466),
.Y(n_461)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_463),
.Y(n_465)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_476),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_484),
.Y(n_494)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_489),
.A2(n_490),
.B(n_491),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_494),
.B(n_495),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_539),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_536),
.Y(n_497)
);

NOR2xp67_ASAP7_75t_L g540 ( 
.A(n_498),
.B(n_536),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_522),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_520),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_516),
.B2(n_517),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

XOR2x1_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_512),
.Y(n_504)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_506),
.Y(n_511)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx8_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_533),
.Y(n_522)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_526),
.Y(n_532)
);

NAND2x1_ASAP7_75t_SL g526 ( 
.A(n_527),
.B(n_528),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_535),
.Y(n_533)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_540),
.Y(n_539)
);


endmodule