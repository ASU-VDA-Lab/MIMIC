module fake_jpeg_16445_n_89 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_89);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_89;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_22),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_16),
.A2(n_6),
.B1(n_9),
.B2(n_3),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_19),
.B1(n_2),
.B2(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_1),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_31),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_16),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_29),
.B1(n_16),
.B2(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_12),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_17),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_34),
.B(n_36),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_26),
.B1(n_24),
.B2(n_10),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_12),
.B(n_21),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_50),
.B(n_51),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_45),
.B1(n_26),
.B2(n_7),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_18),
.B1(n_17),
.B2(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx24_ASAP7_75t_SL g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_24),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_27),
.A2(n_18),
.B(n_6),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_4),
.C(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_56),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_57),
.B1(n_60),
.B2(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_64),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_9),
.B1(n_37),
.B2(n_43),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_42),
.B1(n_44),
.B2(n_50),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_51),
.B1(n_39),
.B2(n_48),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_67),
.Y(n_77)
);

INVxp33_ASAP7_75t_SL g67 ( 
.A(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_69),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_72),
.B1(n_57),
.B2(n_52),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_48),
.B(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_60),
.Y(n_74)
);

XNOR2x1_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_79),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_58),
.B(n_69),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

XNOR2x1_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_65),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_68),
.C(n_66),
.Y(n_81)
);

MAJx2_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_75),
.C(n_80),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_73),
.C(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_82),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_87),
.B1(n_82),
.B2(n_85),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);


endmodule