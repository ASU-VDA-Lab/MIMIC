module fake_jpeg_32192_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_42),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_14),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_21),
.B(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_55),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_51),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_77),
.A2(n_59),
.B1(n_52),
.B2(n_56),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_58),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_87),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_78),
.A2(n_68),
.B1(n_65),
.B2(n_72),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_92),
.B1(n_60),
.B2(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_65),
.B1(n_68),
.B2(n_71),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_55),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_68),
.B1(n_71),
.B2(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_69),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_64),
.B1(n_56),
.B2(n_62),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_64),
.B1(n_54),
.B2(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_58),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_96),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_70),
.B(n_66),
.C(n_57),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_109),
.B1(n_6),
.B2(n_9),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_103),
.Y(n_123)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_110),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_82),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_120),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_109),
.A2(n_81),
.B1(n_7),
.B2(n_8),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_50),
.B1(n_37),
.B2(n_38),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_95),
.C(n_96),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_100),
.C(n_97),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_34),
.Y(n_142)
);

NOR2x1p5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_10),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_19),
.B(n_22),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_11),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_17),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_11),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_12),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_130),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_118),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_135),
.B1(n_140),
.B2(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_13),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_133),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_118),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_138),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_127),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_124),
.B(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_123),
.B(n_121),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_143),
.A2(n_119),
.B1(n_126),
.B2(n_123),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_144),
.A2(n_41),
.B1(n_43),
.B2(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_148),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_149),
.Y(n_156)
);

AO22x1_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_122),
.B1(n_112),
.B2(n_46),
.Y(n_149)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_134),
.C(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_155),
.B(n_144),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_159),
.A2(n_160),
.B1(n_147),
.B2(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_151),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_152),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_153),
.C(n_158),
.Y(n_165)
);

AOI321xp33_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_150),
.A3(n_154),
.B1(n_156),
.B2(n_138),
.C(n_147),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_154),
.Y(n_167)
);


endmodule