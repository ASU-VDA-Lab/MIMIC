module fake_jpeg_1305_n_678 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_678);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_678;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_17),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_65),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_0),
.C(n_1),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_66),
.A2(n_57),
.B(n_27),
.C(n_29),
.Y(n_158)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_67),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_68),
.B(n_70),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_26),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_69),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_21),
.B(n_0),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_71),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_26),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_72),
.B(n_77),
.Y(n_134)
);

NAND2x1_ASAP7_75t_SL g73 ( 
.A(n_26),
.B(n_59),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_73),
.B(n_45),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_74),
.Y(n_223)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_75),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_76),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_32),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_32),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_78),
.B(n_79),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_32),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_81),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_82),
.Y(n_187)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_83),
.Y(n_176)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_85),
.Y(n_196)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_87),
.Y(n_200)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_88),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g214 ( 
.A(n_89),
.Y(n_214)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_90),
.Y(n_174)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_91),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g202 ( 
.A(n_92),
.B(n_119),
.Y(n_202)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_93),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_30),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_27),
.B(n_0),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_105),
.Y(n_149)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_100),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_28),
.B(n_1),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_106),
.Y(n_199)
);

BUFx12_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g173 ( 
.A(n_107),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_31),
.B(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_131),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_116),
.Y(n_146)
);

BUFx4f_ASAP7_75t_SL g111 ( 
.A(n_41),
.Y(n_111)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_41),
.Y(n_112)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_112),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_22),
.Y(n_115)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_33),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_123),
.Y(n_147)
);

BUFx12f_ASAP7_75t_SL g119 ( 
.A(n_44),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_31),
.Y(n_120)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_120),
.Y(n_204)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_23),
.Y(n_121)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_33),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_54),
.B(n_1),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_125),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_23),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_22),
.Y(n_126)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_126),
.Y(n_201)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_22),
.Y(n_128)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_128),
.Y(n_213)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_23),
.Y(n_129)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_129),
.Y(n_224)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_130),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_51),
.B(n_1),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_48),
.Y(n_132)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_133),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_81),
.A2(n_55),
.B1(n_40),
.B2(n_50),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_135),
.A2(n_165),
.B1(n_187),
.B2(n_214),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_66),
.A2(n_55),
.B1(n_57),
.B2(n_29),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_138),
.A2(n_152),
.B1(n_160),
.B2(n_184),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_90),
.A2(n_40),
.B1(n_45),
.B2(n_44),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_141),
.A2(n_161),
.B1(n_170),
.B2(n_186),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_52),
.B1(n_56),
.B2(n_53),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g288 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_73),
.B(n_45),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_82),
.A2(n_40),
.B1(n_56),
.B2(n_52),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_119),
.A2(n_45),
.B1(n_43),
.B2(n_37),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_91),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_75),
.A2(n_45),
.B1(n_43),
.B2(n_37),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_92),
.B(n_34),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_180),
.B(n_192),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_89),
.A2(n_34),
.B1(n_47),
.B2(n_41),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_101),
.A2(n_47),
.B1(n_41),
.B2(n_4),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_185),
.A2(n_209),
.B1(n_217),
.B2(n_220),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_75),
.A2(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_83),
.B(n_2),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_188),
.B(n_229),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_111),
.B(n_102),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_60),
.A2(n_47),
.B1(n_3),
.B2(n_6),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g269 ( 
.A1(n_195),
.A2(n_211),
.B1(n_141),
.B2(n_186),
.Y(n_269)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_86),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_198),
.Y(n_262)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_98),
.Y(n_207)
);

INVx3_ASAP7_75t_SL g294 ( 
.A(n_207),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_113),
.A2(n_47),
.B1(n_7),
.B2(n_8),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_64),
.A2(n_2),
.B1(n_7),
.B2(n_9),
.Y(n_211)
);

AO22x1_ASAP7_75t_L g212 ( 
.A1(n_121),
.A2(n_2),
.B1(n_7),
.B2(n_9),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_17),
.Y(n_252)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_215),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_114),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_122),
.B(n_10),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_219),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_61),
.A2(n_76),
.B1(n_74),
.B2(n_71),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_129),
.A2(n_12),
.B(n_14),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_221),
.B(n_228),
.Y(n_303)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_88),
.Y(n_222)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_67),
.Y(n_225)
);

BUFx4f_ASAP7_75t_SL g287 ( 
.A(n_225),
.Y(n_287)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_117),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_175),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_111),
.B(n_16),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_87),
.B(n_16),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_94),
.B(n_17),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_231),
.B(n_210),
.Y(n_277)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_232),
.Y(n_329)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_233),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_145),
.B(n_108),
.C(n_133),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_234),
.B(n_236),
.C(n_244),
.Y(n_334)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_235),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_149),
.B(n_132),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_237),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_238),
.Y(n_359)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_239),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_147),
.B(n_112),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_241),
.B(n_250),
.Y(n_357)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_156),
.B(n_112),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_245),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_177),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_246),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_SL g247 ( 
.A1(n_202),
.A2(n_107),
.B(n_126),
.C(n_115),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_SL g370 ( 
.A1(n_247),
.A2(n_269),
.B(n_272),
.C(n_285),
.Y(n_370)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_249),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_230),
.Y(n_250)
);

OAI22x1_ASAP7_75t_L g251 ( 
.A1(n_157),
.A2(n_102),
.B1(n_107),
.B2(n_128),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_251),
.A2(n_273),
.B1(n_293),
.B2(n_260),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_252),
.B(n_263),
.Y(n_340)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_134),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_254),
.B(n_256),
.Y(n_320)
);

BUFx12f_ASAP7_75t_L g255 ( 
.A(n_154),
.Y(n_255)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_255),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_166),
.B(n_18),
.Y(n_256)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_181),
.A2(n_18),
.B(n_19),
.C(n_97),
.D(n_158),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_257),
.A2(n_263),
.B(n_313),
.Y(n_354)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_174),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g350 ( 
.A(n_258),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_137),
.B(n_18),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_259),
.B(n_268),
.Y(n_325)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_187),
.Y(n_260)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_260),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_219),
.B(n_18),
.Y(n_263)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_159),
.Y(n_264)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_264),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_155),
.B(n_19),
.C(n_183),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_265),
.B(n_263),
.C(n_310),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_161),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_266),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_19),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_267),
.B(n_282),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_179),
.B(n_194),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g272 ( 
.A1(n_184),
.A2(n_217),
.B1(n_170),
.B2(n_160),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_144),
.A2(n_146),
.B1(n_135),
.B2(n_211),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_168),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_275),
.B(n_276),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_199),
.B(n_208),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_277),
.B(n_278),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_162),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_279),
.A2(n_295),
.B1(n_297),
.B2(n_251),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_204),
.B(n_150),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_280),
.B(n_284),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_151),
.Y(n_281)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_281),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_171),
.B(n_196),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_193),
.B(n_136),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_283),
.B(n_291),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_168),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_214),
.Y(n_285)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_148),
.B(n_164),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_286),
.B(n_289),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_172),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_143),
.Y(n_290)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_143),
.B(n_153),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_153),
.Y(n_292)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_195),
.A2(n_189),
.B1(n_178),
.B2(n_223),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_205),
.A2(n_140),
.B1(n_223),
.B2(n_216),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_189),
.B(n_178),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_296),
.B(n_300),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_163),
.A2(n_213),
.B1(n_201),
.B2(n_200),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_142),
.Y(n_298)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_298),
.Y(n_336)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_159),
.Y(n_299)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_299),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_190),
.B(n_191),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_142),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_301),
.B(n_314),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_140),
.B(n_216),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_302),
.B(n_312),
.Y(n_365)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_191),
.Y(n_304)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_139),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_305),
.Y(n_333)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_218),
.Y(n_306)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_306),
.Y(n_347)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_218),
.Y(n_307)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_307),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_206),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_308),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_163),
.B(n_201),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_310),
.B(n_315),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_226),
.B(n_200),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_311),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_167),
.B(n_213),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_159),
.B(n_169),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_313),
.B(n_245),
.Y(n_368)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_167),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_169),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_245),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_236),
.B(n_169),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_316),
.B(n_339),
.C(n_343),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_266),
.A2(n_279),
.B1(n_267),
.B2(n_288),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_318),
.A2(n_321),
.B1(n_331),
.B2(n_352),
.Y(n_381)
);

OAI22xp33_ASAP7_75t_L g321 ( 
.A1(n_272),
.A2(n_283),
.B1(n_242),
.B2(n_309),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_252),
.A2(n_270),
.B1(n_261),
.B2(n_272),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_271),
.B(n_244),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_257),
.A2(n_303),
.B(n_252),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_342),
.B(n_373),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_244),
.B(n_282),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_272),
.A2(n_247),
.B1(n_296),
.B2(n_302),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_344),
.A2(n_367),
.B1(n_370),
.B2(n_376),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_345),
.A2(n_299),
.B1(n_377),
.B2(n_370),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_349),
.B(n_238),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_242),
.A2(n_269),
.B1(n_291),
.B2(n_293),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_354),
.Y(n_401)
);

OA22x2_ASAP7_75t_L g358 ( 
.A1(n_242),
.A2(n_269),
.B1(n_243),
.B2(n_304),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_358),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_366),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_242),
.A2(n_269),
.B1(n_239),
.B2(n_234),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_368),
.B(n_340),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_265),
.B(n_240),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_245),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_375),
.A2(n_314),
.B1(n_262),
.B2(n_274),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_305),
.A2(n_308),
.B1(n_290),
.B2(n_243),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_248),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_378),
.B(n_383),
.C(n_395),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_338),
.Y(n_380)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_380),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_355),
.B(n_249),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_382),
.B(n_386),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_316),
.B(n_334),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_328),
.Y(n_384)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_385),
.B(n_415),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_363),
.B(n_253),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_353),
.Y(n_387)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_387),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_341),
.B(n_232),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_388),
.B(n_394),
.Y(n_457)
);

BUFx12_ASAP7_75t_L g389 ( 
.A(n_335),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_389),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_320),
.B(n_233),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_392),
.B(n_393),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_372),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_341),
.B(n_351),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_334),
.B(n_235),
.C(n_246),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_321),
.A2(n_292),
.B1(n_306),
.B2(n_307),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_396),
.A2(n_403),
.B1(n_405),
.B2(n_409),
.Y(n_434)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_335),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_397),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_326),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_398),
.B(n_400),
.Y(n_459)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_399),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_351),
.B(n_287),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_366),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_402),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_364),
.B(n_287),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_404),
.B(n_408),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_375),
.A2(n_352),
.B1(n_331),
.B2(n_367),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_L g406 ( 
.A(n_318),
.B(n_262),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_406),
.A2(n_333),
.B(n_361),
.Y(n_450)
);

AND2x2_ASAP7_75t_SL g407 ( 
.A(n_364),
.B(n_274),
.Y(n_407)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_407),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_287),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_370),
.A2(n_294),
.B1(n_278),
.B2(n_298),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_327),
.B(n_294),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_410),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_371),
.B(n_281),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_411),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_377),
.A2(n_258),
.B(n_255),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_413),
.A2(n_391),
.B(n_362),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_343),
.B(n_255),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_419),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_365),
.B(n_255),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_416),
.B(n_422),
.C(n_323),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_353),
.Y(n_417)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_417),
.Y(n_444)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_338),
.Y(n_418)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_418),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_349),
.B(n_264),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_421),
.A2(n_358),
.B(n_354),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_373),
.B(n_368),
.C(n_358),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_340),
.B(n_337),
.Y(n_423)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_423),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_357),
.B(n_374),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_424),
.Y(n_441)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_425),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_366),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_426),
.Y(n_454)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_319),
.Y(n_427)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_427),
.Y(n_466)
);

OA21x2_ASAP7_75t_L g437 ( 
.A1(n_381),
.A2(n_358),
.B(n_370),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_437),
.A2(n_442),
.B(n_449),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_439),
.Y(n_472)
);

NAND2x1_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_340),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_448),
.A2(n_406),
.B(n_413),
.Y(n_500)
);

OA21x2_ASAP7_75t_L g449 ( 
.A1(n_381),
.A2(n_342),
.B(n_376),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_450),
.A2(n_468),
.B(n_393),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_405),
.A2(n_325),
.B1(n_336),
.B2(n_322),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_452),
.A2(n_463),
.B1(n_387),
.B2(n_427),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_412),
.A2(n_353),
.B1(n_324),
.B2(n_369),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_456),
.A2(n_461),
.B1(n_465),
.B2(n_417),
.Y(n_483)
);

OAI32xp33_ASAP7_75t_L g460 ( 
.A1(n_394),
.A2(n_346),
.A3(n_360),
.B1(n_347),
.B2(n_332),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_454),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_412),
.A2(n_369),
.B1(n_356),
.B2(n_329),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_400),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_462),
.B(n_467),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_379),
.A2(n_317),
.B1(n_348),
.B2(n_329),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_379),
.A2(n_356),
.B1(n_317),
.B2(n_348),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_404),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_SL g468 ( 
.A1(n_409),
.A2(n_396),
.B1(n_391),
.B2(n_426),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_469),
.B(n_419),
.C(n_383),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_441),
.B(n_398),
.Y(n_470)
);

CKINVDCx14_ASAP7_75t_R g517 ( 
.A(n_470),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_459),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_471),
.B(n_474),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_473),
.B(n_480),
.C(n_486),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_459),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_445),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_475),
.B(n_478),
.Y(n_527)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_431),
.Y(n_476)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_476),
.Y(n_514)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_431),
.Y(n_477)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_477),
.Y(n_525)
);

NOR2x1_ASAP7_75t_L g478 ( 
.A(n_450),
.B(n_414),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_433),
.A2(n_423),
.B1(n_408),
.B2(n_415),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_479),
.A2(n_483),
.B1(n_487),
.B2(n_505),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_458),
.B(n_395),
.C(n_378),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_466),
.Y(n_481)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_481),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_441),
.B(n_411),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_482),
.B(n_488),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_390),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_484),
.B(n_453),
.Y(n_532)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_466),
.Y(n_485)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_485),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_432),
.B(n_420),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_437),
.A2(n_385),
.B1(n_388),
.B2(n_401),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_443),
.B(n_410),
.Y(n_488)
);

AO21x1_ASAP7_75t_L g533 ( 
.A1(n_490),
.A2(n_504),
.B(n_489),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_491),
.B(n_494),
.Y(n_535)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_438),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_492),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_390),
.C(n_420),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_493),
.B(n_444),
.C(n_453),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_462),
.A2(n_420),
.B1(n_407),
.B2(n_425),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_438),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_495),
.B(n_497),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_443),
.B(n_429),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_496),
.B(n_499),
.Y(n_518)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_460),
.Y(n_497)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_451),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_500),
.B(n_464),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_430),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_501),
.B(n_502),
.Y(n_528)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_451),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_435),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_503),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_457),
.B(n_407),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_437),
.A2(n_407),
.B1(n_384),
.B2(n_418),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_464),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_506),
.B(n_429),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_507),
.A2(n_439),
.B(n_442),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_449),
.A2(n_399),
.B1(n_380),
.B2(n_397),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_508),
.A2(n_434),
.B1(n_463),
.B2(n_467),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_484),
.B(n_448),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_509),
.B(n_516),
.Y(n_553)
);

XNOR2x1_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_432),
.Y(n_510)
);

XNOR2x1_ASAP7_75t_L g550 ( 
.A(n_510),
.B(n_521),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_473),
.B(n_448),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_SL g555 ( 
.A(n_512),
.B(n_519),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_513),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_480),
.B(n_435),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_493),
.B(n_455),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_497),
.A2(n_474),
.B1(n_471),
.B2(n_490),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_520),
.A2(n_505),
.B1(n_491),
.B2(n_500),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_472),
.A2(n_440),
.B(n_454),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_522),
.B(n_456),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_494),
.B(n_455),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_530),
.B(n_531),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_506),
.B(n_457),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_532),
.B(n_539),
.C(n_543),
.Y(n_554)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_533),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_487),
.B(n_489),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_534),
.B(n_538),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_536),
.A2(n_434),
.B1(n_483),
.B2(n_508),
.Y(n_552)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_537),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_504),
.B(n_449),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_478),
.B(n_444),
.C(n_440),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_475),
.B(n_433),
.Y(n_544)
);

NAND3xp33_ASAP7_75t_L g557 ( 
.A(n_544),
.B(n_511),
.C(n_527),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_501),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_545),
.B(n_481),
.Y(n_565)
);

CKINVDCx14_ASAP7_75t_R g546 ( 
.A(n_518),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_546),
.B(n_549),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_547),
.A2(n_530),
.B1(n_524),
.B2(n_502),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_542),
.A2(n_535),
.B1(n_523),
.B2(n_527),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_548),
.A2(n_552),
.B1(n_574),
.B2(n_515),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_517),
.B(n_452),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_523),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_556),
.B(n_557),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_528),
.B(n_492),
.Y(n_558)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_558),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_526),
.B(n_478),
.C(n_507),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_561),
.B(n_568),
.C(n_571),
.Y(n_577)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_529),
.Y(n_562)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_562),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_542),
.A2(n_428),
.B1(n_472),
.B2(n_485),
.Y(n_563)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_563),
.Y(n_598)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_529),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_564),
.B(n_569),
.Y(n_590)
);

CKINVDCx14_ASAP7_75t_R g579 ( 
.A(n_565),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_520),
.B(n_495),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_566),
.B(n_570),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_526),
.B(n_447),
.C(n_498),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_533),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_531),
.B(n_476),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_516),
.B(n_447),
.C(n_498),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_572),
.A2(n_446),
.B(n_380),
.Y(n_599)
);

CKINVDCx16_ASAP7_75t_R g573 ( 
.A(n_522),
.Y(n_573)
);

INVx8_ASAP7_75t_L g600 ( 
.A(n_573),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_535),
.A2(n_428),
.B1(n_477),
.B2(n_461),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_514),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_575),
.A2(n_541),
.B(n_525),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_578),
.A2(n_582),
.B1(n_585),
.B2(n_567),
.Y(n_617)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_581),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_548),
.A2(n_534),
.B1(n_538),
.B2(n_540),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_568),
.B(n_539),
.C(n_532),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_583),
.B(n_591),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_553),
.B(n_509),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_584),
.B(n_589),
.C(n_595),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_556),
.A2(n_543),
.B1(n_521),
.B2(n_513),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_587),
.A2(n_572),
.B1(n_547),
.B2(n_574),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_553),
.B(n_510),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_554),
.B(n_512),
.C(n_519),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_571),
.B(n_524),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_593),
.B(n_597),
.C(n_587),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_554),
.B(n_430),
.C(n_499),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_561),
.B(n_576),
.C(n_555),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_596),
.B(n_597),
.C(n_601),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_550),
.B(n_465),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_599),
.A2(n_572),
.B(n_562),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_550),
.B(n_446),
.Y(n_601)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_602),
.Y(n_624)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_603),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_578),
.A2(n_559),
.B1(n_566),
.B2(n_551),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_606),
.A2(n_617),
.B1(n_362),
.B2(n_323),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_586),
.Y(n_608)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_608),
.Y(n_625)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_594),
.Y(n_609)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_609),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_595),
.B(n_576),
.C(n_551),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_611),
.B(n_613),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_579),
.B(n_560),
.Y(n_612)
);

AOI21xp33_ASAP7_75t_L g632 ( 
.A1(n_612),
.A2(n_619),
.B(n_580),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_588),
.B(n_560),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_583),
.B(n_555),
.C(n_564),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_614),
.B(n_616),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_590),
.A2(n_559),
.B(n_598),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_615),
.A2(n_612),
.B(n_619),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_593),
.B(n_558),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_577),
.B(n_584),
.C(n_591),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_618),
.B(n_620),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_592),
.B(n_570),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_577),
.B(n_596),
.C(n_589),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_585),
.A2(n_567),
.B1(n_572),
.B2(n_436),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_621),
.B(n_436),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_622),
.B(n_580),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_627),
.B(n_639),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_618),
.B(n_582),
.C(n_599),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_628),
.B(n_630),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_604),
.A2(n_600),
.B(n_581),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g650 ( 
.A(n_631),
.B(n_620),
.Y(n_650)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_632),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_611),
.B(n_601),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_633),
.B(n_634),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_622),
.B(n_600),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_636),
.A2(n_637),
.B1(n_625),
.B2(n_639),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_615),
.A2(n_389),
.B(n_359),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_608),
.B(n_359),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_SL g649 ( 
.A(n_640),
.B(n_610),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_629),
.B(n_607),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_641),
.B(n_645),
.Y(n_656)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_623),
.A2(n_603),
.B(n_602),
.Y(n_644)
);

AOI21x1_ASAP7_75t_L g658 ( 
.A1(n_644),
.A2(n_652),
.B(n_635),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_638),
.B(n_625),
.Y(n_645)
);

FAx1_ASAP7_75t_SL g648 ( 
.A(n_628),
.B(n_606),
.CI(n_614),
.CON(n_648),
.SN(n_648)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_648),
.B(n_650),
.Y(n_663)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_649),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_651),
.Y(n_661)
);

NAND3xp33_ASAP7_75t_L g652 ( 
.A(n_627),
.B(n_610),
.C(n_605),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_637),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_653),
.B(n_654),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_634),
.B(n_605),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_SL g655 ( 
.A1(n_642),
.A2(n_626),
.B(n_624),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_655),
.A2(n_648),
.B(n_389),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_643),
.B(n_631),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_657),
.B(n_658),
.C(n_664),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_650),
.B(n_633),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_659),
.Y(n_666)
);

AO21x2_ASAP7_75t_L g662 ( 
.A1(n_651),
.A2(n_389),
.B(n_350),
.Y(n_662)
);

AO21x1_ASAP7_75t_L g665 ( 
.A1(n_662),
.A2(n_647),
.B(n_646),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_665),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_663),
.A2(n_652),
.B(n_647),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_667),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_656),
.Y(n_668)
);

AOI311xp33_ASAP7_75t_L g673 ( 
.A1(n_668),
.A2(n_669),
.A3(n_670),
.B(n_660),
.C(n_661),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_673),
.A2(n_672),
.B(n_671),
.Y(n_674)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_674),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_672),
.A2(n_657),
.B(n_666),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_676),
.A2(n_675),
.B(n_662),
.Y(n_677)
);

HAxp5_ASAP7_75t_SL g678 ( 
.A(n_677),
.B(n_662),
.CON(n_678),
.SN(n_678)
);


endmodule