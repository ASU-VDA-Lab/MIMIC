module fake_jpeg_31308_n_109 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_109);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_109;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVxp33_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_15),
.C(n_32),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_47),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_14),
.B(n_30),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_54),
.B1(n_37),
.B2(n_39),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_16),
.B(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_49),
.B(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_52),
.Y(n_58)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_44),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_65),
.B1(n_45),
.B2(n_5),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_11),
.B(n_12),
.Y(n_80)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_20),
.Y(n_74)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_41),
.B1(n_36),
.B2(n_45),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_79),
.B(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_3),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_6),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_59),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_25),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_6),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_78),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_21),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_55),
.B(n_18),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_91),
.B(n_92),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_28),
.B1(n_91),
.B2(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_89),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_34),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_26),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_86),
.C(n_85),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_85),
.B(n_87),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_98),
.C(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_99),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_101),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_108),
.A2(n_97),
.B(n_96),
.Y(n_109)
);


endmodule