module fake_jpeg_27807_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx2_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_4),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_0),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_0),
.B(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_11),
.B(n_0),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_15),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_18),
.B1(n_13),
.B2(n_19),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_25),
.B1(n_18),
.B2(n_13),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_22),
.B(n_21),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_25),
.B(n_21),
.C(n_30),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_22),
.C(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_27),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_5),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_39),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_20),
.B1(n_16),
.B2(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_44),
.B1(n_38),
.B2(n_20),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_34),
.C(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_27),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_54),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_55),
.C(n_56),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_16),
.C(n_8),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_60),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_49),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_7),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_61),
.B(n_7),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_57),
.B(n_8),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_9),
.C(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_69),
.Y(n_71)
);

BUFx24_ASAP7_75t_SL g72 ( 
.A(n_71),
.Y(n_72)
);


endmodule