module fake_netlist_1_4879_n_380 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_3, n_18, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_380);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_3;
input n_18;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_380;
wire n_117;
wire n_361;
wire n_185;
wire n_57;
wire n_284;
wire n_278;
wire n_60;
wire n_114;
wire n_94;
wire n_125;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_163;
wire n_105;
wire n_227;
wire n_231;
wire n_298;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_100;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_62;
wire n_255;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_247;
wire n_304;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_243;
wire n_235;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_59;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_61;
wire n_259;
wire n_308;
wire n_93;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_88;
wire n_107;
wire n_254;
wire n_262;
wire n_239;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_342;
wire n_370;
wire n_217;
wire n_139;
wire n_193;
wire n_273;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_374;
wire n_111;
wire n_64;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_168;
wire n_134;
wire n_233;
wire n_82;
wire n_106;
wire n_173;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_63;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_356;
wire n_281;
wire n_341;
wire n_58;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_159;
wire n_337;
wire n_176;
wire n_68;
wire n_123;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_332;
wire n_350;
wire n_164;
wire n_175;
wire n_145;
wire n_290;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_151;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g57 ( .A(n_55), .Y(n_57) );
INVx1_ASAP7_75t_L g58 ( .A(n_6), .Y(n_58) );
CKINVDCx20_ASAP7_75t_R g59 ( .A(n_14), .Y(n_59) );
INVx1_ASAP7_75t_L g60 ( .A(n_2), .Y(n_60) );
CKINVDCx16_ASAP7_75t_R g61 ( .A(n_13), .Y(n_61) );
INVx1_ASAP7_75t_L g62 ( .A(n_10), .Y(n_62) );
INVx1_ASAP7_75t_L g63 ( .A(n_3), .Y(n_63) );
INVx1_ASAP7_75t_L g64 ( .A(n_49), .Y(n_64) );
INVx2_ASAP7_75t_L g65 ( .A(n_27), .Y(n_65) );
INVxp67_ASAP7_75t_SL g66 ( .A(n_52), .Y(n_66) );
INVx1_ASAP7_75t_L g67 ( .A(n_41), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_28), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_37), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_29), .Y(n_70) );
INVxp33_ASAP7_75t_L g71 ( .A(n_38), .Y(n_71) );
INVxp67_ASAP7_75t_L g72 ( .A(n_40), .Y(n_72) );
CKINVDCx5p33_ASAP7_75t_R g73 ( .A(n_51), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_14), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_18), .Y(n_75) );
INVxp33_ASAP7_75t_SL g76 ( .A(n_47), .Y(n_76) );
INVxp33_ASAP7_75t_SL g77 ( .A(n_21), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_56), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_33), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_17), .Y(n_80) );
INVxp33_ASAP7_75t_L g81 ( .A(n_50), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_22), .Y(n_82) );
CKINVDCx14_ASAP7_75t_R g83 ( .A(n_23), .Y(n_83) );
NOR2xp67_ASAP7_75t_L g84 ( .A(n_42), .B(n_39), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_35), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_45), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_48), .Y(n_87) );
BUFx6f_ASAP7_75t_SL g88 ( .A(n_46), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_12), .Y(n_89) );
INVxp33_ASAP7_75t_SL g90 ( .A(n_8), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_31), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_65), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_57), .Y(n_93) );
NOR2xp33_ASAP7_75t_L g94 ( .A(n_90), .B(n_0), .Y(n_94) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_65), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g96 ( .A(n_58), .B(n_60), .Y(n_96) );
INVx3_ASAP7_75t_L g97 ( .A(n_91), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_57), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_64), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_61), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_58), .B(n_0), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_64), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_83), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_67), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_76), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_60), .B(n_1), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_67), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_68), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_68), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_69), .Y(n_110) );
NOR2xp33_ASAP7_75t_R g111 ( .A(n_73), .B(n_26), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_69), .Y(n_112) );
INVx3_ASAP7_75t_L g113 ( .A(n_70), .Y(n_113) );
INVx5_ASAP7_75t_L g114 ( .A(n_88), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_70), .Y(n_115) );
INVx4_ASAP7_75t_L g116 ( .A(n_114), .Y(n_116) );
INVx5_ASAP7_75t_L g117 ( .A(n_114), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_108), .Y(n_118) );
NAND3x1_ASAP7_75t_L g119 ( .A(n_96), .B(n_91), .C(n_78), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g120 ( .A(n_114), .B(n_78), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_108), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_108), .Y(n_122) );
INVxp33_ASAP7_75t_L g123 ( .A(n_94), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_93), .A2(n_62), .B1(n_63), .B2(n_80), .Y(n_124) );
AOI21x1_ASAP7_75t_L g125 ( .A1(n_93), .A2(n_79), .B(n_82), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_114), .B(n_71), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_108), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_108), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_95), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_97), .B(n_62), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_95), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_108), .Y(n_133) );
NAND3xp33_ASAP7_75t_L g134 ( .A(n_98), .B(n_79), .C(n_82), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_108), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_95), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_112), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_112), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_97), .B(n_85), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_95), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_131), .B(n_99), .Y(n_141) );
NOR2xp33_ASAP7_75t_R g142 ( .A(n_125), .B(n_100), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_139), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_132), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
NOR2xp33_ASAP7_75t_R g146 ( .A(n_125), .B(n_103), .Y(n_146) );
NOR3xp33_ASAP7_75t_SL g147 ( .A(n_134), .B(n_105), .C(n_106), .Y(n_147) );
BUFx4f_ASAP7_75t_L g148 ( .A(n_139), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_130), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_130), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_130), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_132), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_139), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_131), .A2(n_99), .B1(n_109), .B2(n_106), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_130), .B(n_97), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_126), .B(n_97), .Y(n_156) );
INVx2_ASAP7_75t_SL g157 ( .A(n_130), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_139), .Y(n_158) );
OR2x2_ASAP7_75t_L g159 ( .A(n_123), .B(n_96), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_126), .B(n_113), .Y(n_160) );
NOR3xp33_ASAP7_75t_SL g161 ( .A(n_134), .B(n_101), .C(n_75), .Y(n_161) );
BUFx2_ASAP7_75t_L g162 ( .A(n_139), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_139), .Y(n_163) );
NOR3xp33_ASAP7_75t_SL g164 ( .A(n_120), .B(n_101), .C(n_74), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_124), .B(n_114), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_139), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_139), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_132), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_119), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_124), .B(n_113), .Y(n_171) );
AOI221xp5_ASAP7_75t_L g172 ( .A1(n_120), .A2(n_89), .B1(n_80), .B2(n_63), .C(n_107), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_119), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_119), .B(n_113), .Y(n_174) );
INVxp67_ASAP7_75t_L g175 ( .A(n_159), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_159), .B(n_113), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_157), .A2(n_59), .B1(n_81), .B2(n_77), .Y(n_177) );
AOI221xp5_ASAP7_75t_L g178 ( .A1(n_149), .A2(n_89), .B1(n_110), .B2(n_107), .C(n_102), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_143), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_174), .A2(n_102), .B1(n_110), .B2(n_107), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_150), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_155), .B(n_102), .Y(n_182) );
CKINVDCx11_ASAP7_75t_R g183 ( .A(n_143), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_142), .Y(n_184) );
AOI21xp33_ASAP7_75t_L g185 ( .A1(n_169), .A2(n_72), .B(n_66), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_157), .A2(n_110), .B1(n_104), .B2(n_88), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_154), .B(n_104), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_174), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_151), .B(n_86), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_144), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_155), .B(n_104), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_174), .A2(n_88), .B1(n_87), .B2(n_85), .Y(n_192) );
BUFx12f_ASAP7_75t_L g193 ( .A(n_143), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_144), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_141), .B(n_92), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_158), .A2(n_92), .B1(n_112), .B2(n_115), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_173), .A2(n_112), .B1(n_115), .B2(n_84), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_162), .B(n_112), .Y(n_198) );
BUFx12f_ASAP7_75t_L g199 ( .A(n_143), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_162), .Y(n_200) );
NAND2x1p5_ASAP7_75t_L g201 ( .A(n_148), .B(n_117), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_161), .B(n_171), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_143), .B(n_112), .Y(n_203) );
INVx3_ASAP7_75t_SL g204 ( .A(n_158), .Y(n_204) );
OR2x6_ASAP7_75t_L g205 ( .A(n_145), .B(n_116), .Y(n_205) );
AOI221x1_ASAP7_75t_L g206 ( .A1(n_156), .A2(n_95), .B1(n_112), .B2(n_115), .C(n_140), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_145), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_193), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_202), .A2(n_160), .B(n_165), .Y(n_209) );
BUFx4f_ASAP7_75t_L g210 ( .A(n_193), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_175), .B(n_148), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_190), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_182), .B(n_148), .Y(n_213) );
AOI22xp33_ASAP7_75t_SL g214 ( .A1(n_177), .A2(n_146), .B1(n_115), .B2(n_166), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_183), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_182), .A2(n_172), .B1(n_115), .B2(n_95), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_188), .B(n_145), .Y(n_217) );
OAI211xp5_ASAP7_75t_SL g218 ( .A1(n_176), .A2(n_147), .B(n_164), .C(n_135), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_199), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_199), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_181), .B(n_145), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_184), .B(n_166), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_180), .A2(n_167), .B1(n_115), .B2(n_153), .Y(n_223) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_206), .A2(n_136), .B(n_137), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_181), .A2(n_115), .B1(n_95), .B2(n_163), .Y(n_225) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_197), .A2(n_136), .B(n_137), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_195), .A2(n_152), .B(n_168), .Y(n_227) );
OR2x2_ASAP7_75t_L g228 ( .A(n_191), .B(n_187), .Y(n_228) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_206), .A2(n_136), .B(n_118), .Y(n_229) );
OR2x2_ASAP7_75t_L g230 ( .A(n_200), .B(n_163), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_200), .B(n_145), .Y(n_231) );
AO31x2_ASAP7_75t_L g232 ( .A1(n_196), .A2(n_118), .A3(n_121), .B(n_122), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_211), .B(n_228), .Y(n_233) );
AO31x2_ASAP7_75t_L g234 ( .A1(n_209), .A2(n_189), .A3(n_190), .B(n_194), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_212), .Y(n_235) );
AOI222xp33_ASAP7_75t_L g236 ( .A1(n_211), .A2(n_178), .B1(n_184), .B2(n_183), .C1(n_198), .C2(n_204), .Y(n_236) );
AOI21x1_ASAP7_75t_L g237 ( .A1(n_224), .A2(n_203), .B(n_127), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_228), .A2(n_192), .B1(n_186), .B2(n_204), .Y(n_238) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_229), .A2(n_121), .B(n_122), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_210), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_212), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_211), .A2(n_204), .B1(n_185), .B2(n_167), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_212), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_221), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_221), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_218), .A2(n_198), .B1(n_203), .B2(n_205), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_218), .A2(n_203), .B1(n_205), .B2(n_179), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_208), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_213), .A2(n_153), .B1(n_205), .B2(n_207), .Y(n_249) );
AOI221xp5_ASAP7_75t_L g250 ( .A1(n_209), .A2(n_111), .B1(n_135), .B2(n_127), .C(n_128), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_210), .Y(n_251) );
AOI221x1_ASAP7_75t_SL g252 ( .A1(n_248), .A2(n_1), .B1(n_2), .B2(n_3), .C(n_4), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_241), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_241), .B(n_221), .Y(n_254) );
NAND3xp33_ASAP7_75t_L g255 ( .A(n_236), .B(n_214), .C(n_247), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_245), .B(n_232), .Y(n_256) );
OR2x6_ASAP7_75t_L g257 ( .A(n_244), .B(n_231), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_233), .A2(n_214), .B1(n_215), .B2(n_210), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_243), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_238), .A2(n_215), .B1(n_213), .B2(n_208), .Y(n_260) );
NOR4xp25_ASAP7_75t_SL g261 ( .A(n_251), .B(n_219), .C(n_215), .D(n_232), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_235), .B(n_232), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_245), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_244), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_234), .B(n_232), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_237), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_240), .A2(n_215), .B1(n_220), .B2(n_230), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_240), .Y(n_268) );
OR2x6_ASAP7_75t_L g269 ( .A(n_259), .B(n_237), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_259), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_253), .Y(n_271) );
OAI31xp33_ASAP7_75t_L g272 ( .A1(n_258), .A2(n_220), .A3(n_223), .B(n_231), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_256), .B(n_234), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_253), .Y(n_274) );
OAI211xp5_ASAP7_75t_SL g275 ( .A1(n_260), .A2(n_242), .B(n_246), .C(n_216), .Y(n_275) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_262), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_263), .B(n_251), .Y(n_277) );
AOI221xp5_ASAP7_75t_SL g278 ( .A1(n_258), .A2(n_222), .B1(n_223), .B2(n_250), .C(n_225), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_266), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_262), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_265), .B(n_239), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_265), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_265), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_266), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_254), .B(n_231), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_266), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_254), .B(n_232), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_264), .B(n_239), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_257), .B(n_239), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g290 ( .A(n_255), .B(n_249), .C(n_225), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_280), .B(n_252), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_272), .B(n_267), .Y(n_292) );
INVx3_ASAP7_75t_SL g293 ( .A(n_269), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_282), .B(n_267), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_282), .B(n_257), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_276), .B(n_257), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_283), .B(n_257), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_271), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_283), .B(n_257), .Y(n_299) );
NAND2xp33_ASAP7_75t_SL g300 ( .A(n_274), .B(n_261), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_270), .B(n_268), .Y(n_301) );
NAND2xp33_ASAP7_75t_SL g302 ( .A(n_273), .B(n_268), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_277), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_288), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_273), .B(n_226), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_281), .B(n_226), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_285), .B(n_4), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_281), .B(n_226), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_279), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_287), .B(n_5), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_275), .B(n_6), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_289), .B(n_224), .Y(n_312) );
NOR3xp33_ASAP7_75t_L g313 ( .A(n_290), .B(n_128), .C(n_138), .Y(n_313) );
AOI221xp5_ASAP7_75t_L g314 ( .A1(n_311), .A2(n_278), .B1(n_289), .B2(n_284), .C(n_286), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_292), .A2(n_269), .B1(n_217), .B2(n_230), .Y(n_315) );
OAI21xp5_ASAP7_75t_L g316 ( .A1(n_313), .A2(n_227), .B(n_217), .Y(n_316) );
AOI21xp33_ASAP7_75t_SL g317 ( .A1(n_293), .A2(n_7), .B(n_9), .Y(n_317) );
AOI222xp33_ASAP7_75t_L g318 ( .A1(n_291), .A2(n_217), .B1(n_11), .B2(n_12), .C1(n_13), .C2(n_15), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_304), .B(n_15), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_307), .A2(n_224), .B1(n_229), .B2(n_140), .Y(n_320) );
OAI222xp33_ASAP7_75t_L g321 ( .A1(n_296), .A2(n_16), .B1(n_17), .B2(n_18), .C1(n_19), .C2(n_201), .Y(n_321) );
AOI21xp33_ASAP7_75t_SL g322 ( .A1(n_293), .A2(n_16), .B(n_19), .Y(n_322) );
NAND2x1_ASAP7_75t_L g323 ( .A(n_296), .B(n_207), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_299), .B(n_20), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_310), .A2(n_207), .B1(n_179), .B2(n_201), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_302), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_297), .A2(n_201), .B1(n_153), .B2(n_140), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_303), .B(n_24), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_298), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_301), .B(n_25), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_297), .A2(n_153), .B1(n_129), .B2(n_138), .Y(n_331) );
NAND3xp33_ASAP7_75t_L g332 ( .A(n_300), .B(n_129), .C(n_133), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_306), .B(n_308), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_295), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_312), .B(n_30), .Y(n_335) );
INVxp67_ASAP7_75t_L g336 ( .A(n_302), .Y(n_336) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_294), .A2(n_129), .B(n_153), .C(n_34), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g338 ( .A1(n_305), .A2(n_133), .B(n_32), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_333), .B(n_334), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_329), .Y(n_340) );
XNOR2x1_ASAP7_75t_L g341 ( .A(n_319), .B(n_305), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_314), .B(n_309), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_315), .B(n_36), .Y(n_343) );
NOR2xp33_ASAP7_75t_R g344 ( .A(n_326), .B(n_43), .Y(n_344) );
INVxp67_ASAP7_75t_L g345 ( .A(n_317), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_323), .Y(n_346) );
XOR2x2_ASAP7_75t_L g347 ( .A(n_332), .B(n_44), .Y(n_347) );
NOR2xp33_ASAP7_75t_SL g348 ( .A(n_321), .B(n_53), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_336), .B(n_54), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g350 ( .A1(n_345), .A2(n_318), .B1(n_322), .B2(n_338), .C(n_330), .Y(n_350) );
XNOR2xp5_ASAP7_75t_L g351 ( .A(n_341), .B(n_324), .Y(n_351) );
O2A1O1Ixp5_ASAP7_75t_L g352 ( .A1(n_342), .A2(n_325), .B(n_327), .C(n_335), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_348), .A2(n_325), .B1(n_327), .B2(n_320), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_341), .A2(n_328), .B1(n_331), .B2(n_337), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_340), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_344), .B(n_316), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_339), .B(n_170), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_347), .A2(n_116), .B1(n_117), .B2(n_346), .Y(n_358) );
INVxp33_ASAP7_75t_L g359 ( .A(n_344), .Y(n_359) );
NOR3xp33_ASAP7_75t_L g360 ( .A(n_352), .B(n_349), .C(n_343), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_357), .Y(n_361) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_351), .Y(n_362) );
XNOR2x1_ASAP7_75t_L g363 ( .A(n_358), .B(n_354), .Y(n_363) );
AOI211xp5_ASAP7_75t_L g364 ( .A1(n_359), .A2(n_353), .B(n_350), .C(n_356), .Y(n_364) );
NOR3xp33_ASAP7_75t_SL g365 ( .A(n_350), .B(n_353), .C(n_356), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_355), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_359), .A2(n_353), .B1(n_356), .B2(n_350), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_352), .A2(n_351), .B1(n_359), .B2(n_345), .C(n_350), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_362), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_365), .B(n_364), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_366), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_367), .B(n_363), .Y(n_372) );
NOR2x1p5_ASAP7_75t_L g373 ( .A(n_369), .B(n_361), .Y(n_373) );
XOR2x2_ASAP7_75t_L g374 ( .A(n_370), .B(n_368), .Y(n_374) );
AND2x2_ASAP7_75t_SL g375 ( .A(n_372), .B(n_360), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_373), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_373), .B(n_369), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_377), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_378), .A2(n_374), .B1(n_377), .B2(n_375), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_379), .A2(n_376), .B(n_371), .Y(n_380) );
endmodule