module fake_jpeg_12074_n_411 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_411);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_52),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_56),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

HAxp5_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_0),
.CON(n_57),
.SN(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_75),
.B(n_28),
.C(n_40),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_59),
.Y(n_90)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_64),
.Y(n_108)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_73),
.Y(n_109)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx9p33_ASAP7_75t_R g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_38),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_43),
.A2(n_0),
.B(n_1),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_80),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_82),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_84),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_24),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_124),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_93),
.B(n_52),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_26),
.B1(n_42),
.B2(n_35),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_94),
.A2(n_121),
.B1(n_84),
.B2(n_31),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_47),
.A2(n_26),
.B1(n_22),
.B2(n_29),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_104),
.A2(n_122),
.B1(n_74),
.B2(n_50),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_57),
.A2(n_37),
.B1(n_29),
.B2(n_40),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_66),
.A2(n_29),
.B1(n_41),
.B2(n_40),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_66),
.A2(n_28),
.B1(n_41),
.B2(n_21),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_49),
.B(n_42),
.C(n_27),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_31),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_63),
.A2(n_41),
.B1(n_21),
.B2(n_23),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_126),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_80),
.A2(n_36),
.B1(n_35),
.B2(n_27),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_54),
.A2(n_22),
.B1(n_28),
.B2(n_23),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_36),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_20),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_30),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_85),
.A2(n_51),
.B1(n_61),
.B2(n_23),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_124),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_132),
.B(n_134),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_133),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_30),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_77),
.B1(n_71),
.B2(n_58),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_135),
.A2(n_165),
.B1(n_99),
.B2(n_86),
.Y(n_188)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_120),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_111),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_139),
.B(n_140),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_64),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_142),
.B(n_144),
.Y(n_189)
);

INVx6_ASAP7_75t_SL g143 ( 
.A(n_98),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_143),
.Y(n_180)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_151),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_104),
.A2(n_83),
.B1(n_81),
.B2(n_60),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_155),
.B1(n_159),
.B2(n_166),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_82),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_88),
.A2(n_93),
.B(n_118),
.C(n_109),
.Y(n_152)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_152),
.B(n_127),
.CI(n_31),
.CON(n_174),
.SN(n_174)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_72),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_156),
.C(n_158),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_154),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_89),
.B(n_0),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_87),
.B(n_15),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_59),
.B1(n_78),
.B2(n_76),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_89),
.B(n_2),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_163),
.C(n_167),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_92),
.B(n_3),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_92),
.A2(n_67),
.B1(n_46),
.B2(n_68),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_101),
.B(n_3),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_106),
.B(n_12),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_117),
.B(n_90),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_137),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_184),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_164),
.A2(n_99),
.B1(n_91),
.B2(n_90),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_175),
.A2(n_154),
.B1(n_91),
.B2(n_96),
.Y(n_216)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_119),
.B1(n_101),
.B2(n_130),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_165),
.B1(n_142),
.B2(n_139),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_143),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_131),
.A2(n_130),
.B1(n_115),
.B2(n_116),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_196),
.B1(n_150),
.B2(n_166),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_151),
.Y(n_222)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_131),
.A2(n_116),
.B1(n_86),
.B2(n_95),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_209),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_186),
.B(n_132),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_201),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_152),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_161),
.B(n_149),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_203),
.A2(n_173),
.B(n_171),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_146),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_208),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_196),
.B1(n_188),
.B2(n_178),
.Y(n_232)
);

AO22x1_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_141),
.B1(n_159),
.B2(n_149),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_207),
.A2(n_211),
.B(n_217),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_146),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_195),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_140),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_212),
.B(n_168),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_158),
.C(n_146),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_214),
.C(n_163),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_144),
.Y(n_214)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_216),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_177),
.A2(n_167),
.B(n_156),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_195),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_199),
.B1(n_219),
.B2(n_209),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_181),
.B(n_134),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_223),
.B(n_160),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_243),
.B(n_171),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_187),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_230),
.B(n_239),
.C(n_249),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_232),
.A2(n_245),
.B1(n_190),
.B2(n_191),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_202),
.B(n_222),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_250),
.B(n_198),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_234),
.B(n_248),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_212),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_240),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_174),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_242),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_215),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_214),
.Y(n_242)
);

AO21x2_ASAP7_75t_L g244 ( 
.A1(n_207),
.A2(n_178),
.B(n_182),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_210),
.B1(n_218),
.B2(n_147),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_206),
.A2(n_180),
.B1(n_184),
.B2(n_194),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_180),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_237),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_201),
.C(n_208),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_202),
.A2(n_207),
.B(n_205),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_251),
.A2(n_269),
.B(n_278),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_259),
.Y(n_291)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_226),
.A2(n_221),
.B1(n_220),
.B2(n_198),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_257),
.A2(n_268),
.B1(n_270),
.B2(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_234),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_261),
.Y(n_303)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_235),
.Y(n_288)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_272),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_210),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_266),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_267),
.A2(n_271),
.B1(n_273),
.B2(n_197),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_226),
.A2(n_183),
.B1(n_193),
.B2(n_133),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_192),
.B(n_176),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_230),
.B1(n_233),
.B2(n_227),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_193),
.B1(n_133),
.B2(n_147),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_229),
.Y(n_274)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_193),
.B1(n_197),
.B2(n_119),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_229),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_227),
.B(n_157),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_243),
.A2(n_197),
.B(n_191),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_247),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_231),
.B1(n_250),
.B2(n_235),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_239),
.C(n_249),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_299),
.C(n_300),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_292),
.B1(n_296),
.B2(n_305),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_270),
.A2(n_244),
.B1(n_232),
.B2(n_231),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_302),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_255),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_244),
.B1(n_225),
.B2(n_242),
.Y(n_292)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_294),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_273),
.A2(n_241),
.B1(n_248),
.B2(n_119),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_306),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_254),
.B(n_241),
.C(n_172),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_172),
.C(n_97),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_97),
.C(n_145),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_272),
.C(n_265),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_275),
.A2(n_154),
.B1(n_95),
.B2(n_96),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_261),
.A2(n_102),
.B1(n_115),
.B2(n_128),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_252),
.B(n_102),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_284),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_315),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_283),
.B1(n_292),
.B2(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_312),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_291),
.Y(n_315)
);

AOI211xp5_ASAP7_75t_L g316 ( 
.A1(n_295),
.A2(n_276),
.B(n_269),
.C(n_279),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_316),
.A2(n_328),
.B1(n_289),
.B2(n_296),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_259),
.B1(n_263),
.B2(n_253),
.Y(n_317)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_252),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_318),
.B(n_321),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_300),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_266),
.C(n_251),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_299),
.C(n_306),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_324),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_325),
.B(n_326),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_288),
.B(n_263),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_327),
.Y(n_334)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_304),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_329),
.B(n_348),
.Y(n_354)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_331),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_314),
.A2(n_310),
.B1(n_257),
.B2(n_323),
.Y(n_332)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_332),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_311),
.C(n_319),
.Y(n_353)
);

OAI322xp33_ASAP7_75t_L g336 ( 
.A1(n_314),
.A2(n_320),
.A3(n_321),
.B1(n_282),
.B2(n_316),
.C1(n_318),
.C2(n_328),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_336),
.B(n_11),
.Y(n_360)
);

BUFx12_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_337),
.B(n_322),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_309),
.B(n_289),
.C(n_286),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_339),
.B(n_340),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_278),
.C(n_304),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_310),
.B(n_271),
.Y(n_341)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_341),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_327),
.A2(n_268),
.B1(n_305),
.B2(n_262),
.Y(n_343)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_343),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_311),
.B(n_282),
.Y(n_348)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_SL g375 ( 
.A(n_353),
.B(n_355),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_308),
.C(n_260),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_258),
.C(n_256),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_353),
.C(n_344),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_330),
.A2(n_302),
.B(n_128),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_357),
.B(n_334),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_348),
.B(n_11),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_359),
.B(n_329),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_364),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_335),
.A2(n_346),
.B1(n_340),
.B2(n_341),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_363),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_68),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_347),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_337),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_366),
.B(n_369),
.Y(n_387)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_368),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_349),
.A2(n_341),
.B1(n_334),
.B2(n_338),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_370),
.A2(n_376),
.B(n_377),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_350),
.A2(n_345),
.B1(n_337),
.B2(n_6),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_372),
.B(n_373),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_10),
.C(n_17),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_10),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_14),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_359),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_388),
.Y(n_393)
);

INVx13_ASAP7_75t_L g381 ( 
.A(n_374),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_381),
.B(n_383),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_375),
.A2(n_362),
.B(n_361),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_354),
.C(n_358),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_387),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_351),
.C(n_363),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_18),
.C(n_4),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_367),
.A2(n_8),
.B(n_16),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_384),
.B(n_371),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_391),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_385),
.A2(n_378),
.B1(n_366),
.B2(n_6),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_382),
.B(n_7),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_392),
.B(n_394),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_380),
.A2(n_7),
.B1(n_15),
.B2(n_16),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_395),
.Y(n_400)
);

A2O1A1O1Ixp25_ASAP7_75t_L g398 ( 
.A1(n_396),
.A2(n_388),
.B(n_381),
.C(n_379),
.D(n_18),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_398),
.B(n_5),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_389),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_393),
.Y(n_403)
);

A2O1A1Ixp33_ASAP7_75t_SL g402 ( 
.A1(n_393),
.A2(n_386),
.B(n_396),
.C(n_4),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_402),
.B(n_4),
.C(n_5),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_403),
.A2(n_405),
.B(n_406),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_404),
.B(n_402),
.C(n_397),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_5),
.Y(n_405)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_407),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_408),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_401),
.Y(n_411)
);


endmodule