module fake_netlist_6_309_n_198 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_198);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_198;

wire n_52;
wire n_91;
wire n_146;
wire n_46;
wire n_163;
wire n_119;
wire n_193;
wire n_147;
wire n_154;
wire n_191;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_131;
wire n_105;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_195;
wire n_189;
wire n_32;
wire n_85;
wire n_99;
wire n_130;
wire n_78;
wire n_84;
wire n_66;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_197;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_151;
wire n_110;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_108;
wire n_97;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_175;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_196;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_194;
wire n_171;
wire n_192;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_43),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2x1_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_1),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_36),
.B1(n_38),
.B2(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_51),
.B1(n_54),
.B2(n_7),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

AO22x2_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_81)
);

OAI221xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_2),
.B1(n_9),
.B2(n_31),
.C(n_13),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

AO22x2_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_9),
.B1(n_10),
.B2(n_18),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

OAI221xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.C(n_25),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_72),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_100),
.Y(n_105)
);

OAI31xp33_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_82),
.A3(n_92),
.B(n_58),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_79),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

O2A1O1Ixp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_57),
.B(n_87),
.C(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_104),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_104),
.Y(n_117)
);

AO21x2_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_92),
.B(n_82),
.Y(n_118)
);

AND2x4_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_94),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_98),
.B(n_101),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_64),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_107),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

AOI211xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_98),
.B(n_101),
.C(n_63),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_113),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

NAND4xp25_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_61),
.C(n_71),
.D(n_62),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_117),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_117),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_117),
.Y(n_141)
);

NAND2x1_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_115),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_90),
.Y(n_143)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_133),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_132),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_137),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_150),
.Y(n_156)
);

AND3x1_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_106),
.C(n_66),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_131),
.Y(n_158)
);

OAI31xp33_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_106),
.A3(n_97),
.B(n_70),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_81),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_57),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_75),
.C(n_70),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_57),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_67),
.Y(n_169)
);

NAND3x1_ASAP7_75t_SL g170 ( 
.A(n_159),
.B(n_81),
.C(n_97),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

OAI221xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_154),
.B1(n_160),
.B2(n_61),
.C(n_73),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_158),
.Y(n_176)
);

NAND3x1_ASAP7_75t_SL g177 ( 
.A(n_170),
.B(n_116),
.C(n_97),
.Y(n_177)
);

CKINVDCx6p67_ASAP7_75t_R g178 ( 
.A(n_166),
.Y(n_178)
);

AND2x4_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_142),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_168),
.B1(n_73),
.B2(n_169),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

AND2x4_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_73),
.Y(n_182)
);

NAND4xp75_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_111),
.C(n_105),
.D(n_97),
.Y(n_183)
);

NAND5xp2_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_75),
.C(n_19),
.D(n_118),
.E(n_65),
.Y(n_184)
);

OAI31xp33_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_75),
.A3(n_119),
.B(n_128),
.Y(n_185)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_178),
.B1(n_173),
.B2(n_172),
.Y(n_187)
);

AOI211xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_172),
.B(n_65),
.C(n_119),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_128),
.B1(n_119),
.B2(n_118),
.Y(n_190)
);

OAI322xp33_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_181),
.A3(n_185),
.B1(n_93),
.B2(n_94),
.C1(n_118),
.C2(n_110),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_114),
.B(n_185),
.C(n_189),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_114),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_114),
.B1(n_188),
.B2(n_187),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

NAND2x1p5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_114),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

AOI221xp5_ASAP7_75t_SL g198 ( 
.A1(n_195),
.A2(n_114),
.B1(n_191),
.B2(n_197),
.C(n_196),
.Y(n_198)
);


endmodule