module fake_netlist_6_3107_n_146 (n_16, n_1, n_34, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_0, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_146);

input n_16;
input n_1;
input n_34;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_0;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_146;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_138;
wire n_68;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_144;
wire n_127;
wire n_125;
wire n_77;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_75;
wire n_109;
wire n_122;
wire n_45;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_82;
wire n_38;
wire n_110;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

NOR2xp67_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_24),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

OA21x2_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_1),
.B(n_2),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_1),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_2),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_48),
.Y(n_77)
);

NAND2x1p5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_77),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_65),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_45),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_81),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_73),
.B(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_47),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_89),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_68),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

NAND2x1p5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_100),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_61),
.B1(n_82),
.B2(n_86),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

OAI21x1_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_97),
.B(n_103),
.Y(n_113)
);

OA21x2_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_99),
.B(n_96),
.Y(n_114)
);

AOI21x1_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_17),
.B(n_35),
.Y(n_115)
);

NAND2x1p5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_107),
.B(n_18),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_114),
.B(n_110),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_109),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_119),
.B1(n_115),
.B2(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_124),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_124),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_6),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_129),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);

AOI221x1_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_125),
.B1(n_132),
.B2(n_9),
.C(n_10),
.Y(n_137)
);

OAI211xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_7),
.B(n_12),
.C(n_13),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_21),
.Y(n_139)
);

NOR2x1_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_22),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_141),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_142),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_23),
.B1(n_25),
.B2(n_27),
.Y(n_144)
);

AOI22x1_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_145),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_146)
);


endmodule