module fake_jpeg_20707_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_0),
.B(n_1),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_52),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_29),
.B1(n_22),
.B2(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_29),
.B1(n_22),
.B2(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_29),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_30),
.B1(n_23),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_33),
.B1(n_40),
.B2(n_34),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_41),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_57),
.C(n_58),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_56),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_41),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_34),
.C(n_41),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_40),
.B1(n_32),
.B2(n_39),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_73),
.B1(n_64),
.B2(n_57),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_27),
.B1(n_26),
.B2(n_15),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_67),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_70),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_51),
.C(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_72),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_23),
.A3(n_26),
.B1(n_19),
.B2(n_20),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_39),
.B1(n_41),
.B2(n_21),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_0),
.B(n_1),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_74),
.B(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_24),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_2),
.Y(n_103)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_53),
.B1(n_47),
.B2(n_43),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_98),
.B1(n_99),
.B2(n_80),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_86),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_59),
.B1(n_66),
.B2(n_77),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g90 ( 
.A(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_96),
.Y(n_107)
);

AOI32xp33_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_54),
.A3(n_19),
.B1(n_20),
.B2(n_17),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_24),
.B1(n_21),
.B2(n_20),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_24),
.B1(n_21),
.B2(n_28),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_17),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_103),
.Y(n_119)
);

AOI22x1_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_74),
.B1(n_96),
.B2(n_93),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_113),
.B1(n_86),
.B2(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_108),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_57),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_118),
.B(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_28),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_83),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_71),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_125),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_79),
.B1(n_68),
.B2(n_67),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_28),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_122),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_2),
.B(n_3),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_4),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_124),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_88),
.B(n_14),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_88),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_119),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_143),
.B1(n_110),
.B2(n_106),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_137),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_100),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_139),
.B(n_133),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_91),
.B(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_119),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_98),
.B1(n_99),
.B2(n_91),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_121),
.Y(n_152)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_115),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_151),
.A2(n_159),
.B1(n_143),
.B2(n_129),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_141),
.B(n_133),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_120),
.C(n_112),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_135),
.C(n_138),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_104),
.B1(n_107),
.B2(n_106),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_139),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_130),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_97),
.Y(n_157)
);

NOR2xp67_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_145),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_144),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_104),
.B1(n_92),
.B2(n_97),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_160),
.B(n_159),
.Y(n_175)
);

OAI322xp33_ASAP7_75t_L g162 ( 
.A1(n_155),
.A2(n_126),
.A3(n_132),
.B1(n_141),
.B2(n_145),
.C1(n_135),
.C2(n_140),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_171),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_156),
.C(n_151),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_128),
.C(n_142),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_153),
.B(n_148),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_160),
.B1(n_158),
.B2(n_150),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_176),
.B1(n_172),
.B2(n_175),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_174),
.A2(n_171),
.B(n_169),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_163),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_168),
.A2(n_159),
.B1(n_147),
.B2(n_130),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_12),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_146),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_164),
.B(n_128),
.C(n_142),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_166),
.C(n_165),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_183),
.Y(n_188)
);

OAI31xp33_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_186),
.A3(n_6),
.B(n_7),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_184),
.B(n_185),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_180),
.A2(n_14),
.B(n_12),
.Y(n_186)
);

AOI31xp67_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_5),
.A3(n_6),
.B(n_7),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_176),
.B1(n_177),
.B2(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_192),
.B(n_7),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_189),
.A2(n_188),
.B(n_184),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_195),
.C(n_196),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_177),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_8),
.C(n_9),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_8),
.C(n_9),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_201),
.B(n_200),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_11),
.Y(n_203)
);


endmodule