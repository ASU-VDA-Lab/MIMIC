module fake_jpeg_12949_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_2),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_21),
.Y(n_31)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx5_ASAP7_75t_SL g30 ( 
.A(n_19),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_6),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_23),
.B(n_24),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_0),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_25),
.B(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_10),
.B(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_11),
.A2(n_13),
.B1(n_14),
.B2(n_12),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_10),
.B1(n_19),
.B2(n_24),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_25),
.B1(n_21),
.B2(n_16),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_31),
.Y(n_38)
);

AO22x1_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_34),
.B1(n_30),
.B2(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_36),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_37),
.C(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_39),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_30),
.B(n_37),
.Y(n_43)
);


endmodule