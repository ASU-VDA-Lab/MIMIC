module fake_jpeg_9241_n_180 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_20),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_34),
.B1(n_27),
.B2(n_22),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_36),
.A2(n_49),
.B1(n_44),
.B2(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_13),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_22),
.B1(n_25),
.B2(n_21),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_29),
.B(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_27),
.B1(n_18),
.B2(n_25),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_27),
.B1(n_21),
.B2(n_18),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_44),
.B1(n_41),
.B2(n_24),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_30),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_68),
.B1(n_44),
.B2(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_55),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_0),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_30),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_26),
.B1(n_13),
.B2(n_16),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_68),
.Y(n_78)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_42),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_29),
.C(n_28),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_50),
.B(n_1),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_2),
.B(n_3),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_84),
.B1(n_64),
.B2(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_30),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_50),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_89),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_31),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_0),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_1),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_54),
.B1(n_85),
.B2(n_87),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_103),
.B1(n_96),
.B2(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_100),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_53),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_104),
.B(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_105),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_65),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_78),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_59),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_108),
.B(n_90),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_113),
.C(n_119),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_116),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_79),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_70),
.C(n_76),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_74),
.B1(n_81),
.B2(n_71),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_104),
.B1(n_91),
.B2(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_108),
.B(n_101),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_82),
.C(n_86),
.Y(n_119)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_102),
.B1(n_101),
.B2(n_104),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_77),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_29),
.C(n_31),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_69),
.C(n_56),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_124),
.B(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_2),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_99),
.B(n_98),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_114),
.C(n_115),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_138),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_117),
.A2(n_19),
.B1(n_14),
.B2(n_24),
.Y(n_132)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_134),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_129),
.C(n_113),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_121),
.A2(n_14),
.B1(n_19),
.B2(n_23),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_23),
.B1(n_14),
.B2(n_19),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_137),
.B(n_23),
.Y(n_147)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_130),
.B(n_132),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_131),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_140),
.B(n_142),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_135),
.B(n_111),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_149),
.C(n_29),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_122),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_144),
.B(n_28),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_138),
.B1(n_134),
.B2(n_128),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_109),
.C(n_114),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_133),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_156),
.Y(n_165)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_155),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_141),
.B(n_126),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_145),
.B(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_38),
.B1(n_37),
.B2(n_28),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_38),
.B1(n_4),
.B2(n_5),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_3),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_3),
.C(n_4),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_162),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_161),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_4),
.C(n_5),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_151),
.B(n_154),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_168),
.C(n_6),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_153),
.B1(n_156),
.B2(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_5),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_6),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_173),
.Y(n_175)
);

AOI21x1_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_165),
.B(n_162),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_169),
.C(n_7),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_175),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_177),
.A2(n_6),
.B(n_8),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);


endmodule