module fake_jpeg_5052_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_22),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_56),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g103 ( 
.A(n_40),
.Y(n_103)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_46),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_43),
.B(n_47),
.Y(n_87)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_30),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_8),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_48),
.B(n_57),
.Y(n_94)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_59),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_15),
.B(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_34),
.B1(n_20),
.B2(n_21),
.Y(n_68)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_61),
.Y(n_88)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_62),
.A2(n_25),
.B1(n_11),
.B2(n_14),
.Y(n_109)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_71),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_20),
.B1(n_21),
.B2(n_34),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_65),
.A2(n_73),
.B(n_75),
.C(n_106),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_68),
.A2(n_78),
.B1(n_84),
.B2(n_100),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_18),
.B(n_23),
.C(n_24),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_69),
.B(n_102),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_21),
.B1(n_20),
.B2(n_30),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_82),
.B1(n_83),
.B2(n_91),
.Y(n_118)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_18),
.B1(n_23),
.B2(n_24),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_27),
.B(n_33),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_96),
.Y(n_115)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_79),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_30),
.B1(n_23),
.B2(n_24),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_86),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_31),
.B1(n_37),
.B2(n_36),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_15),
.B1(n_37),
.B2(n_36),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_31),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_16),
.Y(n_90)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_44),
.A2(n_16),
.B1(n_37),
.B2(n_17),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_95),
.Y(n_126)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_41),
.B(n_35),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_101),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_61),
.A2(n_16),
.B1(n_17),
.B2(n_25),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_41),
.Y(n_102)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_35),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_109),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_56),
.A2(n_27),
.B(n_33),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_62),
.A2(n_25),
.B1(n_17),
.B2(n_35),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_110),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_58),
.A2(n_32),
.B1(n_28),
.B2(n_38),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_62),
.A2(n_32),
.B1(n_28),
.B2(n_38),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_33),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_33),
.C(n_32),
.Y(n_129)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_116),
.Y(n_145)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_1),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_67),
.B(n_2),
.Y(n_124)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_128),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_81),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_103),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_33),
.B(n_32),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_28),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_81),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_132),
.Y(n_160)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_138),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_67),
.B(n_3),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_79),
.Y(n_148)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_81),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_139),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_98),
.Y(n_178)
);

NAND2x1p5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_67),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_144),
.A2(n_164),
.B(n_169),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_140),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_151),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_148),
.B(n_177),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_110),
.B1(n_109),
.B2(n_107),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_152),
.B1(n_159),
.B2(n_161),
.Y(n_180)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_69),
.B1(n_70),
.B2(n_111),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_157),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_119),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_158),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_102),
.C(n_74),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_114),
.C(n_125),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_94),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_65),
.B1(n_77),
.B2(n_86),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_108),
.B1(n_85),
.B2(n_93),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_126),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_173),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_170),
.C(n_174),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_134),
.B(n_123),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_97),
.B1(n_87),
.B2(n_99),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_132),
.B1(n_116),
.B2(n_112),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_87),
.A3(n_63),
.B1(n_95),
.B2(n_71),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_168),
.Y(n_204)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_115),
.B(n_88),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_101),
.B(n_33),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_120),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_118),
.A2(n_80),
.B1(n_99),
.B2(n_104),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_171),
.A2(n_117),
.B1(n_139),
.B2(n_10),
.Y(n_202)
);

XOR2x2_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_28),
.Y(n_172)
);

XOR2x2_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_118),
.Y(n_190)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

AND2x6_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_92),
.Y(n_174)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_3),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_3),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_121),
.B(n_114),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_181),
.A2(n_214),
.B(n_182),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_183),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_184),
.B(n_198),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g188 ( 
.A(n_146),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_194),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_191),
.C(n_192),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_146),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_92),
.C(n_64),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_170),
.C(n_168),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_193),
.A2(n_202),
.B1(n_151),
.B2(n_117),
.Y(n_235)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_98),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_145),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_200),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_10),
.Y(n_205)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_207),
.Y(n_233)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_152),
.A2(n_117),
.B1(n_5),
.B2(n_6),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_12),
.B1(n_14),
.B2(n_8),
.Y(n_237)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_210),
.B(n_211),
.Y(n_223)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_166),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_172),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_218),
.C(n_182),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_172),
.B(n_177),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_217),
.A2(n_224),
.B(n_230),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_155),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_222),
.Y(n_242)
);

A2O1A1O1Ixp25_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_177),
.B(n_149),
.C(n_164),
.D(n_159),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_220),
.A2(n_231),
.B(n_238),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_163),
.B(n_158),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_229),
.B(n_184),
.Y(n_259)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_193),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_203),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_207),
.A2(n_148),
.B(n_157),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_187),
.A2(n_162),
.B(n_153),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_237),
.B1(n_186),
.B2(n_183),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_187),
.A2(n_154),
.B(n_176),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_201),
.B1(n_214),
.B2(n_210),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_241),
.A2(n_257),
.B1(n_240),
.B2(n_229),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_245),
.C(n_251),
.Y(n_264)
);

OAI32xp33_ASAP7_75t_L g244 ( 
.A1(n_225),
.A2(n_180),
.A3(n_208),
.B1(n_206),
.B2(n_192),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_253),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_191),
.C(n_180),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_194),
.Y(n_246)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_221),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_249),
.A2(n_250),
.B(n_255),
.Y(n_265)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_189),
.C(n_181),
.Y(n_251)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_209),
.C(n_200),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_211),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_232),
.Y(n_256)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_232),
.A2(n_199),
.B1(n_186),
.B2(n_196),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_258),
.A2(n_222),
.B1(n_219),
.B2(n_231),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_260),
.B(n_217),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_173),
.C(n_154),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_262),
.A2(n_248),
.B(n_246),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_223),
.B1(n_224),
.B2(n_230),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_268),
.B1(n_271),
.B2(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_269),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_223),
.B1(n_237),
.B2(n_220),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_216),
.B1(n_218),
.B2(n_234),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_249),
.A2(n_236),
.B1(n_215),
.B2(n_212),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_215),
.B1(n_212),
.B2(n_226),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_273),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_282),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_245),
.B1(n_240),
.B2(n_251),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_281),
.B1(n_261),
.B2(n_270),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_241),
.B1(n_257),
.B2(n_248),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_275),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_244),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_268),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_243),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_286),
.C(n_287),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_260),
.C(n_242),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_262),
.C(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_247),
.C(n_213),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_5),
.C(n_7),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_294),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_272),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_5),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_286),
.Y(n_304)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_289),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_299),
.Y(n_305)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_8),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_284),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_11),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_292),
.A2(n_279),
.B1(n_276),
.B2(n_281),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_304),
.B1(n_5),
.B2(n_7),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_297),
.B(n_287),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_307),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_9),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_293),
.C(n_291),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_301),
.A2(n_300),
.B1(n_293),
.B2(n_10),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_311),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_312),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_313),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_305),
.Y(n_319)
);


endmodule