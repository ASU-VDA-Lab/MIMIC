module real_aes_9137_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_725;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g467 ( .A1(n_0), .A2(n_145), .B(n_468), .C(n_471), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_1), .B(n_462), .Y(n_473) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g183 ( .A(n_3), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_4), .B(n_146), .Y(n_545) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_5), .A2(n_124), .B1(n_125), .B2(n_431), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_5), .Y(n_431) );
OAI22xp5_ASAP7_75t_SL g738 ( .A1(n_5), .A2(n_95), .B1(n_431), .B2(n_739), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_6), .A2(n_447), .B(n_494), .Y(n_493) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_7), .A2(n_152), .B(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_8), .A2(n_36), .B1(n_149), .B2(n_201), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_9), .B(n_152), .Y(n_169) );
AND2x6_ASAP7_75t_L g154 ( .A(n_10), .B(n_155), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_11), .A2(n_154), .B(n_450), .C(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_12), .B(n_38), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_12), .B(n_38), .Y(n_436) );
INVx1_ASAP7_75t_L g136 ( .A(n_13), .Y(n_136) );
INVx1_ASAP7_75t_L g175 ( .A(n_14), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_15), .B(n_142), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_16), .B(n_146), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_17), .B(n_132), .Y(n_131) );
AO32x2_ASAP7_75t_L g212 ( .A1(n_18), .A2(n_152), .A3(n_153), .B1(n_172), .B2(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_19), .B(n_149), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_20), .B(n_132), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_21), .A2(n_54), .B1(n_149), .B2(n_201), .Y(n_215) );
AOI22xp33_ASAP7_75t_SL g209 ( .A1(n_22), .A2(n_80), .B1(n_142), .B2(n_149), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_23), .B(n_149), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_24), .A2(n_153), .B(n_450), .C(n_452), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_25), .A2(n_153), .B(n_450), .C(n_528), .Y(n_527) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_26), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_27), .A2(n_96), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_27), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_28), .B(n_191), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_29), .A2(n_447), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_30), .B(n_191), .Y(n_228) );
INVx2_ASAP7_75t_L g144 ( .A(n_31), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_32), .A2(n_482), .B(n_483), .C(n_487), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_33), .B(n_149), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_34), .B(n_191), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_35), .B(n_197), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_37), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_39), .B(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_40), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_41), .B(n_146), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_42), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_43), .B(n_447), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_44), .A2(n_482), .B(n_487), .C(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_45), .B(n_149), .Y(n_162) );
INVx1_ASAP7_75t_L g469 ( .A(n_46), .Y(n_469) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_47), .A2(n_737), .B1(n_740), .B2(n_741), .Y(n_736) );
INVx1_ASAP7_75t_L g741 ( .A(n_47), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_48), .A2(n_89), .B1(n_201), .B2(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g508 ( .A(n_49), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_50), .B(n_149), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_51), .B(n_149), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_52), .B(n_447), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_53), .B(n_167), .Y(n_166) );
AOI22xp33_ASAP7_75t_SL g148 ( .A1(n_55), .A2(n_59), .B1(n_142), .B2(n_149), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_56), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_57), .B(n_149), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_58), .B(n_149), .Y(n_248) );
INVx1_ASAP7_75t_L g155 ( .A(n_60), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_61), .B(n_447), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_62), .B(n_462), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_63), .A2(n_167), .B(n_178), .C(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_64), .B(n_149), .Y(n_184) );
INVx1_ASAP7_75t_L g135 ( .A(n_65), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_66), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_67), .B(n_146), .Y(n_485) );
AO32x2_ASAP7_75t_L g205 ( .A1(n_68), .A2(n_152), .A3(n_153), .B1(n_206), .B2(n_210), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_69), .B(n_147), .Y(n_519) );
INVx1_ASAP7_75t_L g247 ( .A(n_70), .Y(n_247) );
INVx1_ASAP7_75t_L g223 ( .A(n_71), .Y(n_223) );
CKINVDCx16_ASAP7_75t_R g465 ( .A(n_72), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_73), .B(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_74), .A2(n_103), .B1(n_116), .B2(n_748), .Y(n_102) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_75), .A2(n_450), .B(n_487), .C(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_76), .B(n_142), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_77), .Y(n_495) );
INVx1_ASAP7_75t_L g115 ( .A(n_78), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_79), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_81), .B(n_201), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_82), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_83), .B(n_142), .Y(n_227) );
INVx2_ASAP7_75t_L g133 ( .A(n_84), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_85), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_86), .B(n_139), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_87), .B(n_142), .Y(n_163) );
INVx2_ASAP7_75t_L g112 ( .A(n_88), .Y(n_112) );
OR2x2_ASAP7_75t_L g434 ( .A(n_88), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g735 ( .A(n_88), .B(n_729), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_90), .A2(n_101), .B1(n_142), .B2(n_143), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_91), .B(n_447), .Y(n_480) );
INVx1_ASAP7_75t_L g484 ( .A(n_92), .Y(n_484) );
INVxp67_ASAP7_75t_L g498 ( .A(n_93), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_94), .B(n_142), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_95), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_96), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_97), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g515 ( .A(n_98), .Y(n_515) );
INVx1_ASAP7_75t_L g544 ( .A(n_99), .Y(n_544) );
AND2x2_ASAP7_75t_L g510 ( .A(n_100), .B(n_191), .Y(n_510) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx9p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g749 ( .A(n_106), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_112), .C(n_113), .Y(n_110) );
AND2x2_ASAP7_75t_L g435 ( .A(n_111), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g721 ( .A(n_112), .B(n_435), .Y(n_721) );
NOR2x2_ASAP7_75t_L g728 ( .A(n_112), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AO221x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_730), .B1(n_733), .B2(n_742), .C(n_744), .Y(n_116) );
OAI222xp33_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_121), .B1(n_722), .B2(n_723), .C1(n_726), .C2(n_727), .Y(n_117) );
INVx1_ASAP7_75t_L g722 ( .A(n_118), .Y(n_722) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_432), .B1(n_437), .B2(n_719), .Y(n_122) );
INVx1_ASAP7_75t_L g725 ( .A(n_123), .Y(n_725) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
XNOR2xp5_ASAP7_75t_L g737 ( .A(n_125), .B(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_SL g125 ( .A(n_126), .B(n_365), .Y(n_125) );
NOR5xp2_ASAP7_75t_L g126 ( .A(n_127), .B(n_278), .C(n_324), .D(n_337), .E(n_349), .Y(n_126) );
OAI211xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_186), .B(n_232), .C(n_259), .Y(n_127) );
INVx1_ASAP7_75t_SL g360 ( .A(n_128), .Y(n_360) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_156), .Y(n_128) );
AND2x2_ASAP7_75t_L g284 ( .A(n_129), .B(n_157), .Y(n_284) );
AND2x2_ASAP7_75t_L g312 ( .A(n_129), .B(n_258), .Y(n_312) );
AND2x2_ASAP7_75t_L g320 ( .A(n_129), .B(n_263), .Y(n_320) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g250 ( .A(n_130), .B(n_158), .Y(n_250) );
INVx2_ASAP7_75t_L g262 ( .A(n_130), .Y(n_262) );
AND2x2_ASAP7_75t_L g387 ( .A(n_130), .B(n_329), .Y(n_387) );
OR2x2_ASAP7_75t_L g389 ( .A(n_130), .B(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_137), .Y(n_130) );
INVx1_ASAP7_75t_L g256 ( .A(n_131), .Y(n_256) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_132), .Y(n_152) );
INVx1_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g191 ( .A(n_133), .B(n_134), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
NAND3xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_151), .C(n_153), .Y(n_137) );
AO21x1_ASAP7_75t_L g255 ( .A1(n_138), .A2(n_151), .B(n_256), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_141), .B1(n_145), .B2(n_148), .Y(n_138) );
INVx2_ASAP7_75t_L g202 ( .A(n_139), .Y(n_202) );
OAI22xp5_ASAP7_75t_SL g206 ( .A1(n_139), .A2(n_147), .B1(n_207), .B2(n_209), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_139), .A2(n_145), .B1(n_214), .B2(n_215), .Y(n_213) );
INVx4_ASAP7_75t_L g470 ( .A(n_139), .Y(n_470) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g147 ( .A(n_140), .Y(n_147) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_140), .Y(n_180) );
INVx1_ASAP7_75t_L g197 ( .A(n_140), .Y(n_197) );
AND2x2_ASAP7_75t_L g448 ( .A(n_140), .B(n_168), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_140), .Y(n_451) );
INVx2_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g150 ( .A(n_144), .Y(n_150) );
INVx1_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_145), .A2(n_165), .B(n_166), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_145), .A2(n_182), .B(n_183), .C(n_184), .Y(n_181) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_146), .A2(n_162), .B(n_163), .Y(n_161) );
O2A1O1Ixp5_ASAP7_75t_SL g221 ( .A1(n_146), .A2(n_222), .B(n_223), .C(n_224), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_146), .A2(n_244), .B(n_245), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_146), .B(n_498), .Y(n_497) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g222 ( .A(n_149), .Y(n_222) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_149), .Y(n_546) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g201 ( .A(n_150), .Y(n_201) );
BUFx3_ASAP7_75t_L g208 ( .A(n_150), .Y(n_208) );
AND2x6_ASAP7_75t_L g450 ( .A(n_150), .B(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g462 ( .A(n_151), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_151), .B(n_489), .Y(n_488) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_151), .A2(n_514), .B(n_521), .Y(n_513) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_151), .A2(n_541), .B(n_548), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_151), .B(n_549), .Y(n_548) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_152), .A2(n_160), .B(n_169), .Y(n_159) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_152), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_152), .A2(n_526), .B(n_527), .Y(n_525) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_153), .A2(n_243), .B(n_246), .Y(n_242) );
BUFx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OAI21xp5_ASAP7_75t_L g160 ( .A1(n_154), .A2(n_161), .B(n_164), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g173 ( .A1(n_154), .A2(n_174), .B(n_181), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_154), .A2(n_193), .B(n_198), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_154), .A2(n_221), .B(n_225), .Y(n_220) );
AND2x4_ASAP7_75t_L g447 ( .A(n_154), .B(n_448), .Y(n_447) );
INVx4_ASAP7_75t_SL g472 ( .A(n_154), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g516 ( .A(n_154), .B(n_448), .Y(n_516) );
INVx2_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g300 ( .A(n_157), .B(n_272), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_157), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g414 ( .A(n_157), .B(n_254), .Y(n_414) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_170), .Y(n_157) );
AND2x2_ASAP7_75t_L g257 ( .A(n_158), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g304 ( .A(n_158), .Y(n_304) );
AND2x2_ASAP7_75t_L g329 ( .A(n_158), .B(n_241), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_158), .B(n_362), .Y(n_399) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g263 ( .A(n_159), .B(n_241), .Y(n_263) );
AND2x2_ASAP7_75t_L g277 ( .A(n_159), .B(n_240), .Y(n_277) );
AND2x2_ASAP7_75t_L g294 ( .A(n_159), .B(n_170), .Y(n_294) );
AND2x2_ASAP7_75t_L g351 ( .A(n_159), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_159), .B(n_258), .Y(n_364) );
AND2x2_ASAP7_75t_L g416 ( .A(n_159), .B(n_341), .Y(n_416) );
INVx2_ASAP7_75t_L g182 ( .A(n_167), .Y(n_182) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g239 ( .A(n_170), .B(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g258 ( .A(n_170), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_170), .B(n_241), .Y(n_335) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_173), .B(n_185), .Y(n_170) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_171), .A2(n_242), .B(n_249), .Y(n_241) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_172), .B(n_522), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_178), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_176), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_176), .A2(n_529), .B(n_530), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_178), .A2(n_544), .B(n_545), .C(n_546), .Y(n_543) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_179), .A2(n_226), .B(n_227), .Y(n_225) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g454 ( .A(n_180), .Y(n_454) );
O2A1O1Ixp5_ASAP7_75t_L g246 ( .A1(n_182), .A2(n_202), .B(n_247), .C(n_248), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_182), .A2(n_453), .B(n_455), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_216), .B(n_229), .Y(n_186) );
INVx1_ASAP7_75t_SL g348 ( .A(n_187), .Y(n_348) );
AND2x4_ASAP7_75t_L g187 ( .A(n_188), .B(n_204), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_SL g236 ( .A(n_189), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g231 ( .A(n_190), .Y(n_231) );
INVx1_ASAP7_75t_L g268 ( .A(n_190), .Y(n_268) );
AND2x2_ASAP7_75t_L g289 ( .A(n_190), .B(n_211), .Y(n_289) );
AND2x2_ASAP7_75t_L g323 ( .A(n_190), .B(n_212), .Y(n_323) );
OR2x2_ASAP7_75t_L g342 ( .A(n_190), .B(n_218), .Y(n_342) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_190), .Y(n_356) );
AND2x2_ASAP7_75t_L g369 ( .A(n_190), .B(n_370), .Y(n_369) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_203), .Y(n_190) );
INVx2_ASAP7_75t_L g210 ( .A(n_191), .Y(n_210) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_191), .A2(n_220), .B(n_228), .Y(n_219) );
INVx1_ASAP7_75t_L g460 ( .A(n_191), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_191), .A2(n_480), .B(n_481), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_191), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_196), .Y(n_193) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_202), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_204), .A2(n_291), .B1(n_292), .B2(n_301), .Y(n_290) );
AND2x2_ASAP7_75t_L g374 ( .A(n_204), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_211), .Y(n_204) );
INVx1_ASAP7_75t_L g235 ( .A(n_205), .Y(n_235) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_205), .Y(n_272) );
INVx1_ASAP7_75t_L g283 ( .A(n_205), .Y(n_283) );
AND2x2_ASAP7_75t_L g298 ( .A(n_205), .B(n_212), .Y(n_298) );
INVx2_ASAP7_75t_L g471 ( .A(n_208), .Y(n_471) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_208), .Y(n_486) );
INVx1_ASAP7_75t_L g457 ( .A(n_210), .Y(n_457) );
OR2x2_ASAP7_75t_L g252 ( .A(n_211), .B(n_237), .Y(n_252) );
AND2x2_ASAP7_75t_L g282 ( .A(n_211), .B(n_283), .Y(n_282) );
NOR2xp67_ASAP7_75t_L g370 ( .A(n_211), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g230 ( .A(n_212), .B(n_231), .Y(n_230) );
BUFx2_ASAP7_75t_L g339 ( .A(n_212), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_216), .B(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g317 ( .A(n_217), .B(n_283), .Y(n_317) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g229 ( .A(n_218), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g288 ( .A(n_218), .Y(n_288) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g237 ( .A(n_219), .Y(n_237) );
OR2x2_ASAP7_75t_L g267 ( .A(n_219), .B(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_219), .Y(n_322) );
AOI32xp33_ASAP7_75t_L g359 ( .A1(n_229), .A2(n_289), .A3(n_360), .B1(n_361), .B2(n_363), .Y(n_359) );
AND2x2_ASAP7_75t_L g285 ( .A(n_230), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_230), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_230), .B(n_317), .Y(n_403) );
INVx1_ASAP7_75t_L g408 ( .A(n_230), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_238), .B1(n_251), .B2(n_253), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_236), .Y(n_233) );
AND2x2_ASAP7_75t_L g338 ( .A(n_234), .B(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_235), .B(n_237), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_236), .A2(n_260), .B1(n_264), .B2(n_274), .Y(n_259) );
AND2x2_ASAP7_75t_L g281 ( .A(n_236), .B(n_282), .Y(n_281) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_236), .A2(n_250), .B(n_298), .C(n_333), .Y(n_332) );
OAI332xp33_ASAP7_75t_L g337 ( .A1(n_236), .A2(n_338), .A3(n_340), .B1(n_342), .B2(n_343), .B3(n_345), .C1(n_346), .C2(n_348), .Y(n_337) );
INVx2_ASAP7_75t_L g378 ( .A(n_236), .Y(n_378) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_237), .Y(n_296) );
INVx1_ASAP7_75t_L g371 ( .A(n_237), .Y(n_371) );
AND2x2_ASAP7_75t_L g425 ( .A(n_237), .B(n_289), .Y(n_425) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_250), .Y(n_238) );
AND2x2_ASAP7_75t_L g305 ( .A(n_240), .B(n_255), .Y(n_305) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g254 ( .A(n_241), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g353 ( .A(n_241), .B(n_255), .Y(n_353) );
INVx1_ASAP7_75t_L g362 ( .A(n_241), .Y(n_362) );
INVx1_ASAP7_75t_L g336 ( .A(n_250), .Y(n_336) );
INVxp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g420 ( .A(n_252), .B(n_272), .Y(n_420) );
INVx1_ASAP7_75t_SL g331 ( .A(n_253), .Y(n_331) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_257), .Y(n_253) );
AND2x2_ASAP7_75t_L g358 ( .A(n_254), .B(n_316), .Y(n_358) );
INVx1_ASAP7_75t_L g377 ( .A(n_254), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_254), .B(n_344), .Y(n_379) );
INVx1_ASAP7_75t_L g276 ( .A(n_255), .Y(n_276) );
AND2x2_ASAP7_75t_L g280 ( .A(n_257), .B(n_261), .Y(n_280) );
AND2x2_ASAP7_75t_L g347 ( .A(n_257), .B(n_305), .Y(n_347) );
INVx2_ASAP7_75t_L g390 ( .A(n_257), .Y(n_390) );
INVx2_ASAP7_75t_L g273 ( .A(n_258), .Y(n_273) );
AND2x2_ASAP7_75t_L g275 ( .A(n_258), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
INVx1_ASAP7_75t_L g291 ( .A(n_261), .Y(n_291) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_262), .B(n_335), .Y(n_341) );
OR2x2_ASAP7_75t_L g405 ( .A(n_262), .B(n_364), .Y(n_405) );
INVx1_ASAP7_75t_L g429 ( .A(n_262), .Y(n_429) );
INVx1_ASAP7_75t_L g385 ( .A(n_263), .Y(n_385) );
AND2x2_ASAP7_75t_L g430 ( .A(n_263), .B(n_273), .Y(n_430) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_269), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_267), .A2(n_293), .B1(n_295), .B2(n_299), .Y(n_292) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OAI322xp33_ASAP7_75t_SL g376 ( .A1(n_270), .A2(n_377), .A3(n_378), .B1(n_379), .B2(n_380), .C1(n_383), .C2(n_385), .Y(n_376) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
AND2x2_ASAP7_75t_L g373 ( .A(n_271), .B(n_289), .Y(n_373) );
OR2x2_ASAP7_75t_L g407 ( .A(n_271), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g410 ( .A(n_271), .B(n_342), .Y(n_410) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g355 ( .A(n_272), .B(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g411 ( .A(n_272), .B(n_342), .Y(n_411) );
INVx3_ASAP7_75t_L g344 ( .A(n_273), .Y(n_344) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g400 ( .A(n_275), .Y(n_400) );
AOI222xp33_ASAP7_75t_L g279 ( .A1(n_277), .A2(n_280), .B1(n_281), .B2(n_284), .C1(n_285), .C2(n_287), .Y(n_279) );
INVx1_ASAP7_75t_L g310 ( .A(n_277), .Y(n_310) );
NAND3xp33_ASAP7_75t_SL g278 ( .A(n_279), .B(n_290), .C(n_307), .Y(n_278) );
AND2x2_ASAP7_75t_L g395 ( .A(n_282), .B(n_296), .Y(n_395) );
BUFx2_ASAP7_75t_L g286 ( .A(n_283), .Y(n_286) );
INVx1_ASAP7_75t_L g327 ( .A(n_283), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_284), .A2(n_320), .B1(n_373), .B2(n_374), .C(n_376), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_286), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_289), .Y(n_313) );
AND2x2_ASAP7_75t_L g326 ( .A(n_289), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_294), .B(n_305), .Y(n_306) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
OAI21xp33_ASAP7_75t_L g301 ( .A1(n_296), .A2(n_302), .B(n_306), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_296), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g393 ( .A(n_298), .B(n_375), .Y(n_393) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g316 ( .A(n_304), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_305), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g422 ( .A(n_305), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_313), .B1(n_314), .B2(n_317), .C(n_318), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_309), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g418 ( .A(n_317), .B(n_323), .Y(n_418) );
INVxp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
OAI31xp33_ASAP7_75t_SL g386 ( .A1(n_321), .A2(n_360), .A3(n_387), .B(n_388), .Y(n_386) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g375 ( .A(n_322), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_323), .B(n_327), .Y(n_426) );
OAI221xp5_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_328), .B1(n_330), .B2(n_331), .C(n_332), .Y(n_324) );
INVx1_ASAP7_75t_L g330 ( .A(n_326), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_329), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g345 ( .A(n_338), .Y(n_345) );
INVx2_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g367 ( .A(n_344), .B(n_353), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g417 ( .A1(n_344), .A2(n_361), .B(n_418), .C(n_419), .Y(n_417) );
OAI221xp5_ASAP7_75t_SL g349 ( .A1(n_345), .A2(n_350), .B1(n_354), .B2(n_357), .C(n_359), .Y(n_349) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_L g412 ( .A1(n_348), .A2(n_413), .B(n_415), .C(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_351), .A2(n_402), .B1(n_404), .B2(n_406), .C(n_409), .Y(n_401) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
NOR4xp25_ASAP7_75t_L g365 ( .A(n_366), .B(n_391), .C(n_412), .D(n_423), .Y(n_365) );
OAI211xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_368), .B(n_372), .C(n_386), .Y(n_366) );
INVx1_ASAP7_75t_SL g421 ( .A(n_373), .Y(n_421) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_SL g384 ( .A(n_382), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_389), .A2(n_398), .B1(n_410), .B2(n_411), .Y(n_409) );
A2O1A1Ixp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_396), .C(n_401), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI31xp33_ASAP7_75t_L g423 ( .A1(n_394), .A2(n_424), .A3(n_426), .B(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B(n_422), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_434), .A2(n_438), .B1(n_721), .B2(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g729 ( .A(n_435), .Y(n_729) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_SL g438 ( .A(n_439), .B(n_655), .Y(n_438) );
NOR5xp2_ASAP7_75t_L g439 ( .A(n_440), .B(n_586), .C(n_615), .D(n_635), .E(n_642), .Y(n_439) );
OAI211xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_474), .B(n_531), .C(n_573), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_442), .A2(n_658), .B1(n_660), .B2(n_661), .Y(n_657) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_461), .Y(n_442) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_443), .Y(n_534) );
AND2x4_ASAP7_75t_L g566 ( .A(n_443), .B(n_567), .Y(n_566) );
INVx5_ASAP7_75t_L g584 ( .A(n_443), .Y(n_584) );
AND2x2_ASAP7_75t_L g593 ( .A(n_443), .B(n_585), .Y(n_593) );
AND2x2_ASAP7_75t_L g605 ( .A(n_443), .B(n_478), .Y(n_605) );
AND2x2_ASAP7_75t_L g701 ( .A(n_443), .B(n_569), .Y(n_701) );
OR2x6_ASAP7_75t_L g443 ( .A(n_444), .B(n_458), .Y(n_443) );
AOI21xp5_ASAP7_75t_SL g444 ( .A1(n_445), .A2(n_449), .B(n_457), .Y(n_444) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx5_ASAP7_75t_L g466 ( .A(n_450), .Y(n_466) );
INVx2_ASAP7_75t_L g456 ( .A(n_454), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_456), .A2(n_484), .B(n_485), .C(n_486), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_456), .A2(n_486), .B(n_508), .C(n_509), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVx2_ASAP7_75t_L g567 ( .A(n_461), .Y(n_567) );
AND2x2_ASAP7_75t_L g585 ( .A(n_461), .B(n_540), .Y(n_585) );
AND2x2_ASAP7_75t_L g604 ( .A(n_461), .B(n_539), .Y(n_604) );
AND2x2_ASAP7_75t_L g644 ( .A(n_461), .B(n_584), .Y(n_644) );
OA21x2_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B(n_473), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_466), .B(n_467), .C(n_472), .Y(n_464) );
INVx2_ASAP7_75t_L g482 ( .A(n_466), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_466), .A2(n_472), .B(n_495), .C(n_496), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g487 ( .A(n_472), .Y(n_487) );
INVxp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_500), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AOI322xp5_ASAP7_75t_L g703 ( .A1(n_477), .A2(n_511), .A3(n_558), .B1(n_566), .B2(n_620), .C1(n_704), .C2(n_707), .Y(n_703) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_490), .Y(n_477) );
INVx5_ASAP7_75t_L g536 ( .A(n_478), .Y(n_536) );
AND2x2_ASAP7_75t_L g552 ( .A(n_478), .B(n_538), .Y(n_552) );
BUFx2_ASAP7_75t_L g630 ( .A(n_478), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_478), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g707 ( .A(n_478), .B(n_614), .Y(n_707) );
OR2x6_ASAP7_75t_L g478 ( .A(n_479), .B(n_488), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_490), .B(n_502), .Y(n_561) );
INVx1_ASAP7_75t_L g588 ( .A(n_490), .Y(n_588) );
AND2x2_ASAP7_75t_L g601 ( .A(n_490), .B(n_523), .Y(n_601) );
AND2x2_ASAP7_75t_L g702 ( .A(n_490), .B(n_620), .Y(n_702) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g556 ( .A(n_491), .B(n_502), .Y(n_556) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_491), .Y(n_564) );
OR2x2_ASAP7_75t_L g571 ( .A(n_491), .B(n_523), .Y(n_571) );
AND2x2_ASAP7_75t_L g581 ( .A(n_491), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_491), .B(n_513), .Y(n_610) );
INVxp67_ASAP7_75t_L g634 ( .A(n_491), .Y(n_634) );
AND2x2_ASAP7_75t_L g641 ( .A(n_491), .B(n_511), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_491), .B(n_523), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_491), .B(n_512), .Y(n_667) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B(n_499), .Y(n_491) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_511), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_502), .B(n_524), .Y(n_611) );
OR2x2_ASAP7_75t_L g633 ( .A(n_502), .B(n_512), .Y(n_633) );
AND2x2_ASAP7_75t_L g646 ( .A(n_502), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_502), .B(n_601), .Y(n_652) );
OAI211xp5_ASAP7_75t_SL g656 ( .A1(n_502), .A2(n_657), .B(n_662), .C(n_671), .Y(n_656) );
AND2x2_ASAP7_75t_L g717 ( .A(n_502), .B(n_523), .Y(n_717) );
INVx5_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g570 ( .A(n_503), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_503), .B(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_503), .B(n_565), .Y(n_577) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_503), .Y(n_579) );
OR2x2_ASAP7_75t_L g590 ( .A(n_503), .B(n_512), .Y(n_590) );
AND2x2_ASAP7_75t_SL g595 ( .A(n_503), .B(n_581), .Y(n_595) );
AND2x2_ASAP7_75t_L g620 ( .A(n_503), .B(n_512), .Y(n_620) );
AND2x2_ASAP7_75t_L g640 ( .A(n_503), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g678 ( .A(n_503), .B(n_511), .Y(n_678) );
OR2x2_ASAP7_75t_L g681 ( .A(n_503), .B(n_667), .Y(n_681) );
OR2x6_ASAP7_75t_L g503 ( .A(n_504), .B(n_510), .Y(n_503) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_523), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g624 ( .A1(n_512), .A2(n_625), .B(n_628), .C(n_634), .Y(n_624) );
INVx5_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_513), .B(n_523), .Y(n_555) );
AND2x2_ASAP7_75t_L g559 ( .A(n_513), .B(n_524), .Y(n_559) );
OR2x2_ASAP7_75t_L g565 ( .A(n_513), .B(n_523), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
INVx1_ASAP7_75t_SL g582 ( .A(n_523), .Y(n_582) );
OR2x2_ASAP7_75t_L g710 ( .A(n_523), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_550), .B(n_553), .C(n_562), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AOI31xp33_ASAP7_75t_L g635 ( .A1(n_533), .A2(n_636), .A3(n_638), .B(n_639), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_534), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_535), .B(n_566), .Y(n_572) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_536), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g592 ( .A(n_536), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g597 ( .A(n_536), .B(n_567), .Y(n_597) );
AND2x2_ASAP7_75t_L g607 ( .A(n_536), .B(n_566), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_536), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g627 ( .A(n_536), .B(n_584), .Y(n_627) );
AND2x2_ASAP7_75t_L g632 ( .A(n_536), .B(n_604), .Y(n_632) );
OR2x2_ASAP7_75t_L g651 ( .A(n_536), .B(n_538), .Y(n_651) );
OR2x2_ASAP7_75t_L g653 ( .A(n_536), .B(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_536), .Y(n_700) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g600 ( .A(n_538), .B(n_567), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_538), .B(n_584), .Y(n_623) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g569 ( .A(n_540), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_547), .Y(n_541) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g660 ( .A(n_552), .B(n_584), .Y(n_660) );
AOI322xp5_ASAP7_75t_L g662 ( .A1(n_552), .A2(n_566), .A3(n_604), .B1(n_663), .B2(n_664), .C1(n_665), .C2(n_668), .Y(n_662) );
INVx1_ASAP7_75t_L g670 ( .A(n_552), .Y(n_670) );
NAND2xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
INVx1_ASAP7_75t_SL g664 ( .A(n_554), .Y(n_664) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
OR2x2_ASAP7_75t_L g616 ( .A(n_555), .B(n_561), .Y(n_616) );
INVx1_ASAP7_75t_L g647 ( .A(n_555), .Y(n_647) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OAI32xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_566), .A3(n_568), .B1(n_570), .B2(n_572), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AOI21xp33_ASAP7_75t_SL g602 ( .A1(n_565), .A2(n_580), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_SL g617 ( .A(n_566), .Y(n_617) );
AND2x4_ASAP7_75t_L g614 ( .A(n_567), .B(n_584), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_567), .B(n_650), .Y(n_649) );
AOI322xp5_ASAP7_75t_L g679 ( .A1(n_568), .A2(n_595), .A3(n_614), .B1(n_647), .B2(n_680), .C1(n_682), .C2(n_683), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_568), .A2(n_645), .B1(n_709), .B2(n_710), .C(n_712), .Y(n_708) );
AND2x2_ASAP7_75t_L g596 ( .A(n_569), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_SL g576 ( .A(n_571), .Y(n_576) );
OR2x2_ASAP7_75t_L g648 ( .A(n_571), .B(n_633), .Y(n_648) );
OAI31xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_577), .A3(n_578), .B(n_583), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_574), .A2(n_607), .B1(n_608), .B2(n_612), .Y(n_606) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g619 ( .A(n_576), .B(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_578), .A2(n_619), .B1(n_672), .B2(n_675), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g661 ( .A(n_581), .B(n_630), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_581), .B(n_620), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_582), .B(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g695 ( .A(n_582), .B(n_633), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_583), .A2(n_678), .B1(n_691), .B2(n_694), .Y(n_690) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx2_ASAP7_75t_L g599 ( .A(n_584), .Y(n_599) );
AND2x2_ASAP7_75t_L g682 ( .A(n_584), .B(n_604), .Y(n_682) );
OR2x2_ASAP7_75t_L g684 ( .A(n_584), .B(n_651), .Y(n_684) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_584), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_585), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_585), .B(n_630), .Y(n_638) );
OAI211xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_591), .B(n_594), .C(n_606), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_598), .B2(n_601), .C(n_602), .Y(n_594) );
INVxp67_ASAP7_75t_L g706 ( .A(n_597), .Y(n_706) );
INVx1_ASAP7_75t_L g673 ( .A(n_598), .Y(n_673) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g637 ( .A(n_599), .B(n_604), .Y(n_637) );
INVx1_ASAP7_75t_L g654 ( .A(n_600), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_600), .B(n_627), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g669 ( .A(n_604), .Y(n_669) );
AND2x2_ASAP7_75t_L g675 ( .A(n_604), .B(n_630), .Y(n_675) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_SL g663 ( .A(n_611), .Y(n_663) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_614), .B(n_650), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_618), .B2(n_621), .C(n_624), .Y(n_615) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g711 ( .A(n_620), .Y(n_711) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g629 ( .A(n_623), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_627), .B(n_686), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B(n_633), .Y(n_628) );
OAI211xp5_ASAP7_75t_SL g676 ( .A1(n_631), .A2(n_677), .B(n_679), .C(n_685), .Y(n_676) );
INVx1_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g688 ( .A(n_633), .Y(n_688) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI222xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B1(n_648), .B2(n_649), .C1(n_652), .C2(n_653), .Y(n_642) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g718 ( .A(n_649), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_650), .B(n_693), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_650), .A2(n_697), .B1(n_699), .B2(n_702), .Y(n_696) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
NOR4xp25_ASAP7_75t_L g655 ( .A(n_656), .B(n_676), .C(n_689), .D(n_708), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_658), .B(n_688), .Y(n_698) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g665 ( .A(n_663), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_666), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_673), .B(n_674), .Y(n_672) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_696), .C(n_703), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx2_ASAP7_75t_L g705 ( .A(n_701), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
OAI21xp5_ASAP7_75t_SL g712 ( .A1(n_713), .A2(n_715), .B(n_718), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
BUFx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_SL g743 ( .A(n_731), .Y(n_743) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g747 ( .A(n_735), .Y(n_747) );
INVx1_ASAP7_75t_L g740 ( .A(n_737), .Y(n_740) );
BUFx3_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
endmodule