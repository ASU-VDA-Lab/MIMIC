module fake_netlist_5_1131_n_781 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_781);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_781;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_753;
wire n_621;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_779;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_607;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

INVx1_ASAP7_75t_L g158 ( 
.A(n_39),
.Y(n_158)
);

BUFx8_ASAP7_75t_SL g159 ( 
.A(n_18),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_89),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_28),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_17),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_43),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_38),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_68),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_9),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_56),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_26),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_60),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_9),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

BUFx8_ASAP7_75t_SL g178 ( 
.A(n_50),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_33),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_13),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_111),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_62),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_25),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_23),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_12),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_76),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_149),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_87),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_19),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_55),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_37),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_12),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_66),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_67),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_48),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_90),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_84),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_141),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_58),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_31),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_65),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_140),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_53),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_54),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_82),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_34),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_63),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_80),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_1),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_107),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_0),
.Y(n_216)
);

AND2x6_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_20),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_2),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_165),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_3),
.Y(n_223)
);

OAI22x1_ASAP7_75t_SL g224 ( 
.A1(n_187),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_6),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_7),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_158),
.B(n_7),
.Y(n_233)
);

AOI22x1_ASAP7_75t_SL g234 ( 
.A1(n_213),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_234)
);

BUFx8_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_178),
.Y(n_238)
);

BUFx8_ASAP7_75t_SL g239 ( 
.A(n_161),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

CKINVDCx6p67_ASAP7_75t_R g244 ( 
.A(n_186),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_176),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_160),
.B(n_8),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

OAI22x1_ASAP7_75t_SL g251 ( 
.A1(n_180),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_175),
.B(n_14),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_163),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_208),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_188),
.B(n_207),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_217),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

AND2x6_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_177),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_223),
.B(n_164),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_212),
.C(n_211),
.Y(n_269)
);

AOI21x1_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_179),
.B(n_209),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_230),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_230),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_225),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_226),
.A2(n_196),
.B1(n_169),
.B2(n_206),
.Y(n_275)
);

AOI21x1_ASAP7_75t_L g276 ( 
.A1(n_232),
.A2(n_242),
.B(n_237),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_230),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_231),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_231),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_231),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_219),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_231),
.Y(n_283)
);

AOI21x1_ASAP7_75t_L g284 ( 
.A1(n_232),
.A2(n_242),
.B(n_237),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

AO22x2_ASAP7_75t_L g287 ( 
.A1(n_218),
.A2(n_181),
.B1(n_197),
.B2(n_203),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_219),
.B(n_204),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_239),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_256),
.Y(n_298)
);

BUFx6f_ASAP7_75t_SL g299 ( 
.A(n_220),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

AO22x2_ASAP7_75t_L g301 ( 
.A1(n_227),
.A2(n_207),
.B1(n_15),
.B2(n_16),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_256),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_246),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_246),
.B(n_168),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_248),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_243),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_228),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_282),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_276),
.Y(n_309)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_263),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_228),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_276),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_259),
.B(n_227),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_282),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_241),
.Y(n_316)
);

BUFx6f_ASAP7_75t_SL g317 ( 
.A(n_258),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_228),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_269),
.B(n_240),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_263),
.B(n_228),
.Y(n_320)
);

AO221x1_ASAP7_75t_L g321 ( 
.A1(n_301),
.A2(n_287),
.B1(n_303),
.B2(n_221),
.C(n_260),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_265),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_263),
.B(n_220),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_259),
.B(n_216),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_285),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_263),
.B(n_172),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_259),
.B(n_207),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_241),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_284),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_251),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g332 ( 
.A(n_275),
.B(n_252),
.C(n_233),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_266),
.A2(n_252),
.B1(n_233),
.B2(n_222),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_285),
.B(n_207),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_L g335 ( 
.A(n_290),
.B(n_210),
.C(n_184),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_268),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_263),
.B(n_174),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_261),
.B(n_244),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_306),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_263),
.B(n_189),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_286),
.B(n_192),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_274),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_287),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_273),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_294),
.B(n_193),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_268),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_298),
.B(n_198),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_270),
.B(n_207),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_273),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_270),
.B(n_207),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_262),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_300),
.B(n_199),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_262),
.Y(n_354)
);

BUFx6f_ASAP7_75t_SL g355 ( 
.A(n_258),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_268),
.B(n_240),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_289),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_264),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_289),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_277),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_277),
.B(n_200),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_296),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_277),
.B(n_295),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_264),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_267),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_299),
.B(n_235),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_295),
.B(n_243),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_299),
.B(n_235),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_267),
.B(n_202),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_295),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_271),
.B(n_249),
.Y(n_371)
);

NOR3xp33_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_239),
.C(n_287),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_336),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_312),
.B(n_271),
.Y(n_374)
);

OAI21xp33_ASAP7_75t_L g375 ( 
.A1(n_333),
.A2(n_287),
.B(n_301),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_313),
.A2(n_301),
.B(n_302),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_313),
.A2(n_301),
.B(n_302),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_329),
.B(n_258),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_321),
.A2(n_299),
.B1(n_217),
.B2(n_249),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_312),
.B(n_272),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_309),
.A2(n_297),
.B(n_293),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_312),
.B(n_309),
.Y(n_382)
);

BUFx4f_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

AO21x1_ASAP7_75t_L g385 ( 
.A1(n_349),
.A2(n_254),
.B(n_293),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_312),
.B(n_314),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_338),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_314),
.A2(n_330),
.B(n_318),
.Y(n_388)
);

O2A1O1Ixp33_ASAP7_75t_L g389 ( 
.A1(n_344),
.A2(n_325),
.B(n_349),
.C(n_351),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_330),
.B(n_272),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_338),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_324),
.B(n_278),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_324),
.B(n_278),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_325),
.A2(n_297),
.B(n_292),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_351),
.A2(n_292),
.B(n_291),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_311),
.A2(n_323),
.B(n_328),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_316),
.A2(n_217),
.B1(n_254),
.B2(n_224),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_343),
.B(n_279),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_367),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_317),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_328),
.A2(n_291),
.B(n_288),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_361),
.A2(n_288),
.B(n_283),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_345),
.B(n_279),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_363),
.A2(n_283),
.B(n_280),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_350),
.B(n_280),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_319),
.B(n_217),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_371),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_315),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_334),
.B(n_234),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_357),
.B(n_217),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_336),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_359),
.B(n_21),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_356),
.B(n_14),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_339),
.B(n_15),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_334),
.B(n_16),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_307),
.B(n_22),
.Y(n_417)
);

AOI21x1_ASAP7_75t_L g418 ( 
.A1(n_371),
.A2(n_99),
.B(n_155),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_340),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_342),
.B(n_17),
.Y(n_421)
);

O2A1O1Ixp33_ASAP7_75t_SL g422 ( 
.A1(n_327),
.A2(n_18),
.B(n_19),
.C(n_24),
.Y(n_422)
);

BUFx12f_ASAP7_75t_L g423 ( 
.A(n_317),
.Y(n_423)
);

AO21x1_ASAP7_75t_L g424 ( 
.A1(n_369),
.A2(n_27),
.B(n_29),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_346),
.A2(n_30),
.B(n_32),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_347),
.B(n_35),
.Y(n_426)
);

NOR3xp33_ASAP7_75t_L g427 ( 
.A(n_362),
.B(n_36),
.C(n_40),
.Y(n_427)
);

A2O1A1Ixp33_ASAP7_75t_L g428 ( 
.A1(n_360),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_348),
.B(n_45),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_337),
.A2(n_46),
.B(n_47),
.Y(n_430)
);

NOR2x2_ASAP7_75t_L g431 ( 
.A(n_331),
.B(n_49),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_347),
.B(n_51),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_341),
.A2(n_310),
.B(n_320),
.Y(n_433)
);

NAND3xp33_ASAP7_75t_L g434 ( 
.A(n_369),
.B(n_52),
.C(n_57),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_352),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_353),
.A2(n_310),
.B(n_370),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_310),
.A2(n_59),
.B(n_61),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_352),
.Y(n_438)
);

AOI21x1_ASAP7_75t_L g439 ( 
.A1(n_354),
.A2(n_365),
.B(n_364),
.Y(n_439)
);

NOR3xp33_ASAP7_75t_L g440 ( 
.A(n_366),
.B(n_64),
.C(n_69),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_347),
.B(n_70),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_375),
.A2(n_355),
.B1(n_368),
.B2(n_366),
.Y(n_442)
);

NAND2x1p5_ASAP7_75t_L g443 ( 
.A(n_373),
.B(n_354),
.Y(n_443)
);

OAI21x1_ASAP7_75t_L g444 ( 
.A1(n_439),
.A2(n_365),
.B(n_364),
.Y(n_444)
);

AO31x2_ASAP7_75t_L g445 ( 
.A1(n_385),
.A2(n_358),
.A3(n_368),
.B(n_335),
.Y(n_445)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_388),
.A2(n_358),
.B(n_72),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_382),
.B(n_71),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_386),
.B(n_73),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_381),
.A2(n_75),
.B(n_77),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_436),
.A2(n_78),
.B(n_79),
.Y(n_451)
);

AOI21x1_ASAP7_75t_L g452 ( 
.A1(n_374),
.A2(n_81),
.B(n_83),
.Y(n_452)
);

AOI21x1_ASAP7_75t_L g453 ( 
.A1(n_380),
.A2(n_86),
.B(n_88),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_409),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_436),
.A2(n_91),
.B(n_92),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_423),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_376),
.A2(n_355),
.B(n_94),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_393),
.B(n_93),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_416),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_400),
.B(n_95),
.Y(n_460)
);

AO31x2_ASAP7_75t_L g461 ( 
.A1(n_376),
.A2(n_377),
.A3(n_424),
.B(n_421),
.Y(n_461)
);

INVx6_ASAP7_75t_SL g462 ( 
.A(n_383),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_377),
.A2(n_389),
.B(n_390),
.Y(n_463)
);

O2A1O1Ixp5_ASAP7_75t_L g464 ( 
.A1(n_397),
.A2(n_96),
.B(n_97),
.C(n_98),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_408),
.B(n_100),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_396),
.A2(n_101),
.B(n_102),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_417),
.B(n_103),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_415),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_420),
.B(n_104),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_387),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_412),
.B(n_105),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_414),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_412),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_378),
.B(n_106),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_391),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_419),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g477 ( 
.A1(n_396),
.A2(n_108),
.B(n_109),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_373),
.B(n_110),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_395),
.A2(n_156),
.B(n_113),
.Y(n_479)
);

OAI21x1_ASAP7_75t_L g480 ( 
.A1(n_395),
.A2(n_154),
.B(n_114),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_433),
.A2(n_112),
.B(n_115),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_429),
.B(n_116),
.Y(n_482)
);

AOI21x1_ASAP7_75t_L g483 ( 
.A1(n_402),
.A2(n_117),
.B(n_118),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_438),
.B(n_119),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_392),
.A2(n_120),
.B(n_121),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_383),
.Y(n_486)
);

AOI211x1_ASAP7_75t_L g487 ( 
.A1(n_430),
.A2(n_153),
.B(n_123),
.C(n_124),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_372),
.B(n_122),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_403),
.A2(n_150),
.B(n_127),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_405),
.A2(n_148),
.B(n_128),
.Y(n_490)
);

A2O1A1Ixp33_ASAP7_75t_L g491 ( 
.A1(n_379),
.A2(n_126),
.B(n_129),
.C(n_131),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_394),
.B(n_132),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_435),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_404),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_411),
.A2(n_133),
.B(n_134),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_398),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_399),
.A2(n_135),
.B(n_136),
.Y(n_497)
);

OAI21x1_ASAP7_75t_SL g498 ( 
.A1(n_413),
.A2(n_137),
.B(n_143),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_446),
.A2(n_441),
.B(n_432),
.Y(n_499)
);

OAI21x1_ASAP7_75t_SL g500 ( 
.A1(n_498),
.A2(n_437),
.B(n_418),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_449),
.A2(n_426),
.B(n_437),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_450),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_479),
.A2(n_480),
.B(n_477),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_456),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_410),
.Y(n_505)
);

AO21x2_ASAP7_75t_L g506 ( 
.A1(n_481),
.A2(n_406),
.B(n_407),
.Y(n_506)
);

NAND2x1p5_ASAP7_75t_L g507 ( 
.A(n_473),
.B(n_425),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_451),
.A2(n_434),
.B(n_422),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_448),
.A2(n_447),
.B(n_463),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_444),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_493),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_496),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_473),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_454),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_455),
.A2(n_428),
.B(n_440),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_468),
.B(n_401),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_471),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_489),
.A2(n_427),
.B(n_146),
.Y(n_518)
);

NAND2x1p5_ASAP7_75t_L g519 ( 
.A(n_473),
.B(n_144),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_459),
.B(n_147),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_490),
.A2(n_483),
.B(n_463),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_470),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_448),
.A2(n_431),
.B(n_478),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_475),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_465),
.A2(n_481),
.B(n_482),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_452),
.Y(n_526)
);

OAI21x1_ASAP7_75t_SL g527 ( 
.A1(n_466),
.A2(n_457),
.B(n_458),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_442),
.Y(n_528)
);

INVx5_ASAP7_75t_L g529 ( 
.A(n_471),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_453),
.A2(n_469),
.B(n_464),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_457),
.A2(n_466),
.B(n_465),
.Y(n_531)
);

OA21x2_ASAP7_75t_L g532 ( 
.A1(n_469),
.A2(n_482),
.B(n_491),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_492),
.A2(n_443),
.B(n_484),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_443),
.A2(n_495),
.B(n_485),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_459),
.B(n_472),
.Y(n_535)
);

AO21x2_ASAP7_75t_L g536 ( 
.A1(n_460),
.A2(n_497),
.B(n_467),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_461),
.B(n_488),
.Y(n_537)
);

AO21x1_ASAP7_75t_L g538 ( 
.A1(n_442),
.A2(n_488),
.B(n_487),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_486),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_476),
.A2(n_474),
.B(n_445),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_445),
.A2(n_461),
.B(n_462),
.Y(n_541)
);

OA21x2_ASAP7_75t_L g542 ( 
.A1(n_461),
.A2(n_445),
.B(n_462),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_450),
.Y(n_543)
);

AO31x2_ASAP7_75t_L g544 ( 
.A1(n_491),
.A2(n_385),
.A3(n_424),
.B(n_377),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g545 ( 
.A(n_473),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_510),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_537),
.B(n_505),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_513),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_543),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_510),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_503),
.A2(n_521),
.B(n_534),
.Y(n_551)
);

OAI21x1_ASAP7_75t_L g552 ( 
.A1(n_503),
.A2(n_521),
.B(n_534),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_502),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_511),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_511),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_513),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_522),
.Y(n_557)
);

INVxp33_ASAP7_75t_SL g558 ( 
.A(n_516),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_526),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_529),
.B(n_535),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_504),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_517),
.B(n_529),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_525),
.A2(n_540),
.B(n_509),
.Y(n_563)
);

BUFx8_ASAP7_75t_SL g564 ( 
.A(n_504),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_524),
.Y(n_565)
);

AO21x2_ASAP7_75t_L g566 ( 
.A1(n_527),
.A2(n_500),
.B(n_530),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_526),
.Y(n_567)
);

AOI21x1_ASAP7_75t_L g568 ( 
.A1(n_530),
.A2(n_532),
.B(n_501),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_526),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_541),
.Y(n_570)
);

CKINVDCx14_ASAP7_75t_R g571 ( 
.A(n_512),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_541),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_533),
.A2(n_501),
.B(n_508),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_540),
.Y(n_574)
);

NAND2x1p5_ASAP7_75t_L g575 ( 
.A(n_529),
.B(n_513),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_544),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_542),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_514),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_542),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_513),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_517),
.B(n_529),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_542),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_533),
.A2(n_508),
.B(n_499),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_512),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_528),
.A2(n_531),
.B1(n_537),
.B2(n_545),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_544),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_544),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_538),
.A2(n_523),
.B1(n_531),
.B2(n_520),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_531),
.B(n_544),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_547),
.B(n_523),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_558),
.A2(n_539),
.B1(n_532),
.B2(n_519),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_547),
.B(n_519),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_554),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_585),
.B(n_532),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_553),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_553),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_578),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_549),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_556),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_555),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_549),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_546),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_546),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_557),
.B(n_506),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_546),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_557),
.B(n_506),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_565),
.B(n_518),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_560),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_589),
.B(n_518),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_565),
.B(n_515),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_587),
.B(n_515),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_562),
.B(n_539),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_507),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_588),
.B(n_507),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_584),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_562),
.B(n_536),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_548),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_562),
.B(n_536),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_571),
.A2(n_499),
.B1(n_562),
.B2(n_581),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_SL g620 ( 
.A1(n_563),
.A2(n_581),
.B(n_575),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_550),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_581),
.B(n_559),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_576),
.B(n_586),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_589),
.B(n_586),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_576),
.B(n_586),
.Y(n_625)
);

AND2x4_ASAP7_75t_SL g626 ( 
.A(n_556),
.B(n_581),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_550),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_576),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_548),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_SL g630 ( 
.A1(n_561),
.A2(n_548),
.B1(n_556),
.B2(n_575),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_566),
.A2(n_564),
.B1(n_570),
.B2(n_572),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_577),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_577),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_559),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_632),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_590),
.B(n_582),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_595),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_590),
.B(n_582),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_632),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_602),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_602),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_591),
.A2(n_566),
.B1(n_556),
.B2(n_580),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_608),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_608),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_598),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_633),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_613),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_633),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g649 ( 
.A(n_595),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_604),
.B(n_579),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_625),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_612),
.B(n_580),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_604),
.B(n_579),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_624),
.B(n_625),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_603),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_624),
.B(n_566),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_597),
.B(n_569),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_603),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_615),
.B(n_569),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_628),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_630),
.A2(n_580),
.B1(n_575),
.B2(n_572),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_592),
.A2(n_580),
.B1(n_570),
.B2(n_567),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_601),
.B(n_569),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_628),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_606),
.B(n_574),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_609),
.B(n_574),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_623),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_592),
.B(n_567),
.Y(n_668)
);

NOR2x1_ASAP7_75t_SL g669 ( 
.A(n_620),
.B(n_567),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_596),
.B(n_568),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_606),
.B(n_610),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_671),
.B(n_611),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_652),
.B(n_619),
.C(n_631),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_647),
.B(n_667),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_671),
.B(n_611),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_654),
.B(n_616),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_656),
.B(n_594),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_635),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_643),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_645),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_643),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_635),
.Y(n_682)
);

NAND2x1p5_ASAP7_75t_L g683 ( 
.A(n_644),
.B(n_613),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_639),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_647),
.B(n_610),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_667),
.B(n_618),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_656),
.B(n_670),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_645),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_657),
.B(n_596),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_639),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_636),
.B(n_623),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_659),
.B(n_598),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_637),
.B(n_622),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_644),
.B(n_607),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_648),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_648),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_679),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_690),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_672),
.B(n_638),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_690),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_678),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_688),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_674),
.B(n_669),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_682),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_672),
.B(n_638),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_692),
.B(n_649),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_681),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_684),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_695),
.Y(n_709)
);

NAND4xp75_ASAP7_75t_L g710 ( 
.A(n_689),
.B(n_661),
.C(n_642),
.D(n_663),
.Y(n_710)
);

AOI211xp5_ASAP7_75t_L g711 ( 
.A1(n_710),
.A2(n_673),
.B(n_693),
.C(n_594),
.Y(n_711)
);

AND2x2_ASAP7_75t_SL g712 ( 
.A(n_703),
.B(n_674),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_701),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_702),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_706),
.B(n_687),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_SL g716 ( 
.A1(n_707),
.A2(n_669),
.B(n_680),
.Y(n_716)
);

OAI22xp33_ASAP7_75t_L g717 ( 
.A1(n_710),
.A2(n_683),
.B1(n_677),
.B2(n_676),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_701),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_704),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_700),
.Y(n_720)
);

AOI32xp33_ASAP7_75t_L g721 ( 
.A1(n_703),
.A2(n_674),
.A3(n_685),
.B1(n_686),
.B2(n_675),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_712),
.B(n_705),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_711),
.A2(n_703),
.B(n_708),
.Y(n_723)
);

AOI22x1_ASAP7_75t_L g724 ( 
.A1(n_714),
.A2(n_697),
.B1(n_680),
.B2(n_683),
.Y(n_724)
);

AOI211xp5_ASAP7_75t_L g725 ( 
.A1(n_717),
.A2(n_687),
.B(n_697),
.C(n_694),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_711),
.A2(n_668),
.B(n_677),
.Y(n_726)
);

AOI222xp33_ASAP7_75t_L g727 ( 
.A1(n_723),
.A2(n_717),
.B1(n_686),
.B2(n_719),
.C1(n_718),
.C2(n_713),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_722),
.B(n_715),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_726),
.B(n_721),
.Y(n_729)
);

AOI211xp5_ASAP7_75t_L g730 ( 
.A1(n_725),
.A2(n_716),
.B(n_698),
.C(n_686),
.Y(n_730)
);

AOI211x1_ASAP7_75t_L g731 ( 
.A1(n_724),
.A2(n_705),
.B(n_699),
.C(n_675),
.Y(n_731)
);

AOI221xp5_ASAP7_75t_L g732 ( 
.A1(n_723),
.A2(n_720),
.B1(n_709),
.B2(n_704),
.C(n_699),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_729),
.B(n_709),
.Y(n_733)
);

NOR4xp25_ASAP7_75t_L g734 ( 
.A(n_732),
.B(n_700),
.C(n_696),
.D(n_607),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_731),
.B(n_691),
.Y(n_735)
);

AOI211xp5_ASAP7_75t_L g736 ( 
.A1(n_730),
.A2(n_614),
.B(n_617),
.C(n_629),
.Y(n_736)
);

NAND4xp25_ASAP7_75t_SL g737 ( 
.A(n_727),
.B(n_685),
.C(n_691),
.D(n_662),
.Y(n_737)
);

OAI322xp33_ASAP7_75t_L g738 ( 
.A1(n_733),
.A2(n_728),
.A3(n_646),
.B1(n_666),
.B2(n_664),
.C1(n_660),
.C2(n_654),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_735),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_737),
.A2(n_614),
.B1(n_617),
.B2(n_636),
.Y(n_740)
);

NOR2x1_ASAP7_75t_L g741 ( 
.A(n_738),
.B(n_736),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_739),
.B(n_617),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_740),
.B(n_734),
.Y(n_743)
);

NAND4xp75_ASAP7_75t_L g744 ( 
.A(n_741),
.B(n_665),
.C(n_664),
.D(n_660),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_742),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_743),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_742),
.B(n_617),
.Y(n_747)
);

NAND4xp75_ASAP7_75t_L g748 ( 
.A(n_741),
.B(n_665),
.C(n_653),
.D(n_650),
.Y(n_748)
);

XNOR2xp5_ASAP7_75t_L g749 ( 
.A(n_741),
.B(n_626),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_746),
.A2(n_617),
.B1(n_626),
.B2(n_650),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_745),
.B(n_653),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_747),
.Y(n_752)
);

NOR2x1_ASAP7_75t_L g753 ( 
.A(n_744),
.B(n_599),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_747),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_748),
.A2(n_641),
.B1(n_658),
.B2(n_655),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_749),
.Y(n_756)
);

AO22x2_ASAP7_75t_L g757 ( 
.A1(n_752),
.A2(n_599),
.B1(n_658),
.B2(n_655),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_751),
.Y(n_758)
);

OA21x2_ASAP7_75t_L g759 ( 
.A1(n_754),
.A2(n_583),
.B(n_573),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_756),
.A2(n_641),
.B1(n_640),
.B2(n_599),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_750),
.B(n_666),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_753),
.A2(n_651),
.B1(n_640),
.B2(n_609),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_758),
.Y(n_763)
);

XOR2xp5_ASAP7_75t_L g764 ( 
.A(n_760),
.B(n_762),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_759),
.Y(n_765)
);

XNOR2xp5_ASAP7_75t_L g766 ( 
.A(n_761),
.B(n_755),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_757),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_758),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_758),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_763),
.A2(n_651),
.B1(n_621),
.B2(n_634),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_768),
.A2(n_769),
.B1(n_763),
.B2(n_766),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_764),
.A2(n_583),
.B(n_573),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_767),
.A2(n_551),
.B(n_552),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_765),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_774),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_771),
.B(n_651),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_775),
.B(n_770),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_776),
.A2(n_772),
.B(n_773),
.Y(n_778)
);

XNOR2xp5_ASAP7_75t_L g779 ( 
.A(n_777),
.B(n_568),
.Y(n_779)
);

AOI221xp5_ASAP7_75t_L g780 ( 
.A1(n_779),
.A2(n_778),
.B1(n_627),
.B2(n_605),
.C(n_600),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_780),
.A2(n_627),
.B1(n_605),
.B2(n_593),
.Y(n_781)
);


endmodule