module fake_jpeg_14383_n_266 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_266);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_266;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_155;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_25),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_47),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_50),
.B(n_59),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_4),
.C(n_5),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_26),
.Y(n_109)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g93 ( 
.A(n_54),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_79),
.Y(n_91)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_21),
.B(n_4),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_22),
.B(n_33),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_70),
.Y(n_103)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_66),
.Y(n_105)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_22),
.B(n_33),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_75),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_23),
.A2(n_36),
.B(n_35),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_31),
.C(n_36),
.Y(n_99)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_23),
.B(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_84),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_41),
.Y(n_83)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_32),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_99),
.B(n_112),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_SL g102 ( 
.A(n_80),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_102),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_32),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_104),
.B(n_109),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_47),
.B(n_27),
.C(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_25),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_52),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_69),
.A2(n_38),
.B1(n_17),
.B2(n_29),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_55),
.B1(n_34),
.B2(n_81),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_121),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_65),
.B(n_35),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_126),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_44),
.A2(n_17),
.B1(n_34),
.B2(n_8),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_124),
.A2(n_123),
.B1(n_89),
.B2(n_106),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_5),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_5),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_7),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_83),
.B1(n_60),
.B2(n_46),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_131),
.A2(n_164),
.B1(n_169),
.B2(n_155),
.Y(n_194)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_134),
.B(n_139),
.Y(n_189)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_135),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_58),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_136),
.B(n_137),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_127),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_68),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_155),
.Y(n_170)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

AO22x2_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_54),
.B1(n_48),
.B2(n_51),
.Y(n_141)
);

AO22x1_ASAP7_75t_SL g186 ( 
.A1(n_141),
.A2(n_133),
.B1(n_150),
.B2(n_167),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_81),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_146),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_152),
.B1(n_158),
.B2(n_86),
.Y(n_173)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_97),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_95),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_151),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_7),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_156),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_91),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_109),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_93),
.A2(n_9),
.B(n_10),
.C(n_118),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_159),
.B(n_163),
.Y(n_193)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_111),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_162),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_89),
.A2(n_10),
.B1(n_106),
.B2(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_105),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_160),
.B(n_161),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_123),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_93),
.B(n_86),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_167),
.B(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_107),
.A2(n_125),
.B1(n_119),
.B2(n_93),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_115),
.B(n_116),
.C(n_121),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g213 ( 
.A1(n_171),
.A2(n_196),
.B(n_193),
.C(n_181),
.D(n_184),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_164),
.B1(n_165),
.B2(n_154),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_180),
.B1(n_187),
.B2(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_173),
.B(n_194),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_110),
.B1(n_115),
.B2(n_138),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_160),
.A2(n_115),
.B(n_110),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_198),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_141),
.A2(n_156),
.B1(n_166),
.B2(n_161),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_186),
.B1(n_194),
.B2(n_170),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_140),
.A2(n_159),
.B1(n_168),
.B2(n_144),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_138),
.A2(n_166),
.B1(n_148),
.B2(n_163),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_153),
.C(n_135),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_145),
.A2(n_132),
.B(n_144),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_157),
.C(n_177),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_202),
.A2(n_213),
.B(n_186),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_175),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_198),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_212),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_174),
.B1(n_195),
.B2(n_197),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_216),
.B1(n_182),
.B2(n_190),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_196),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_185),
.Y(n_209)
);

AOI322xp5_ASAP7_75t_SL g223 ( 
.A1(n_209),
.A2(n_176),
.A3(n_179),
.B1(n_182),
.B2(n_190),
.C1(n_191),
.C2(n_205),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_183),
.B(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_191),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_217),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_173),
.A2(n_186),
.B1(n_170),
.B2(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_216),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_223),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_170),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_228),
.C(n_230),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_199),
.B(n_206),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_179),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_205),
.C(n_209),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_213),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_224),
.Y(n_249)
);

NOR2xp67_ASAP7_75t_SL g233 ( 
.A(n_219),
.B(n_201),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_241),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_235),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_199),
.B(n_217),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_236),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_215),
.B(n_211),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_211),
.B(n_229),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_246),
.B(n_249),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_232),
.B(n_228),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_239),
.B1(n_225),
.B2(n_240),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_251),
.B1(n_234),
.B2(n_245),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_225),
.B1(n_240),
.B2(n_236),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_247),
.B(n_242),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_252),
.B(n_221),
.Y(n_258)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_221),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_243),
.C(n_246),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_257),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_256),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_231),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_251),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_250),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_259),
.C(n_260),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_255),
.Y(n_266)
);


endmodule