module fake_netlist_1_6579_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_7), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g14 ( .A(n_8), .B(n_9), .Y(n_14) );
BUFx3_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
BUFx3_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_12), .Y(n_18) );
AOI21xp33_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_0), .B(n_2), .Y(n_19) );
O2A1O1Ixp33_ASAP7_75t_L g20 ( .A1(n_11), .A2(n_2), .B(n_3), .C(n_4), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_16), .A2(n_3), .B(n_4), .Y(n_21) );
BUFx2_ASAP7_75t_L g22 ( .A(n_15), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_17), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_13), .B1(n_11), .B2(n_17), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_21), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_20), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_23), .B(n_18), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_23), .B(n_12), .Y(n_29) );
OAI32xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_25), .A3(n_15), .B1(n_17), .B2(n_26), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_26), .B1(n_24), .B2(n_19), .Y(n_31) );
O2A1O1Ixp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_29), .B(n_19), .C(n_13), .Y(n_32) );
OAI211xp5_ASAP7_75t_SL g33 ( .A1(n_31), .A2(n_14), .B(n_15), .C(n_17), .Y(n_33) );
INVx2_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
XNOR2x1_ASAP7_75t_L g35 ( .A(n_33), .B(n_5), .Y(n_35) );
AOI22x1_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_15), .B1(n_14), .B2(n_7), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_35), .B1(n_34), .B2(n_5), .Y(n_37) );
endmodule