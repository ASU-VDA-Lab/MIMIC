module fake_netlist_6_1791_n_549 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_55, n_94, n_97, n_108, n_58, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_103, n_111, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_549);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_94;
input n_97;
input n_108;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_549;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_507;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_148;
wire n_208;
wire n_161;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_495;
wire n_350;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_114;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_119;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_529;
wire n_445;
wire n_425;
wire n_122;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_490;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_154;
wire n_456;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_513;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_121;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_477;
wire n_533;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_124;
wire n_548;
wire n_282;
wire n_436;
wire n_116;
wire n_211;
wire n_523;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_123;
wire n_136;
wire n_546;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_487;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_17),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_32),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_5),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_41),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_5),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_75),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_12),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_97),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_103),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_50),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_45),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_57),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_26),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_56),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_25),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_14),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_27),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_53),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_59),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_8),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_30),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_63),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_21),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_37),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_31),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_52),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_16),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_29),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_67),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_89),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_43),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_84),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_33),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_54),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_11),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_61),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_10),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_15),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_65),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_1),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_116),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_123),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_114),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_128),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_134),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_119),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_136),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_118),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_137),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_139),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_147),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_124),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_0),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_149),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_151),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_152),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_135),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_141),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_153),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_156),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_143),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_143),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_131),
.B(n_163),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_161),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_173),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

NAND2xp33_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_122),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_172),
.B(n_129),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_179),
.B(n_160),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_180),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_SL g247 ( 
.A(n_197),
.B(n_122),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_205),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_203),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_195),
.Y(n_252)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_178),
.B(n_122),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_184),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_169),
.C(n_168),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_158),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

AND2x6_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_121),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_213),
.B(n_159),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_224),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_228),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_219),
.B(n_142),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_212),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_212),
.B(n_140),
.Y(n_271)
);

BUFx4f_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_127),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_225),
.Y(n_274)
);

NAND3x1_ASAP7_75t_L g275 ( 
.A(n_213),
.B(n_167),
.C(n_162),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_211),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_226),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_226),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_212),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_234),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_235),
.B(n_164),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_214),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_216),
.B(n_148),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_217),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_217),
.B(n_150),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_253),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_227),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_230),
.B(n_165),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_221),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_132),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_223),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_240),
.B(n_243),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_255),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_231),
.B(n_138),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_230),
.B(n_245),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_236),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_246),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_238),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_252),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_145),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_253),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_241),
.B(n_154),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_254),
.Y(n_311)
);

OAI221xp5_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_247),
.B1(n_242),
.B2(n_249),
.C(n_248),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_218),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

AO22x2_ASAP7_75t_L g315 ( 
.A1(n_296),
.A2(n_251),
.B1(n_215),
.B2(n_244),
.Y(n_315)
);

BUFx6f_ASAP7_75t_SL g316 ( 
.A(n_293),
.Y(n_316)
);

BUFx8_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_269),
.Y(n_319)
);

AO22x2_ASAP7_75t_L g320 ( 
.A1(n_299),
.A2(n_251),
.B1(n_253),
.B2(n_3),
.Y(n_320)
);

AO22x2_ASAP7_75t_L g321 ( 
.A1(n_276),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_321)
);

AND2x6_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_254),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_272),
.B(n_2),
.Y(n_323)
);

AO22x2_ASAP7_75t_L g324 ( 
.A1(n_276),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_324)
);

OAI221xp5_ASAP7_75t_L g325 ( 
.A1(n_300),
.A2(n_285),
.B1(n_310),
.B2(n_286),
.C(n_305),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_266),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_267),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_13),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_270),
.B(n_18),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_272),
.B(n_4),
.Y(n_332)
);

BUFx8_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

AO22x2_ASAP7_75t_L g334 ( 
.A1(n_297),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_274),
.Y(n_335)
);

OR2x6_ASAP7_75t_L g336 ( 
.A(n_259),
.B(n_9),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_279),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_280),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_283),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_281),
.B(n_112),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_288),
.B(n_19),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_268),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_268),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_20),
.Y(n_344)
);

BUFx8_ASAP7_75t_L g345 ( 
.A(n_307),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_298),
.B(n_66),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_264),
.B(n_9),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_297),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_298),
.A2(n_69),
.B1(n_22),
.B2(n_23),
.Y(n_349)
);

AO21x1_ASAP7_75t_L g350 ( 
.A1(n_271),
.A2(n_10),
.B(n_24),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_256),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_263),
.Y(n_352)
);

HAxp5_ASAP7_75t_SL g353 ( 
.A(n_275),
.B(n_34),
.CON(n_353),
.SN(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_306),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_273),
.Y(n_355)
);

AO22x2_ASAP7_75t_L g356 ( 
.A1(n_306),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_289),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_289),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_292),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_359)
);

NAND2xp33_ASAP7_75t_SL g360 ( 
.A(n_313),
.B(n_281),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_318),
.B(n_284),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_287),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_354),
.B(n_287),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_347),
.B(n_304),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_290),
.Y(n_365)
);

NOR2x1_ASAP7_75t_L g366 ( 
.A(n_311),
.B(n_292),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_269),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_SL g368 ( 
.A(n_316),
.B(n_309),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_291),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_309),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_346),
.B(n_304),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_314),
.B(n_291),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_341),
.B(n_304),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_326),
.B(n_282),
.Y(n_374)
);

NAND2xp33_ASAP7_75t_SL g375 ( 
.A(n_332),
.B(n_260),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_323),
.B(n_258),
.Y(n_376)
);

NAND2xp33_ASAP7_75t_SL g377 ( 
.A(n_319),
.B(n_271),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_343),
.B(n_262),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_327),
.B(n_261),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_355),
.B(n_257),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_351),
.B(n_257),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_315),
.B(n_44),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_335),
.B(n_329),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_337),
.B(n_47),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_338),
.B(n_48),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_328),
.B(n_330),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_344),
.B(n_51),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_340),
.B(n_55),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_315),
.B(n_60),
.Y(n_389)
);

NAND2xp33_ASAP7_75t_SL g390 ( 
.A(n_353),
.B(n_331),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_352),
.B(n_62),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_349),
.B(n_64),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_386),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_374),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_363),
.B(n_345),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_370),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_322),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_372),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

BUFx10_ASAP7_75t_L g400 ( 
.A(n_368),
.Y(n_400)
);

OAI21x1_ASAP7_75t_L g401 ( 
.A1(n_383),
.A2(n_359),
.B(n_350),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_367),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_369),
.A2(n_325),
.B1(n_356),
.B2(n_312),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_362),
.B(n_322),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_378),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_382),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_379),
.Y(n_407)
);

AO31x2_ASAP7_75t_L g408 ( 
.A1(n_385),
.A2(n_320),
.A3(n_356),
.B(n_324),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_377),
.A2(n_360),
.B(n_373),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_380),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_392),
.A2(n_322),
.B(n_336),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_371),
.A2(n_320),
.B(n_336),
.Y(n_412)
);

A2O1A1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_390),
.A2(n_324),
.B(n_321),
.C(n_334),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_366),
.B(n_70),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_321),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_389),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_392),
.A2(n_334),
.B(n_72),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_376),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_410),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_402),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_418),
.B(n_361),
.Y(n_421)
);

OR2x6_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_391),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_394),
.Y(n_423)
);

NAND3xp33_ASAP7_75t_L g424 ( 
.A(n_417),
.B(n_375),
.C(n_333),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_417),
.B(n_412),
.C(n_413),
.Y(n_425)
);

AO21x2_ASAP7_75t_L g426 ( 
.A1(n_401),
.A2(n_364),
.B(n_387),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_387),
.Y(n_427)
);

INVx4_ASAP7_75t_SL g428 ( 
.A(n_397),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_409),
.A2(n_388),
.B(n_384),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_393),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_403),
.A2(n_416),
.B1(n_411),
.B2(n_415),
.Y(n_431)
);

CKINVDCx11_ASAP7_75t_R g432 ( 
.A(n_400),
.Y(n_432)
);

OAI22xp33_ASAP7_75t_L g433 ( 
.A1(n_415),
.A2(n_416),
.B1(n_406),
.B2(n_403),
.Y(n_433)
);

A2O1A1Ixp33_ASAP7_75t_L g434 ( 
.A1(n_399),
.A2(n_71),
.B(n_73),
.C(n_74),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_405),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_396),
.B(n_76),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_407),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_404),
.A2(n_77),
.B(n_78),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_396),
.Y(n_439)
);

BUFx12f_ASAP7_75t_L g440 ( 
.A(n_400),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_430),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_423),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_423),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_419),
.Y(n_444)
);

AND2x4_ASAP7_75t_SL g445 ( 
.A(n_439),
.B(n_397),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_420),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_419),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_429),
.A2(n_408),
.B(n_414),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_396),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_437),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_424),
.A2(n_414),
.B1(n_317),
.B2(n_408),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_437),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_425),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_439),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_408),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_435),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_433),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_427),
.B(n_79),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_426),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_426),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_440),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_433),
.B(n_82),
.Y(n_462)
);

AO32x2_ASAP7_75t_L g463 ( 
.A1(n_431),
.A2(n_85),
.A3(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_463)
);

OR2x6_ASAP7_75t_L g464 ( 
.A(n_422),
.B(n_90),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_422),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_431),
.B(n_98),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_432),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_428),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_464),
.B(n_428),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_441),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_421),
.Y(n_471)
);

CKINVDCx11_ASAP7_75t_R g472 ( 
.A(n_461),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_R g473 ( 
.A(n_446),
.B(n_438),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_465),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_R g475 ( 
.A(n_464),
.B(n_432),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_452),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_456),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_459),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_R g479 ( 
.A(n_461),
.B(n_440),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_428),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_452),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_454),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_445),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_451),
.B(n_100),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_445),
.B(n_434),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_R g486 ( 
.A(n_455),
.B(n_102),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_442),
.B(n_434),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_R g488 ( 
.A(n_453),
.B(n_110),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_443),
.B(n_104),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_444),
.B(n_109),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_478),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_470),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_453),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_478),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_468),
.B(n_460),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_482),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_476),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_457),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_480),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_457),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_R g501 ( 
.A(n_475),
.B(n_462),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_468),
.B(n_460),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_485),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_451),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_447),
.Y(n_505)
);

AND2x4_ASAP7_75t_SL g506 ( 
.A(n_495),
.B(n_469),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_492),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_496),
.Y(n_508)
);

OAI33xp33_ASAP7_75t_L g509 ( 
.A1(n_498),
.A2(n_466),
.A3(n_458),
.B1(n_463),
.B2(n_473),
.B3(n_450),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g510 ( 
.A1(n_501),
.A2(n_484),
.B1(n_462),
.B2(n_504),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_459),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_495),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_471),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_507),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_508),
.B(n_500),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_511),
.B(n_491),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_512),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_495),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_503),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_513),
.B(n_491),
.Y(n_520)
);

NOR2x1_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_505),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_472),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_497),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_517),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_516),
.B(n_502),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_523),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_525),
.B(n_524),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_518),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_522),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_518),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_526),
.B(n_510),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_527),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_528),
.B(n_519),
.Y(n_533)
);

CKINVDCx6p67_ASAP7_75t_R g534 ( 
.A(n_532),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_529),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_534),
.Y(n_536)
);

NOR3xp33_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_535),
.C(n_533),
.Y(n_537)
);

AOI32xp33_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_528),
.A3(n_530),
.B1(n_501),
.B2(n_469),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_479),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_SL g540 ( 
.A(n_539),
.B(n_488),
.Y(n_540)
);

AOI221xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_509),
.B1(n_486),
.B2(n_490),
.C(n_489),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_541),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_542),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_543),
.A2(n_509),
.B1(n_490),
.B2(n_483),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_105),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_545),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_546),
.Y(n_547)
);

AOI221xp5_ASAP7_75t_L g548 ( 
.A1(n_547),
.A2(n_485),
.B1(n_107),
.B2(n_494),
.C(n_502),
.Y(n_548)
);

AOI211xp5_ASAP7_75t_L g549 ( 
.A1(n_548),
.A2(n_463),
.B(n_448),
.C(n_494),
.Y(n_549)
);


endmodule