module fake_jpeg_9460_n_278 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_39),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_31),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_50),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_22),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_27),
.C(n_19),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_23),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_33),
.B1(n_41),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_49),
.A2(n_66),
.B1(n_21),
.B2(n_19),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_33),
.B1(n_23),
.B2(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_30),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_63),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_24),
.B1(n_29),
.B2(n_20),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_24),
.B1(n_29),
.B2(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_58),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_27),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_29),
.B1(n_25),
.B2(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_32),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_23),
.B1(n_18),
.B2(n_19),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_89),
.Y(n_105)
);

AO22x2_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_23),
.B1(n_43),
.B2(n_31),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_85),
.B1(n_88),
.B2(n_51),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_74),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_32),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_71),
.B(n_76),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_78),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_26),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_81),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_26),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_84),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_25),
.B1(n_21),
.B2(n_43),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_90),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_63),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_1),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_48),
.B(n_1),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_27),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_27),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_45),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_57),
.Y(n_99)
);

INVx2_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_58),
.A2(n_50),
.B(n_61),
.C(n_64),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_18),
.B(n_37),
.Y(n_122)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_37),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_110),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_124),
.B1(n_101),
.B2(n_80),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_98),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_127),
.B(n_18),
.C(n_60),
.D(n_83),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_59),
.B(n_83),
.Y(n_154)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_129),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_64),
.B1(n_59),
.B2(n_60),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_125),
.B(n_3),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_2),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_134),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_118),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_97),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_136),
.C(n_145),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_89),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_128),
.A2(n_70),
.B1(n_68),
.B2(n_92),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_142),
.B(n_144),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_108),
.B(n_86),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_100),
.B(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_79),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_87),
.B(n_67),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_91),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_75),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_146),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_88),
.B1(n_67),
.B2(n_74),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_147),
.A2(n_153),
.B1(n_130),
.B2(n_104),
.Y(n_187)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_80),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_149),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_91),
.Y(n_150)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_152),
.A2(n_157),
.B1(n_131),
.B2(n_112),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_151),
.B(n_114),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_125),
.B(n_4),
.Y(n_166)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_113),
.A2(n_72),
.B1(n_59),
.B2(n_73),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_72),
.B1(n_59),
.B2(n_5),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_160),
.A2(n_114),
.B1(n_107),
.B2(n_109),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_161),
.A2(n_134),
.B1(n_132),
.B2(n_160),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_115),
.B1(n_127),
.B2(n_117),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_163),
.A2(n_186),
.B1(n_147),
.B2(n_150),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_141),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_165),
.B(n_180),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_167),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_168),
.A2(n_130),
.B(n_5),
.Y(n_203)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_109),
.A3(n_107),
.B1(n_120),
.B2(n_125),
.Y(n_169)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_120),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_176),
.C(n_179),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_93),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_112),
.C(n_131),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_187),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_137),
.B1(n_158),
.B2(n_148),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_112),
.B1(n_110),
.B2(n_104),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_199),
.B1(n_185),
.B2(n_161),
.Y(n_215)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_194),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_142),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_176),
.C(n_174),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_203),
.B1(n_168),
.B2(n_186),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_139),
.C(n_145),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_9),
.C(n_11),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_155),
.B(n_5),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_198),
.A2(n_206),
.B1(n_185),
.B2(n_178),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_163),
.A2(n_132),
.B1(n_130),
.B2(n_6),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_167),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_202),
.Y(n_220)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_3),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_208),
.B(n_209),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_181),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_3),
.B(n_8),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_184),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_213),
.C(n_222),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_SL g212 ( 
.A1(n_199),
.A2(n_169),
.A3(n_187),
.B1(n_164),
.B2(n_178),
.C1(n_172),
.C2(n_175),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_217),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_192),
.C(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_171),
.Y(n_218)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_171),
.B1(n_174),
.B2(n_10),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_225),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_8),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_8),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_227),
.C(n_201),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_9),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_203),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_190),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_9),
.C(n_10),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_208),
.Y(n_237)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_240),
.C(n_11),
.Y(n_252)
);

INVx13_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_217),
.B1(n_224),
.B2(n_210),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_205),
.C(n_209),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_216),
.A2(n_196),
.B(n_202),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_241),
.B(n_223),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_200),
.B1(n_196),
.B2(n_219),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_242),
.A2(n_243),
.B(n_250),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_200),
.B(n_211),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_252),
.C(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_235),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_222),
.B1(n_227),
.B2(n_14),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_251),
.B(n_232),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_256),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_255),
.C(n_231),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_236),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_258),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_239),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_237),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_244),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_264),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_263),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_256),
.A2(n_246),
.B(n_248),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_231),
.C(n_252),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_265),
.B(n_250),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_266),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_265),
.A2(n_259),
.B1(n_240),
.B2(n_241),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_12),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_271),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_238),
.C(n_15),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_273),
.C(n_270),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_269),
.Y(n_276)
);

AOI321xp33_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_12),
.A3(n_15),
.B1(n_16),
.B2(n_275),
.C(n_249),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_15),
.Y(n_278)
);


endmodule