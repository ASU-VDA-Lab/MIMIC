module fake_jpeg_15798_n_63 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_63);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_63;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_16),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_20),
.B(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_14),
.B(n_1),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_2),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_9),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_8),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

NOR3xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_12),
.C(n_20),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_25),
.B(n_12),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_10),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_22),
.C(n_10),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_18),
.B1(n_11),
.B2(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_37),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_47),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_35),
.C(n_36),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_50),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_49),
.C(n_46),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_44),
.B(n_52),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_42),
.B(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_43),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_53),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_43),
.B2(n_15),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_59),
.B(n_3),
.Y(n_61)
);

A2O1A1O1Ixp25_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_2),
.B(n_3),
.C(n_4),
.D(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);


endmodule