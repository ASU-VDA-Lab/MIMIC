module fake_jpeg_15157_n_380 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_380);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_380;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_46),
.B(n_60),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_23),
.B(n_6),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_52),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_33),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_50),
.A2(n_27),
.B(n_29),
.Y(n_94)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_61),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_6),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_24),
.B1(n_22),
.B2(n_59),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_68),
.A2(n_82),
.B(n_88),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_90),
.Y(n_122)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_81),
.B(n_84),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_43),
.A2(n_24),
.B1(n_22),
.B2(n_33),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_86),
.B(n_102),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_33),
.B1(n_17),
.B2(n_29),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_64),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_11),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_51),
.A2(n_36),
.B1(n_26),
.B2(n_18),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_101),
.B1(n_106),
.B2(n_112),
.Y(n_143)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

BUFx2_ASAP7_75t_SL g118 ( 
.A(n_98),
.Y(n_118)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_26),
.B1(n_36),
.B2(n_18),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_28),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_50),
.A2(n_28),
.B(n_20),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_4),
.B(n_13),
.C(n_2),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_42),
.A2(n_32),
.B1(n_30),
.B2(n_20),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_47),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_7),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_54),
.A2(n_32),
.B1(n_30),
.B2(n_27),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_47),
.A2(n_35),
.B1(n_34),
.B2(n_27),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_4),
.B1(n_10),
.B2(n_13),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_34),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_114),
.B(n_0),
.Y(n_151)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_45),
.A2(n_35),
.B1(n_25),
.B2(n_8),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_52),
.C(n_25),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_131),
.C(n_165),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_121),
.B(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_126),
.B(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_44),
.B1(n_48),
.B2(n_56),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_128),
.A2(n_140),
.B1(n_147),
.B2(n_159),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_130),
.A2(n_139),
.B(n_156),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_83),
.B(n_44),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_41),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_134),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_71),
.A2(n_61),
.B1(n_49),
.B2(n_10),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_135),
.A2(n_142),
.B1(n_104),
.B2(n_96),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_8),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_136),
.B(n_137),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_57),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_7),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_71),
.A2(n_53),
.B1(n_5),
.B2(n_4),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_92),
.A2(n_5),
.B1(n_11),
.B2(n_10),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_95),
.B(n_5),
.CI(n_11),
.CON(n_145),
.SN(n_145)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_149),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_92),
.A2(n_5),
.B1(n_11),
.B2(n_10),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g186 ( 
.A(n_148),
.B(n_79),
.CI(n_96),
.CON(n_186),
.SN(n_186)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_189)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_152),
.B(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_154),
.A2(n_146),
.B1(n_125),
.B2(n_127),
.Y(n_209)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_155),
.B(n_158),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_0),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_68),
.A2(n_0),
.B1(n_1),
.B2(n_112),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_87),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_110),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_0),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_164),
.Y(n_173)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

FAx1_ASAP7_75t_SL g163 ( 
.A(n_82),
.B(n_1),
.CI(n_87),
.CON(n_163),
.SN(n_163)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_79),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_99),
.B(n_100),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_110),
.B(n_103),
.C(n_80),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

MAJx3_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_131),
.C(n_149),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_169),
.B(n_204),
.C(n_205),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_138),
.A2(n_74),
.B1(n_85),
.B2(n_98),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_179),
.A2(n_189),
.B1(n_195),
.B2(n_201),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_184),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_186),
.B(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_121),
.B(n_73),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_188),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_80),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_193),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_126),
.B(n_75),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_130),
.B(n_93),
.Y(n_193)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_157),
.A2(n_143),
.B1(n_119),
.B2(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_131),
.B(n_156),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_211),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_124),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_199),
.Y(n_236)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_157),
.A2(n_163),
.B(n_136),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_140),
.B1(n_163),
.B2(n_122),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_128),
.A2(n_147),
.B1(n_161),
.B2(n_133),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_134),
.B1(n_158),
.B2(n_146),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_156),
.B(n_145),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_145),
.B(n_128),
.C(n_139),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_120),
.B(n_152),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_139),
.B(n_148),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_207),
.B(n_209),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_166),
.A2(n_162),
.B1(n_129),
.B2(n_125),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_189),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_153),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_123),
.B(n_165),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_216),
.A2(n_218),
.B1(n_227),
.B2(n_245),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_155),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_219),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_172),
.A2(n_129),
.B1(n_167),
.B2(n_144),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_144),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_197),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_211),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_230),
.Y(n_274)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_224),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_185),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_197),
.C(n_178),
.Y(n_259)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_226),
.Y(n_269)
);

AO22x1_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_171),
.B1(n_169),
.B2(n_204),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_229),
.B(n_178),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_193),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_168),
.B(n_169),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_232),
.A2(n_249),
.B1(n_221),
.B2(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_202),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_174),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_175),
.B(n_176),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_242),
.B(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_174),
.B(n_169),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_243),
.B(n_246),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_188),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_195),
.A2(n_207),
.B1(n_171),
.B2(n_186),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_210),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_183),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_220),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_170),
.B(n_179),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_200),
.A2(n_205),
.B1(n_181),
.B2(n_190),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_180),
.B1(n_221),
.B2(n_232),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_251),
.B(n_261),
.Y(n_301)
);

CKINVDCx10_ASAP7_75t_R g253 ( 
.A(n_248),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_253),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_183),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_255),
.A2(n_263),
.B(n_265),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_190),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_256),
.B(n_280),
.Y(n_298)
);

INVx13_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_267),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_259),
.B(n_262),
.C(n_272),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_275),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_238),
.B1(n_235),
.B2(n_240),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_264),
.A2(n_245),
.B1(n_233),
.B2(n_213),
.Y(n_287)
);

INVx4_ASAP7_75t_SL g266 ( 
.A(n_226),
.Y(n_266)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_231),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_268),
.B(n_273),
.Y(n_289)
);

NAND3xp33_ASAP7_75t_L g271 ( 
.A(n_236),
.B(n_237),
.C(n_241),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_SL g291 ( 
.A1(n_271),
.A2(n_227),
.B(n_219),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_229),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_215),
.B(n_222),
.C(n_243),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_215),
.B(n_232),
.C(n_217),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_272),
.Y(n_308)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_223),
.Y(n_279)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g280 ( 
.A(n_250),
.B(n_213),
.CI(n_230),
.CON(n_280),
.SN(n_280)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_218),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_233),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_283),
.A2(n_228),
.B1(n_249),
.B2(n_224),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_284),
.A2(n_293),
.B1(n_297),
.B2(n_304),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_287),
.A2(n_310),
.B1(n_297),
.B2(n_280),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_234),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_309),
.Y(n_325)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_262),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_283),
.A2(n_228),
.B(n_212),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_292),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_255),
.A2(n_240),
.B1(n_227),
.B2(n_224),
.Y(n_293)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

OAI22x1_ASAP7_75t_L g297 ( 
.A1(n_255),
.A2(n_212),
.B1(n_214),
.B2(n_251),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_253),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_299),
.B(n_302),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_301),
.B(n_303),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_270),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_252),
.A2(n_276),
.B(n_264),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_263),
.A2(n_281),
.B1(n_258),
.B2(n_274),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_278),
.Y(n_305)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_278),
.Y(n_306)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_269),
.C(n_254),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_280),
.A2(n_281),
.B(n_256),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_312),
.A2(n_319),
.B(n_288),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_289),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_277),
.B1(n_259),
.B2(n_279),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_314),
.A2(n_320),
.B1(n_306),
.B2(n_286),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_316),
.C(n_317),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_300),
.C(n_294),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_254),
.C(n_267),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_266),
.C(n_257),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_324),
.C(n_316),
.Y(n_344)
);

O2A1O1Ixp33_ASAP7_75t_SL g319 ( 
.A1(n_298),
.A2(n_293),
.B(n_284),
.C(n_292),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_305),
.A2(n_304),
.B1(n_303),
.B2(n_309),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_298),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_321),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_290),
.C(n_286),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_295),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_285),
.Y(n_333)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_332),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_333),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_331),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_336),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_285),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_341),
.Y(n_348)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_311),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_343),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_340),
.A2(n_328),
.B1(n_320),
.B2(n_325),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_330),
.B(n_302),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_342),
.A2(n_326),
.B(n_323),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_299),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_344),
.B(n_345),
.C(n_347),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_317),
.C(n_318),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_325),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_322),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_314),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_349),
.B(n_354),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_342),
.A2(n_312),
.B(n_319),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_356),
.C(n_359),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_327),
.C(n_326),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_358),
.B(n_338),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_327),
.C(n_345),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_351),
.B(n_343),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_363),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_361),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_334),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_350),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_365),
.B(n_366),
.C(n_349),
.Y(n_367)
);

OAI322xp33_ASAP7_75t_L g366 ( 
.A1(n_348),
.A2(n_346),
.A3(n_339),
.B1(n_332),
.B2(n_333),
.C1(n_340),
.C2(n_344),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_364),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_362),
.A2(n_351),
.B1(n_355),
.B2(n_358),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_369),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_368),
.B(n_360),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_371),
.B(n_369),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_373),
.B(n_347),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_374),
.A2(n_375),
.B(n_368),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_376),
.B(n_375),
.Y(n_377)
);

AOI322xp5_ASAP7_75t_L g378 ( 
.A1(n_377),
.A2(n_370),
.A3(n_357),
.B1(n_372),
.B2(n_367),
.C1(n_365),
.C2(n_352),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_378),
.A2(n_352),
.B(n_359),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_356),
.Y(n_380)
);


endmodule