module fake_jpeg_26290_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_40),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_21),
.B1(n_30),
.B2(n_20),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_43),
.A2(n_41),
.B1(n_54),
.B2(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_17),
.B(n_32),
.C(n_31),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_40),
.C(n_44),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_23),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_21),
.B1(n_20),
.B2(n_30),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_59),
.A2(n_62),
.B1(n_34),
.B2(n_61),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_39),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_21),
.B1(n_20),
.B2(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_76),
.Y(n_103)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_81),
.B1(n_16),
.B2(n_26),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_41),
.B1(n_34),
.B2(n_42),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_46),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_42),
.C(n_39),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_58),
.C(n_64),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_41),
.B1(n_34),
.B2(n_25),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_89),
.B1(n_63),
.B2(n_61),
.Y(n_96)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_49),
.B1(n_64),
.B2(n_29),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_86),
.A2(n_61),
.B1(n_53),
.B2(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_25),
.B1(n_28),
.B2(n_32),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_91),
.Y(n_106)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_117),
.B1(n_85),
.B2(n_74),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_107),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_101),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_97),
.B1(n_73),
.B2(n_68),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_65),
.B1(n_56),
.B2(n_49),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_46),
.B(n_51),
.C(n_47),
.Y(n_99)
);

A2O1A1O1Ixp25_ASAP7_75t_L g143 ( 
.A1(n_99),
.A2(n_114),
.B(n_29),
.C(n_25),
.D(n_28),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_39),
.C(n_48),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_39),
.C(n_66),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_115),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_51),
.B(n_64),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_0),
.B(n_1),
.Y(n_133)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_78),
.A2(n_80),
.A3(n_81),
.B1(n_17),
.B2(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_80),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_116),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_69),
.Y(n_118)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_110),
.A2(n_27),
.B1(n_69),
.B2(n_72),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

HAxp5_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_27),
.CON(n_121),
.SN(n_121)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_127),
.B(n_133),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_88),
.B1(n_87),
.B2(n_73),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_130),
.B1(n_137),
.B2(n_139),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_140),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_38),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_128),
.A2(n_144),
.B1(n_146),
.B2(n_98),
.Y(n_174)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_141),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_102),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_103),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_38),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_103),
.B(n_99),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_107),
.A2(n_16),
.B1(n_26),
.B2(n_31),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_28),
.B1(n_25),
.B2(n_18),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_106),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_113),
.Y(n_167)
);

NOR2x1p5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_117),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_28),
.B1(n_18),
.B2(n_19),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_150),
.C(n_154),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_94),
.C(n_99),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_152),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_145),
.B(n_122),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_100),
.C(n_104),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_163),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_96),
.B1(n_100),
.B2(n_92),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_168),
.B1(n_119),
.B2(n_129),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_1),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_128),
.A2(n_116),
.B1(n_105),
.B2(n_118),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_174),
.B1(n_176),
.B2(n_19),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_105),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_113),
.B(n_98),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_192)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_66),
.C(n_95),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_169),
.C(n_170),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_171),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_124),
.A2(n_98),
.B1(n_19),
.B2(n_18),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_132),
.B(n_11),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_38),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_22),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_125),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_126),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_22),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_67),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_143),
.B1(n_120),
.B2(n_140),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_127),
.A3(n_125),
.B1(n_133),
.B2(n_139),
.C1(n_123),
.C2(n_135),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_179),
.A2(n_186),
.B(n_192),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_193),
.Y(n_206)
);

AO22x1_ASAP7_75t_SL g184 ( 
.A1(n_161),
.A2(n_127),
.B1(n_135),
.B2(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_141),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_147),
.B1(n_157),
.B2(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_22),
.Y(n_191)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_19),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_202),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_195),
.A2(n_200),
.B1(n_13),
.B2(n_12),
.Y(n_217)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_197),
.Y(n_215)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_67),
.B1(n_33),
.B2(n_15),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_198),
.A2(n_201),
.B1(n_2),
.B2(n_5),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_156),
.A2(n_0),
.B(n_1),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_199),
.A2(n_156),
.B(n_3),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_0),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_147),
.B(n_14),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_148),
.C(n_150),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_209),
.C(n_211),
.Y(n_228)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_207),
.A2(n_199),
.B(n_201),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_212),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_152),
.C(n_151),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_166),
.C(n_154),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_157),
.B1(n_171),
.B2(n_169),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_191),
.B(n_13),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_217),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_13),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_202),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_11),
.C(n_3),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_221),
.C(n_192),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_2),
.C(n_3),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_226),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_188),
.B1(n_194),
.B2(n_197),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_184),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_208),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_231),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_187),
.B(n_189),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_187),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_189),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_236),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_246),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_185),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_185),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_243),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_184),
.C(n_200),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_240),
.C(n_242),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_212),
.C(n_216),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_184),
.C(n_193),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_221),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_219),
.C(n_206),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_201),
.B(n_190),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_251),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_234),
.A2(n_224),
.B(n_207),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_259),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_255),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_177),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_235),
.A2(n_182),
.B(n_196),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_259),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_210),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_261),
.B(n_243),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_205),
.A3(n_179),
.B1(n_198),
.B2(n_210),
.C1(n_226),
.C2(n_181),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_262),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_238),
.A2(n_224),
.B1(n_218),
.B2(n_182),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_263),
.A2(n_218),
.B1(n_245),
.B2(n_239),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_275),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_236),
.C(n_237),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_228),
.C(n_233),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_177),
.Y(n_269)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_272),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_250),
.A2(n_240),
.B1(n_228),
.B2(n_7),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_5),
.C(n_6),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_6),
.Y(n_285)
);

AOI21x1_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_251),
.B(n_252),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_9),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_274),
.A2(n_253),
.B1(n_263),
.B2(n_254),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_265),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_255),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_283),
.B(n_8),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_257),
.B1(n_258),
.B2(n_8),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_258),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_9),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_288),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_267),
.C(n_278),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_292),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_6),
.B(n_7),
.Y(n_291)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_8),
.C(n_9),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_293),
.B(n_294),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_280),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_295),
.A2(n_296),
.B(n_283),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_302),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_279),
.B(n_10),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_304),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_293),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_303),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_305),
.B(n_301),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_298),
.Y(n_309)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_10),
.CI(n_306),
.CON(n_310),
.SN(n_310)
);


endmodule