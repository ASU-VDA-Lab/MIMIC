module fake_aes_2230_n_41 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_41);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_10), .B(n_13), .Y(n_17) );
OR2x2_ASAP7_75t_L g18 ( .A(n_12), .B(n_14), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_4), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_11), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_0), .Y(n_21) );
INVx3_ASAP7_75t_L g22 ( .A(n_5), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_0), .Y(n_23) );
BUFx3_ASAP7_75t_L g24 ( .A(n_16), .Y(n_24) );
NOR3xp33_ASAP7_75t_SL g25 ( .A(n_15), .B(n_1), .C(n_2), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_19), .B1(n_21), .B2(n_22), .Y(n_26) );
OAI22xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_19), .B1(n_22), .B2(n_20), .Y(n_27) );
BUFx2_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_28), .B(n_26), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
OAI21xp33_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_24), .B(n_23), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_29), .B(n_24), .Y(n_32) );
INVxp67_ASAP7_75t_L g33 ( .A(n_32), .Y(n_33) );
OAI221xp5_ASAP7_75t_L g34 ( .A1(n_31), .A2(n_30), .B1(n_29), .B2(n_16), .C(n_18), .Y(n_34) );
AOI221xp5_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_20), .B1(n_17), .B2(n_18), .C(n_5), .Y(n_35) );
NAND2xp33_ASAP7_75t_R g36 ( .A(n_35), .B(n_2), .Y(n_36) );
AOI22xp33_ASAP7_75t_SL g37 ( .A1(n_34), .A2(n_17), .B1(n_4), .B2(n_6), .Y(n_37) );
OR2x2_ASAP7_75t_L g38 ( .A(n_33), .B(n_3), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_38), .Y(n_39) );
HB1xp67_ASAP7_75t_L g40 ( .A(n_36), .Y(n_40) );
AOI322xp5_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_3), .A3(n_6), .B1(n_7), .B2(n_8), .C1(n_37), .C2(n_39), .Y(n_41) );
endmodule