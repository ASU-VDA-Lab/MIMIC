module real_jpeg_12330_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g104 ( 
.A(n_0),
.Y(n_104)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_3),
.A2(n_38),
.B1(n_64),
.B2(n_66),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_38),
.B1(n_47),
.B2(n_48),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_4),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_122),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_122),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_4),
.A2(n_64),
.B1(n_66),
.B2(n_122),
.Y(n_249)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_54),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_6),
.A2(n_54),
.B1(n_64),
.B2(n_66),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_7),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_151),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_151),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_7),
.A2(n_64),
.B1(n_66),
.B2(n_151),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_10),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_120),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_120),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_10),
.A2(n_64),
.B1(n_66),
.B2(n_120),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_11),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_11),
.B(n_36),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_11),
.B(n_62),
.C(n_64),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_144),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_11),
.A2(n_102),
.B1(n_109),
.B2(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_11),
.B(n_43),
.Y(n_266)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_13),
.A2(n_50),
.B1(n_64),
.B2(n_66),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_50),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_14),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_14),
.A2(n_24),
.B1(n_64),
.B2(n_66),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_14),
.A2(n_24),
.B1(n_34),
.B2(n_35),
.Y(n_161)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_94),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_82),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_82),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_74),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_20),
.A2(n_21),
.B1(n_70),
.B2(n_71),
.Y(n_320)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_22),
.B(n_41),
.C(n_57),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_36),
.B2(n_37),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_23),
.A2(n_36),
.B(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

HAxp5_ASAP7_75t_SL g143 ( 
.A(n_25),
.B(n_144),
.CON(n_143),
.SN(n_143)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_25),
.B(n_32),
.C(n_34),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_28),
.A2(n_37),
.B(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_28),
.A2(n_36),
.B1(n_143),
.B2(n_150),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_28),
.A2(n_86),
.B(n_164),
.Y(n_301)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_29),
.B(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_29),
.A2(n_33),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_29),
.A2(n_33),
.B1(n_119),
.B2(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_29),
.A2(n_121),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_31),
.A2(n_35),
.B(n_143),
.C(n_145),
.Y(n_142)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_33),
.B(n_73),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_56)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g214 ( 
.A(n_35),
.B(n_144),
.CON(n_214),
.SN(n_214)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_35),
.B(n_45),
.C(n_48),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_36),
.B(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_57),
.B2(n_69),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_51),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_42),
.A2(n_77),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_49),
.B(n_55),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_43),
.A2(n_55),
.B1(n_191),
.B2(n_214),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_43),
.A2(n_55),
.B1(n_79),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_53),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_44),
.A2(n_51),
.B(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_44),
.A2(n_77),
.B1(n_147),
.B2(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_44),
.A2(n_77),
.B1(n_182),
.B2(n_190),
.Y(n_189)
);

OA22x2_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_46),
.A2(n_47),
.B(n_214),
.C(n_215),
.Y(n_213)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_48),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_47),
.B(n_240),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_49),
.A2(n_55),
.B(n_81),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_71),
.C(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_57),
.A2(n_69),
.B1(n_76),
.B2(n_316),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_67),
.B(n_68),
.Y(n_57)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_58),
.A2(n_67),
.B1(n_112),
.B2(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_58),
.A2(n_134),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_58),
.A2(n_68),
.B(n_171),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_58),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_58),
.A2(n_67),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_58),
.A2(n_67),
.B1(n_219),
.B2(n_244),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_SL g62 ( 
.A(n_60),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_63),
.B(n_114),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_63),
.A2(n_115),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_63),
.B(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_64),
.Y(n_66)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_66),
.B(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_67),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_67),
.B(n_144),
.Y(n_257)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_68),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_70),
.A2(n_71),
.B1(n_315),
.B2(n_317),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_74),
.A2(n_75),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_76),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_80),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_310),
.B(n_327),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_290),
.B(n_309),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_174),
.B(n_289),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_152),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_98),
.B(n_152),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_125),
.C(n_135),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_99),
.B(n_125),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_116),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_100),
.B(n_117),
.C(n_124),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_111),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_101),
.B(n_111),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_105),
.B(n_107),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_102),
.A2(n_109),
.B(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_102),
.A2(n_109),
.B1(n_247),
.B2(n_255),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_102),
.A2(n_130),
.B(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_103),
.A2(n_108),
.B(n_131),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_103),
.A2(n_104),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_131),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_109),
.A2(n_128),
.B(n_141),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_109),
.B(n_144),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_113),
.B(n_229),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_123),
.B2(n_124),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_132),
.B2(n_133),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_133),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_135),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_146),
.C(n_148),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_136),
.A2(n_137),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_148),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_173),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_165),
.B2(n_166),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_154),
.B(n_166),
.C(n_173),
.Y(n_308)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_156),
.B(n_160),
.C(n_162),
.Y(n_293)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_161),
.Y(n_306)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_172),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_167),
.A2(n_168),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_168),
.B(n_170),
.Y(n_298)
);

AOI21xp33_ASAP7_75t_L g318 ( 
.A1(n_168),
.A2(n_298),
.B(n_301),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_170),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_202),
.B(n_284),
.C(n_288),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_195),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_195),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_185),
.C(n_188),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_177),
.B(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_180),
.C(n_184),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_188),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_189),
.B(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_196),
.B(n_200),
.C(n_201),
.Y(n_285)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_278),
.B(n_283),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_233),
.B(n_277),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_221),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_207),
.B(n_221),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_216),
.C(n_217),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_208),
.A2(n_209),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_210),
.B(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_216),
.B(n_217),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_220),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_222),
.B(n_227),
.C(n_231),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_231),
.B2(n_232),
.Y(n_225)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_226),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_227),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_271),
.B(n_276),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_261),
.B(n_270),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_250),
.B(n_260),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_245),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_245),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_241),
.Y(n_262)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_256),
.B(n_259),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_258),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_263),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_269),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_268),
.C(n_269),
.Y(n_275)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_275),
.Y(n_276)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_282),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_286),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_308),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_308),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_296),
.C(n_303),
.Y(n_323)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_302),
.B2(n_303),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_305),
.B(n_307),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_313),
.C(n_318),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_307),
.A2(n_313),
.B1(n_314),
.B2(n_326),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_307),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_322),
.Y(n_310)
);

AOI21xp33_ASAP7_75t_L g327 ( 
.A1(n_311),
.A2(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_319),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_319),
.Y(n_329)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);


endmodule