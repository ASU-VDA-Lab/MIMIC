module fake_ibex_806_n_2790 (n_151, n_85, n_507, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_8, n_224, n_183, n_508, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_22, n_136, n_261, n_459, n_30, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_483, n_141, n_487, n_222, n_186, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_484, n_480, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_199, n_495, n_410, n_308, n_463, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_479, n_225, n_360, n_272, n_23, n_468, n_223, n_381, n_382, n_502, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_313, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_425, n_2790);

input n_151;
input n_85;
input n_507;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_508;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_22;
input n_136;
input n_261;
input n_459;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_141;
input n_487;
input n_222;
input n_186;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_199;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_479;
input n_225;
input n_360;
input n_272;
input n_23;
input n_468;
input n_223;
input n_381;
input n_382;
input n_502;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2790;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2498;
wire n_1802;
wire n_2235;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1954;
wire n_2183;
wire n_1859;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_708;
wire n_1096;
wire n_2391;
wire n_2151;
wire n_1391;
wire n_667;
wire n_884;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2724;
wire n_2475;
wire n_853;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_2311;
wire n_527;
wire n_893;
wire n_1654;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_523;
wire n_787;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2347;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_554;
wire n_553;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2112;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_971;
wire n_1326;
wire n_702;
wire n_1350;
wire n_906;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_2723;
wire n_1616;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_2224;
wire n_1862;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_2779;
wire n_521;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_660;
wire n_2590;
wire n_524;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_607;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_2095;
wire n_555;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2352;
wire n_2212;
wire n_2716;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_2654;
wire n_2463;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_528;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_916;
wire n_2298;
wire n_2771;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_545;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_961;
wire n_991;
wire n_634;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_2617;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2639;
wire n_2330;
wire n_636;
wire n_1259;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_2688;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2149;
wire n_2268;
wire n_2320;
wire n_2237;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_2758;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2447;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_520;
wire n_775;
wire n_512;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_2608;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_2669;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_2518;
wire n_2784;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1635;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_2734;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_2634;
wire n_1092;
wire n_1808;
wire n_560;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_924;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_2092;
wire n_566;
wire n_581;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_548;
wire n_1158;
wire n_1974;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2704;
wire n_1915;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_2754;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_2738;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

INVx1_ASAP7_75t_L g511 ( 
.A(n_41),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_247),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_296),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_185),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_426),
.Y(n_515)
);

CKINVDCx14_ASAP7_75t_R g516 ( 
.A(n_425),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_481),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_128),
.B(n_279),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_412),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_102),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_203),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_218),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_121),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_371),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_167),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_199),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_102),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_254),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_498),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_114),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_197),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_258),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_159),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_192),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_485),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_207),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_200),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_187),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_143),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_360),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_162),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_475),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_302),
.Y(n_543)
);

INVxp33_ASAP7_75t_L g544 ( 
.A(n_504),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_321),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_208),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_487),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_147),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_215),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_416),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_175),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_328),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_356),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_247),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_491),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_506),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_333),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_261),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_198),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_440),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_472),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_6),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_158),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_488),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_16),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_128),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_444),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_71),
.B(n_397),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_149),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_43),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_346),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_372),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_204),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_36),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_133),
.Y(n_575)
);

NOR2xp67_ASAP7_75t_L g576 ( 
.A(n_459),
.B(n_283),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_375),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_240),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_348),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_95),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_486),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_336),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_510),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_461),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_332),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_300),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_392),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_225),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_273),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g590 ( 
.A(n_413),
.B(n_451),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_409),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_273),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_25),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_434),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_211),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_331),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_239),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_232),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_44),
.B(n_266),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_83),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_44),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_382),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_386),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_123),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_294),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_147),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_238),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_275),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_352),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_445),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_92),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_285),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_32),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_505),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_183),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_473),
.Y(n_616)
);

CKINVDCx16_ASAP7_75t_R g617 ( 
.A(n_183),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_300),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_405),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_420),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_193),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_45),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_344),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_245),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_59),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_215),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_115),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_463),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_297),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_277),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_446),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_452),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_423),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_367),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_464),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_217),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_507),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_210),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_248),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_332),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_254),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_231),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_84),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_32),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_366),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_427),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_419),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_467),
.Y(n_648)
);

BUFx8_ASAP7_75t_SL g649 ( 
.A(n_443),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_442),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_439),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_368),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_410),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_347),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_10),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_492),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_140),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_161),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_278),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_173),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_106),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_122),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_14),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_469),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_249),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_221),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_276),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_272),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_292),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_200),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_466),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_489),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_500),
.B(n_50),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_81),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_441),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_285),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_116),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_373),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_211),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_428),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_138),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_220),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_453),
.Y(n_683)
);

INVxp33_ASAP7_75t_L g684 ( 
.A(n_72),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_308),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_493),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_490),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_338),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_421),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_497),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_479),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_435),
.Y(n_692)
);

CKINVDCx16_ASAP7_75t_R g693 ( 
.A(n_430),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_84),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_195),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_31),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_240),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_454),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_223),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_207),
.Y(n_700)
);

BUFx10_ASAP7_75t_L g701 ( 
.A(n_93),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_389),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_499),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_27),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_187),
.Y(n_705)
);

CKINVDCx16_ASAP7_75t_R g706 ( 
.A(n_50),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_137),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_9),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_28),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_106),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_29),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_380),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_205),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_449),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_438),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_74),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_151),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_252),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_311),
.Y(n_719)
);

NOR2xp67_ASAP7_75t_L g720 ( 
.A(n_431),
.B(n_348),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_414),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_322),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_114),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_457),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_251),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_494),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_227),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_437),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_227),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_337),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_212),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_407),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_56),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_460),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_318),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_468),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_429),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_132),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_161),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_317),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_175),
.Y(n_741)
);

XOR2xp5_ASAP7_75t_R g742 ( 
.A(n_432),
.B(n_3),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_404),
.Y(n_743)
);

CKINVDCx11_ASAP7_75t_R g744 ( 
.A(n_137),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_159),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_150),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_64),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_509),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_145),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_250),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_402),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_323),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_262),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_245),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_8),
.Y(n_755)
);

BUFx10_ASAP7_75t_L g756 ( 
.A(n_80),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_45),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_62),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_139),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_501),
.B(n_334),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_99),
.Y(n_761)
);

CKINVDCx16_ASAP7_75t_R g762 ( 
.A(n_508),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_258),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_28),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_174),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_373),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_36),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_408),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_251),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_318),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_495),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_478),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_75),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_378),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_474),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_502),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_471),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_261),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_417),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_448),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_143),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_304),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_411),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_401),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_477),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_244),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_321),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_436),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_118),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_2),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_104),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_39),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_208),
.Y(n_793)
);

BUFx10_ASAP7_75t_L g794 ( 
.A(n_115),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_296),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_196),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_217),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_424),
.Y(n_798)
);

CKINVDCx14_ASAP7_75t_R g799 ( 
.A(n_480),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_398),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_350),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_95),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_305),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_69),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_319),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_433),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_344),
.Y(n_807)
);

CKINVDCx16_ASAP7_75t_R g808 ( 
.A(n_34),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_269),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_101),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_77),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_470),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_222),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_103),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_312),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_496),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_503),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_476),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_160),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_248),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_23),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_23),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_335),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_133),
.Y(n_824)
);

NOR2xp67_ASAP7_75t_L g825 ( 
.A(n_34),
.B(n_353),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_418),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_219),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_447),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_309),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_456),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_337),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_450),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_326),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_91),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_190),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_105),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_130),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_129),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_268),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_24),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_10),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_660),
.Y(n_842)
);

OAI22x1_ASAP7_75t_SL g843 ( 
.A1(n_521),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_535),
.Y(n_844)
);

INVxp33_ASAP7_75t_L g845 ( 
.A(n_684),
.Y(n_845)
);

BUFx12f_ASAP7_75t_L g846 ( 
.A(n_698),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_678),
.B(n_0),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_684),
.B(n_1),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_660),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_515),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_744),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_562),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_581),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_584),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_649),
.Y(n_855)
);

INVx5_ASAP7_75t_L g856 ( 
.A(n_535),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_562),
.Y(n_857)
);

INVx5_ASAP7_75t_L g858 ( 
.A(n_535),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_755),
.B(n_4),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_527),
.B(n_4),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_689),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_522),
.B(n_5),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_689),
.Y(n_863)
);

OAI21x1_ASAP7_75t_L g864 ( 
.A1(n_691),
.A2(n_391),
.B(n_390),
.Y(n_864)
);

BUFx12f_ASAP7_75t_L g865 ( 
.A(n_744),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_512),
.B(n_6),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_691),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_545),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_528),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_557),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_562),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_649),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_535),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_665),
.B(n_7),
.Y(n_874)
);

OA21x2_ASAP7_75t_L g875 ( 
.A1(n_561),
.A2(n_583),
.B(n_564),
.Y(n_875)
);

INVx4_ASAP7_75t_L g876 ( 
.A(n_542),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_668),
.B(n_11),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_567),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_567),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_567),
.Y(n_880)
);

BUFx12f_ASAP7_75t_L g881 ( 
.A(n_667),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_589),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_607),
.B(n_12),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_589),
.B(n_13),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_675),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_682),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_682),
.B(n_14),
.Y(n_887)
);

OA21x2_ASAP7_75t_L g888 ( 
.A1(n_619),
.A2(n_394),
.B(n_393),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_667),
.Y(n_889)
);

INVx4_ASAP7_75t_L g890 ( 
.A(n_547),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_675),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_694),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_667),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_739),
.B(n_15),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_617),
.B(n_15),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_670),
.Y(n_896)
);

OAI22x1_ASAP7_75t_SL g897 ( 
.A1(n_521),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_897)
);

OAI21x1_ASAP7_75t_L g898 ( 
.A1(n_620),
.A2(n_396),
.B(n_395),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_818),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_701),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_739),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_818),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_670),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_718),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_610),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_830),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_718),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_830),
.B(n_18),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_515),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_544),
.B(n_19),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_774),
.B(n_19),
.Y(n_911)
);

OAI22x1_ASAP7_75t_SL g912 ( 
.A1(n_533),
.A2(n_541),
.B1(n_559),
.B2(n_549),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_540),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_693),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_914)
);

CKINVDCx16_ASAP7_75t_R g915 ( 
.A(n_706),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_701),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_519),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_685),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_610),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_513),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_SL g921 ( 
.A(n_762),
.B(n_399),
.Y(n_921)
);

AND2x2_ASAP7_75t_SL g922 ( 
.A(n_568),
.B(n_400),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_540),
.B(n_20),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_513),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_550),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_631),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_513),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_513),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_578),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_574),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_574),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_578),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_808),
.B(n_21),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_685),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_934)
);

AND2x6_ASAP7_75t_L g935 ( 
.A(n_650),
.B(n_403),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_656),
.Y(n_936)
);

INVx5_ASAP7_75t_L g937 ( 
.A(n_578),
.Y(n_937)
);

BUFx8_ASAP7_75t_SL g938 ( 
.A(n_533),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_578),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_664),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_845),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_845),
.B(n_544),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_844),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_844),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_844),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_876),
.B(n_835),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_844),
.Y(n_947)
);

NOR2x1p5_ASAP7_75t_L g948 ( 
.A(n_881),
.B(n_742),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_873),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_911),
.B(n_671),
.Y(n_950)
);

BUFx6f_ASAP7_75t_SL g951 ( 
.A(n_922),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_911),
.B(n_672),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_860),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_873),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_873),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_935),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_873),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_853),
.B(n_785),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_869),
.B(n_516),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_884),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_884),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_887),
.Y(n_962)
);

BUFx4f_ASAP7_75t_L g963 ( 
.A(n_881),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_878),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_869),
.B(n_837),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_878),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_878),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_878),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_876),
.B(n_828),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_879),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_887),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_879),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_935),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_879),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_918),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_879),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_887),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_L g978 ( 
.A(n_935),
.B(n_555),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_880),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_911),
.B(n_683),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_892),
.B(n_799),
.Y(n_981)
);

AND3x2_ASAP7_75t_L g982 ( 
.A(n_921),
.B(n_793),
.C(n_531),
.Y(n_982)
);

INVx5_ASAP7_75t_L g983 ( 
.A(n_935),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_894),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_880),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_894),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_935),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_926),
.B(n_687),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_923),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_926),
.B(n_703),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_923),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_936),
.B(n_714),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_L g993 ( 
.A(n_885),
.B(n_891),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_896),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_896),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_870),
.Y(n_996)
);

BUFx10_ASAP7_75t_L g997 ( 
.A(n_855),
.Y(n_997)
);

INVx8_ASAP7_75t_L g998 ( 
.A(n_851),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_886),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_918),
.Y(n_1000)
);

XNOR2x2_ASAP7_75t_L g1001 ( 
.A(n_934),
.B(n_518),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_892),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_905),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_890),
.B(n_715),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_852),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_901),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_885),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_891),
.Y(n_1008)
);

INVxp33_ASAP7_75t_L g1009 ( 
.A(n_848),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_905),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_852),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_925),
.B(n_721),
.Y(n_1012)
);

BUFx10_ASAP7_75t_L g1013 ( 
.A(n_855),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_899),
.Y(n_1014)
);

OAI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_914),
.A2(n_882),
.B1(n_868),
.B2(n_915),
.Y(n_1015)
);

BUFx10_ASAP7_75t_L g1016 ( 
.A(n_872),
.Y(n_1016)
);

AOI21x1_ASAP7_75t_L g1017 ( 
.A1(n_864),
.A2(n_732),
.B(n_724),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_936),
.B(n_734),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_857),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_857),
.B(n_889),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_919),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_889),
.B(n_582),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_899),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_902),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_940),
.B(n_736),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_902),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_862),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_919),
.Y(n_1028)
);

NAND2xp33_ASAP7_75t_L g1029 ( 
.A(n_908),
.B(n_529),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_864),
.A2(n_751),
.B(n_743),
.Y(n_1030)
);

AO21x2_ASAP7_75t_L g1031 ( 
.A1(n_898),
.A2(n_760),
.B(n_768),
.Y(n_1031)
);

NOR2x1p5_ASAP7_75t_L g1032 ( 
.A(n_851),
.B(n_836),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_893),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_906),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_893),
.B(n_837),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_920),
.Y(n_1036)
);

INVx5_ASAP7_75t_L g1037 ( 
.A(n_856),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_940),
.B(n_838),
.Y(n_1038)
);

OR2x6_ASAP7_75t_L g1039 ( 
.A(n_865),
.B(n_825),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_920),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_920),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_842),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_909),
.B(n_772),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_849),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_924),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_871),
.B(n_900),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_903),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_916),
.B(n_838),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_924),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_904),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_924),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_927),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_907),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_930),
.B(n_839),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_927),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_930),
.B(n_775),
.Y(n_1056)
);

AO21x2_ASAP7_75t_L g1057 ( 
.A1(n_898),
.A2(n_874),
.B(n_866),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_927),
.Y(n_1058)
);

NAND2xp33_ASAP7_75t_SL g1059 ( 
.A(n_872),
.B(n_517),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_850),
.B(n_776),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_865),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_846),
.B(n_777),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_854),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_909),
.B(n_779),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_928),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_928),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_883),
.Y(n_1067)
);

BUFx10_ASAP7_75t_L g1068 ( 
.A(n_922),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_846),
.B(n_701),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_913),
.B(n_783),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_854),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_928),
.Y(n_1072)
);

AO21x2_ASAP7_75t_L g1073 ( 
.A1(n_877),
.A2(n_800),
.B(n_788),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_929),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_861),
.Y(n_1075)
);

AND3x2_ASAP7_75t_L g1076 ( 
.A(n_895),
.B(n_910),
.C(n_630),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_917),
.B(n_839),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_929),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_932),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_861),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_863),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_863),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_875),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_932),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_932),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_867),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_931),
.B(n_840),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_867),
.B(n_812),
.Y(n_1088)
);

BUFx10_ASAP7_75t_L g1089 ( 
.A(n_939),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_875),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_847),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_937),
.B(n_841),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_L g1093 ( 
.A(n_859),
.B(n_933),
.C(n_697),
.Y(n_1093)
);

BUFx4f_ASAP7_75t_L g1094 ( 
.A(n_888),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_937),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1022),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_1002),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_942),
.B(n_529),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_1046),
.B(n_556),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1046),
.B(n_556),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_941),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_941),
.B(n_711),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_956),
.B(n_560),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1022),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_1000),
.Y(n_1105)
);

OR2x6_ASAP7_75t_L g1106 ( 
.A(n_998),
.B(n_948),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1063),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_975),
.A2(n_587),
.B1(n_591),
.B2(n_517),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_965),
.B(n_532),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1073),
.B(n_817),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_953),
.B(n_832),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_973),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1019),
.B(n_647),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_998),
.B(n_843),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_1054),
.B(n_606),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_959),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1019),
.B(n_680),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_1005),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_983),
.B(n_1091),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_973),
.B(n_594),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_987),
.B(n_628),
.Y(n_1121)
);

NOR2xp67_ASAP7_75t_L g1122 ( 
.A(n_1061),
.B(n_673),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1063),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_994),
.B(n_587),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_981),
.Y(n_1125)
);

INVxp67_ASAP7_75t_L g1126 ( 
.A(n_1038),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_960),
.B(n_633),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_996),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_962),
.B(n_635),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_971),
.B(n_637),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_987),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1033),
.B(n_546),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_995),
.A2(n_730),
.B(n_599),
.C(n_514),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1033),
.B(n_646),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_963),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_977),
.B(n_648),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1007),
.Y(n_1137)
);

INVx8_ASAP7_75t_L g1138 ( 
.A(n_998),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1008),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1005),
.B(n_651),
.Y(n_1140)
);

NOR2xp67_ASAP7_75t_L g1141 ( 
.A(n_1093),
.B(n_856),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_946),
.B(n_653),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1011),
.B(n_1035),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_999),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1006),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1004),
.B(n_690),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1004),
.B(n_692),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1020),
.B(n_1048),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1012),
.B(n_726),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1009),
.B(n_711),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_963),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_984),
.B(n_728),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1090),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_986),
.B(n_748),
.Y(n_1154)
);

INVxp67_ASAP7_75t_L g1155 ( 
.A(n_1069),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1009),
.B(n_711),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_1059),
.Y(n_1157)
);

OR2x6_ASAP7_75t_L g1158 ( 
.A(n_1032),
.B(n_897),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1012),
.B(n_798),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_L g1160 ( 
.A(n_1027),
.B(n_525),
.C(n_520),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_969),
.B(n_958),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1067),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_961),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_961),
.B(n_816),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_958),
.B(n_826),
.Y(n_1165)
);

INVx8_ASAP7_75t_L g1166 ( 
.A(n_1039),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1087),
.B(n_695),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1014),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1023),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1077),
.B(n_536),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1024),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1026),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_1059),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1034),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_989),
.B(n_537),
.Y(n_1175)
);

XOR2xp5_ASAP7_75t_L g1176 ( 
.A(n_1001),
.B(n_912),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_SL g1177 ( 
.A(n_997),
.Y(n_1177)
);

NAND2xp33_ASAP7_75t_SL g1178 ( 
.A(n_951),
.B(n_591),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_991),
.B(n_548),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_950),
.B(n_551),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_950),
.B(n_952),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_993),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1042),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_952),
.B(n_554),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_980),
.B(n_888),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1071),
.Y(n_1186)
);

OR2x6_ASAP7_75t_L g1187 ( 
.A(n_1039),
.B(n_582),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_982),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1075),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1062),
.B(n_570),
.Y(n_1190)
);

AOI221xp5_ASAP7_75t_L g1191 ( 
.A1(n_1015),
.A2(n_524),
.B1(n_526),
.B2(n_523),
.C(n_511),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1068),
.B(n_592),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_951),
.A2(n_616),
.B1(n_632),
.B2(n_614),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_997),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1044),
.B(n_627),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1047),
.B(n_627),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1050),
.B(n_674),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1092),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1053),
.B(n_674),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1029),
.B(n_571),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1080),
.Y(n_1201)
);

NOR2xp67_ASAP7_75t_L g1202 ( 
.A(n_1056),
.B(n_858),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1081),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1029),
.B(n_1060),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1013),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1076),
.B(n_572),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1013),
.B(n_1016),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1083),
.B(n_704),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1082),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1086),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1070),
.A2(n_534),
.B(n_538),
.C(n_530),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1025),
.B(n_988),
.Y(n_1212)
);

AND2x2_ASAP7_75t_SL g1213 ( 
.A(n_978),
.B(n_938),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1015),
.A2(n_616),
.B1(n_632),
.B2(n_614),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1016),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_982),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1039),
.B(n_756),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1076),
.B(n_756),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_988),
.B(n_704),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_1070),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_990),
.B(n_729),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_990),
.B(n_729),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_992),
.B(n_741),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_992),
.B(n_741),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1018),
.B(n_1043),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1089),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1089),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1043),
.B(n_681),
.Y(n_1228)
);

INVxp67_ASAP7_75t_L g1229 ( 
.A(n_1088),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_1064),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1088),
.B(n_822),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1057),
.B(n_789),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1095),
.B(n_773),
.Y(n_1233)
);

NAND2x1p5_ASAP7_75t_L g1234 ( 
.A(n_1037),
.B(n_539),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1031),
.B(n_756),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1037),
.A2(n_543),
.B1(n_553),
.B2(n_552),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1037),
.A2(n_737),
.B1(n_771),
.B2(n_686),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1037),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1017),
.B(n_795),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1030),
.B(n_831),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_943),
.B(n_831),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_945),
.B(n_579),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_943),
.B(n_833),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_944),
.B(n_558),
.Y(n_1244)
);

XOR2xp5_ASAP7_75t_L g1245 ( 
.A(n_1036),
.B(n_686),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1040),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_947),
.B(n_563),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_947),
.B(n_565),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_945),
.B(n_576),
.Y(n_1249)
);

INVx4_ASAP7_75t_L g1250 ( 
.A(n_945),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_954),
.B(n_566),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_949),
.B(n_720),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_949),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1041),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_954),
.B(n_575),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_955),
.B(n_580),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1045),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1045),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_955),
.B(n_586),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_957),
.B(n_593),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_949),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1049),
.B(n_794),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1051),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_957),
.B(n_596),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_949),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_964),
.B(n_598),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_964),
.B(n_600),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1051),
.B(n_794),
.Y(n_1268)
);

INVx8_ASAP7_75t_L g1269 ( 
.A(n_972),
.Y(n_1269)
);

AOI221xp5_ASAP7_75t_L g1270 ( 
.A1(n_966),
.A2(n_603),
.B1(n_611),
.B2(n_609),
.C(n_602),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_966),
.B(n_612),
.Y(n_1271)
);

NAND2xp33_ASAP7_75t_L g1272 ( 
.A(n_972),
.B(n_737),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1052),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_967),
.B(n_613),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_972),
.B(n_595),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_SL g1276 ( 
.A(n_972),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1055),
.A2(n_780),
.B1(n_784),
.B2(n_771),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_L g1278 ( 
.A(n_1058),
.B(n_608),
.C(n_605),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_968),
.B(n_618),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1058),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1021),
.B(n_615),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1065),
.B(n_794),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1065),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1066),
.A2(n_784),
.B1(n_806),
.B2(n_780),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1066),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1072),
.Y(n_1286)
);

AND2x2_ASAP7_75t_SL g1287 ( 
.A(n_1074),
.B(n_938),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_SL g1288 ( 
.A(n_1021),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1078),
.B(n_624),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1079),
.B(n_626),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1079),
.A2(n_806),
.B1(n_636),
.B2(n_638),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_970),
.B(n_623),
.Y(n_1292)
);

INVx4_ASAP7_75t_L g1293 ( 
.A(n_974),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_974),
.B(n_625),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_976),
.B(n_629),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_979),
.B(n_634),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_979),
.B(n_641),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1084),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1138),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1097),
.Y(n_1300)
);

NAND2xp33_ASAP7_75t_L g1301 ( 
.A(n_1112),
.B(n_639),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1185),
.A2(n_590),
.B(n_985),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1138),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1105),
.B(n_541),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1118),
.B(n_642),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1220),
.B(n_643),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1161),
.A2(n_559),
.B1(n_569),
.B2(n_549),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1155),
.B(n_569),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1101),
.B(n_573),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1116),
.B(n_573),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1118),
.B(n_652),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1148),
.B(n_644),
.Y(n_1312)
);

BUFx4f_ASAP7_75t_L g1313 ( 
.A(n_1138),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1194),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1143),
.B(n_658),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1109),
.B(n_645),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1284),
.B(n_577),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1126),
.B(n_1098),
.Y(n_1318)
);

AOI21xp33_ASAP7_75t_L g1319 ( 
.A1(n_1188),
.A2(n_655),
.B(n_654),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1108),
.B(n_577),
.Y(n_1320)
);

NOR2xp67_ASAP7_75t_SL g1321 ( 
.A(n_1205),
.B(n_657),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1181),
.B(n_659),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1215),
.Y(n_1323)
);

NOR3xp33_ASAP7_75t_L g1324 ( 
.A(n_1191),
.B(n_663),
.C(n_662),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1112),
.B(n_666),
.Y(n_1325)
);

NOR2x1_ASAP7_75t_L g1326 ( 
.A(n_1106),
.B(n_585),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1128),
.B(n_676),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1169),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1112),
.B(n_677),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1163),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1204),
.A2(n_1010),
.B(n_1003),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1125),
.A2(n_702),
.B1(n_708),
.B2(n_679),
.Y(n_1332)
);

CKINVDCx10_ASAP7_75t_R g1333 ( 
.A(n_1114),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1162),
.Y(n_1334)
);

INVx4_ASAP7_75t_L g1335 ( 
.A(n_1177),
.Y(n_1335)
);

CKINVDCx8_ASAP7_75t_R g1336 ( 
.A(n_1106),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1144),
.Y(n_1337)
);

INVx5_ASAP7_75t_L g1338 ( 
.A(n_1106),
.Y(n_1338)
);

AND2x2_ASAP7_75t_SL g1339 ( 
.A(n_1237),
.B(n_585),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1145),
.B(n_709),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1167),
.B(n_712),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_SL g1342 ( 
.A(n_1131),
.B(n_588),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1183),
.B(n_713),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1131),
.B(n_716),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1102),
.B(n_717),
.Y(n_1345)
);

NAND2xp33_ASAP7_75t_L g1346 ( 
.A(n_1131),
.B(n_719),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1110),
.A2(n_699),
.B(n_700),
.C(n_696),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1166),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1169),
.B(n_1143),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1127),
.A2(n_1130),
.B(n_1129),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1129),
.A2(n_1028),
.B(n_1084),
.Y(n_1351)
);

OR2x6_ASAP7_75t_L g1352 ( 
.A(n_1166),
.B(n_705),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1198),
.B(n_731),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1234),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1150),
.B(n_733),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1130),
.A2(n_1085),
.B(n_707),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1156),
.B(n_740),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1115),
.B(n_588),
.Y(n_1358)
);

INVx5_ASAP7_75t_L g1359 ( 
.A(n_1207),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1099),
.B(n_745),
.Y(n_1360)
);

AND2x6_ASAP7_75t_L g1361 ( 
.A(n_1235),
.B(n_722),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1135),
.B(n_723),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1136),
.A2(n_727),
.B(n_725),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1136),
.A2(n_738),
.B(n_735),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1096),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1245),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1100),
.B(n_746),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1175),
.B(n_750),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1216),
.B(n_754),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1179),
.B(n_764),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1140),
.B(n_765),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1186),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1110),
.A2(n_749),
.B(n_753),
.C(n_747),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1189),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1234),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1208),
.A2(n_758),
.B(n_759),
.C(n_757),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1124),
.A2(n_601),
.B1(n_604),
.B2(n_597),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1124),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1111),
.A2(n_782),
.B(n_778),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1104),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1184),
.B(n_766),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1208),
.A2(n_791),
.B(n_786),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1111),
.A2(n_807),
.B(n_803),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1212),
.A2(n_821),
.B(n_814),
.Y(n_1384)
);

BUFx4f_ASAP7_75t_L g1385 ( 
.A(n_1166),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1119),
.A2(n_834),
.B(n_829),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1190),
.A2(n_769),
.B1(n_770),
.B2(n_767),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1211),
.A2(n_1133),
.B(n_1272),
.C(n_1221),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1172),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1219),
.A2(n_601),
.B(n_604),
.C(n_597),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1277),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1214),
.B(n_621),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1289),
.Y(n_1393)
);

CKINVDCx8_ASAP7_75t_R g1394 ( 
.A(n_1114),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1225),
.B(n_781),
.Y(n_1395)
);

INVx4_ASAP7_75t_L g1396 ( 
.A(n_1177),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1218),
.A2(n_790),
.B1(n_792),
.B2(n_787),
.Y(n_1397)
);

CKINVDCx6p67_ASAP7_75t_R g1398 ( 
.A(n_1187),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1201),
.Y(n_1399)
);

NOR3xp33_ASAP7_75t_L g1400 ( 
.A(n_1178),
.B(n_797),
.C(n_796),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1165),
.B(n_801),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1225),
.B(n_802),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1157),
.A2(n_622),
.B1(n_640),
.B2(n_621),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1203),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1209),
.A2(n_805),
.B(n_809),
.C(n_804),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1173),
.B(n_622),
.Y(n_1406)
);

BUFx8_ASAP7_75t_L g1407 ( 
.A(n_1151),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1210),
.A2(n_811),
.B(n_813),
.C(n_810),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1153),
.A2(n_819),
.B(n_815),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1229),
.A2(n_823),
.B(n_820),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1103),
.A2(n_827),
.B(n_661),
.Y(n_1411)
);

AO21x1_ASAP7_75t_L g1412 ( 
.A1(n_1249),
.A2(n_26),
.B(n_27),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1152),
.A2(n_661),
.B(n_640),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1291),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1270),
.B(n_688),
.C(n_669),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1154),
.A2(n_688),
.B(n_669),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1137),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1193),
.B(n_710),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1219),
.A2(n_752),
.B(n_710),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1139),
.B(n_752),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1168),
.B(n_761),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1182),
.A2(n_763),
.B(n_761),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1187),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1171),
.B(n_763),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1174),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1170),
.A2(n_824),
.B(n_406),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1195),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1231),
.B(n_824),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1142),
.B(n_26),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1107),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1187),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1123),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1262),
.B(n_29),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1269),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1217),
.B(n_30),
.Y(n_1435)
);

OAI21xp33_ASAP7_75t_L g1436 ( 
.A1(n_1195),
.A2(n_1222),
.B(n_1221),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1268),
.B(n_33),
.Y(n_1437)
);

OAI321xp33_ASAP7_75t_L g1438 ( 
.A1(n_1196),
.A2(n_38),
.A3(n_40),
.B1(n_35),
.B2(n_37),
.C(n_39),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1196),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1114),
.Y(n_1440)
);

INVxp67_ASAP7_75t_L g1441 ( 
.A(n_1134),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1290),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1122),
.B(n_35),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1282),
.B(n_37),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_SL g1445 ( 
.A(n_1213),
.B(n_415),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1160),
.B(n_40),
.Y(n_1446)
);

AND2x6_ASAP7_75t_L g1447 ( 
.A(n_1222),
.B(n_422),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1226),
.Y(n_1448)
);

OAI321xp33_ASAP7_75t_L g1449 ( 
.A1(n_1197),
.A2(n_43),
.A3(n_47),
.B1(n_41),
.B2(n_42),
.C(n_46),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1287),
.B(n_42),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1200),
.B(n_46),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1197),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1180),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1141),
.B(n_48),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1146),
.B(n_49),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1230),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1147),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_1457)
);

AO21x1_ASAP7_75t_L g1458 ( 
.A1(n_1252),
.A2(n_51),
.B(n_52),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1206),
.B(n_53),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1199),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1158),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1132),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_1462)
);

NOR2x1_ASAP7_75t_L g1463 ( 
.A(n_1278),
.B(n_54),
.Y(n_1463)
);

OR2x6_ASAP7_75t_L g1464 ( 
.A(n_1158),
.B(n_55),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1223),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1149),
.B(n_1159),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1199),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1113),
.B(n_58),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1223),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1241),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1164),
.A2(n_1121),
.B(n_1120),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1224),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1117),
.B(n_60),
.Y(n_1473)
);

BUFx4f_ASAP7_75t_L g1474 ( 
.A(n_1158),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1224),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1241),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1192),
.B(n_61),
.Y(n_1477)
);

INVx8_ASAP7_75t_L g1478 ( 
.A(n_1269),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1227),
.Y(n_1479)
);

AO21x1_ASAP7_75t_L g1480 ( 
.A1(n_1244),
.A2(n_63),
.B(n_64),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1269),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1236),
.B(n_65),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1202),
.B(n_66),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1238),
.B(n_67),
.Y(n_1484)
);

NOR3xp33_ASAP7_75t_L g1485 ( 
.A(n_1228),
.B(n_68),
.C(n_69),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1253),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1243),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1242),
.B(n_70),
.Y(n_1488)
);

A2O1A1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1247),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1247),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1275),
.B(n_1281),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1276),
.Y(n_1492)
);

O2A1O1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1248),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_1493)
);

AND2x6_ASAP7_75t_L g1494 ( 
.A(n_1251),
.B(n_1255),
.Y(n_1494)
);

O2A1O1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1255),
.A2(n_1259),
.B(n_1260),
.C(n_1256),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1288),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1265),
.Y(n_1497)
);

INVx4_ASAP7_75t_L g1498 ( 
.A(n_1288),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1256),
.A2(n_1260),
.B(n_1259),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1264),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1293),
.B(n_1233),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1266),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1267),
.A2(n_86),
.B1(n_82),
.B2(n_85),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1267),
.Y(n_1504)
);

A2O1A1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1271),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1271),
.B(n_87),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1274),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1274),
.B(n_89),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1250),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1279),
.Y(n_1510)
);

BUFx4f_ASAP7_75t_L g1511 ( 
.A(n_1298),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1279),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1512)
);

OAI21xp33_ASAP7_75t_L g1513 ( 
.A1(n_1292),
.A2(n_1295),
.B(n_1294),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1292),
.B(n_90),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1294),
.B(n_93),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1250),
.B(n_1261),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1295),
.B(n_94),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1296),
.A2(n_97),
.B(n_94),
.C(n_96),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1261),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1297),
.A2(n_458),
.B(n_455),
.Y(n_1520)
);

AOI21xp33_ASAP7_75t_L g1521 ( 
.A1(n_1293),
.A2(n_1258),
.B(n_1254),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1263),
.B(n_98),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1280),
.A2(n_465),
.B(n_462),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1283),
.B(n_98),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_1286),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1246),
.B(n_100),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1257),
.B(n_101),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1273),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1285),
.Y(n_1529)
);

A2O1A1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1350),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_1530)
);

OA22x2_ASAP7_75t_L g1531 ( 
.A1(n_1317),
.A2(n_111),
.B1(n_107),
.B2(n_110),
.Y(n_1531)
);

OAI22x1_ASAP7_75t_L g1532 ( 
.A1(n_1358),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1337),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1460),
.B(n_1467),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1389),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1300),
.Y(n_1536)
);

AOI21xp33_ASAP7_75t_L g1537 ( 
.A1(n_1318),
.A2(n_113),
.B(n_117),
.Y(n_1537)
);

A2O1A1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1495),
.A2(n_119),
.B(n_113),
.C(n_117),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1334),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1414),
.B(n_119),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1500),
.B(n_120),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1507),
.B(n_120),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1299),
.B(n_121),
.Y(n_1543)
);

O2A1O1Ixp5_ASAP7_75t_L g1544 ( 
.A1(n_1302),
.A2(n_483),
.B(n_484),
.C(n_482),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1314),
.Y(n_1545)
);

NAND2x1p5_ASAP7_75t_L g1546 ( 
.A(n_1313),
.B(n_122),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_SL g1547 ( 
.A1(n_1523),
.A2(n_123),
.B(n_124),
.Y(n_1547)
);

A2O1A1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1388),
.A2(n_126),
.B(n_124),
.C(n_125),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1478),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1313),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1417),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1478),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1425),
.Y(n_1553)
);

OAI22x1_ASAP7_75t_L g1554 ( 
.A1(n_1326),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1352),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1391),
.B(n_130),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1303),
.B(n_131),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1392),
.B(n_132),
.Y(n_1558)
);

AO31x2_ASAP7_75t_L g1559 ( 
.A1(n_1480),
.A2(n_136),
.A3(n_134),
.B(n_135),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1466),
.A2(n_141),
.B(n_142),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1407),
.Y(n_1561)
);

INVx5_ASAP7_75t_L g1562 ( 
.A(n_1478),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1372),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1434),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1339),
.B(n_141),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1393),
.B(n_142),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1356),
.A2(n_144),
.B(n_145),
.Y(n_1567)
);

AOI21xp33_ASAP7_75t_L g1568 ( 
.A1(n_1316),
.A2(n_146),
.B(n_148),
.Y(n_1568)
);

A2O1A1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1436),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_1569)
);

OAI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1469),
.A2(n_152),
.B(n_153),
.Y(n_1570)
);

NAND2x1p5_ASAP7_75t_L g1571 ( 
.A(n_1492),
.B(n_154),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1361),
.B(n_1349),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1472),
.A2(n_155),
.B(n_156),
.Y(n_1573)
);

INVxp67_ASAP7_75t_SL g1574 ( 
.A(n_1342),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1374),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_R g1576 ( 
.A(n_1336),
.B(n_155),
.Y(n_1576)
);

OAI21x1_ASAP7_75t_L g1577 ( 
.A1(n_1331),
.A2(n_156),
.B(n_157),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_L g1578 ( 
.A(n_1441),
.B(n_157),
.C(n_158),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1342),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1361),
.B(n_163),
.Y(n_1580)
);

A2O1A1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1436),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_1581)
);

CKINVDCx16_ASAP7_75t_R g1582 ( 
.A(n_1352),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1361),
.B(n_164),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1442),
.B(n_168),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1347),
.B(n_169),
.Y(n_1585)
);

OAI22x1_ASAP7_75t_L g1586 ( 
.A1(n_1415),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_1586)
);

O2A1O1Ixp5_ASAP7_75t_L g1587 ( 
.A1(n_1483),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1399),
.Y(n_1588)
);

OAI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1499),
.A2(n_176),
.B(n_177),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1373),
.B(n_178),
.Y(n_1590)
);

A2O1A1Ixp33_ASAP7_75t_L g1591 ( 
.A1(n_1493),
.A2(n_179),
.B(n_180),
.C(n_181),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1384),
.B(n_182),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1308),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1404),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1365),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1384),
.B(n_186),
.Y(n_1596)
);

AOI21xp33_ASAP7_75t_L g1597 ( 
.A1(n_1310),
.A2(n_188),
.B(n_189),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1376),
.B(n_189),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1470),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1502),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1481),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1504),
.A2(n_191),
.B(n_193),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1407),
.Y(n_1603)
);

NOR2x1_ASAP7_75t_SL g1604 ( 
.A(n_1352),
.B(n_194),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1363),
.B(n_1364),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1385),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1380),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1315),
.Y(n_1608)
);

A2O1A1Ixp33_ASAP7_75t_L g1609 ( 
.A1(n_1518),
.A2(n_1475),
.B(n_1383),
.C(n_1379),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1315),
.B(n_196),
.Y(n_1610)
);

NAND2x1_ASAP7_75t_L g1611 ( 
.A(n_1328),
.B(n_197),
.Y(n_1611)
);

NAND2x1p5_ASAP7_75t_L g1612 ( 
.A(n_1492),
.B(n_201),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1304),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1415),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.C(n_204),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1324),
.B(n_206),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1476),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1510),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1309),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_1618)
);

AOI221xp5_ASAP7_75t_L g1619 ( 
.A1(n_1390),
.A2(n_213),
.B1(n_214),
.B2(n_216),
.C(n_218),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1323),
.Y(n_1620)
);

AO31x2_ASAP7_75t_L g1621 ( 
.A1(n_1412),
.A2(n_214),
.A3(n_219),
.B(n_221),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1456),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1481),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1513),
.A2(n_224),
.B(n_225),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1312),
.B(n_226),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1487),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1351),
.A2(n_226),
.B(n_228),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1435),
.B(n_229),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1311),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_1629)
);

AOI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1378),
.A2(n_230),
.B1(n_233),
.B2(n_234),
.C(n_235),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1509),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1378),
.B(n_233),
.Y(n_1632)
);

NAND2x1p5_ASAP7_75t_L g1633 ( 
.A(n_1498),
.B(n_236),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1338),
.B(n_236),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1382),
.A2(n_237),
.B(n_238),
.Y(n_1635)
);

AO21x2_ASAP7_75t_L g1636 ( 
.A1(n_1520),
.A2(n_241),
.B(n_242),
.Y(n_1636)
);

AND3x4_ASAP7_75t_L g1637 ( 
.A(n_1333),
.B(n_242),
.C(n_243),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1398),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1403),
.B(n_246),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1395),
.B(n_249),
.Y(n_1640)
);

NAND2x1p5_ASAP7_75t_L g1641 ( 
.A(n_1498),
.B(n_250),
.Y(n_1641)
);

INVx5_ASAP7_75t_L g1642 ( 
.A(n_1509),
.Y(n_1642)
);

A2O1A1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1382),
.A2(n_252),
.B(n_253),
.C(n_255),
.Y(n_1643)
);

AND3x4_ASAP7_75t_L g1644 ( 
.A(n_1400),
.B(n_253),
.C(n_255),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1489),
.A2(n_256),
.B(n_257),
.C(n_259),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1311),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1455),
.A2(n_256),
.B(n_257),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1402),
.B(n_259),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1420),
.B(n_260),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_SL g1650 ( 
.A1(n_1426),
.A2(n_260),
.B(n_262),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1491),
.A2(n_263),
.B(n_264),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1525),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_1652)
);

AND2x2_ASAP7_75t_SL g1653 ( 
.A(n_1445),
.B(n_267),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1496),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1377),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1421),
.B(n_1424),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1494),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1410),
.B(n_274),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1451),
.A2(n_274),
.B(n_275),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1506),
.A2(n_277),
.B(n_278),
.Y(n_1660)
);

AOI222xp33_ASAP7_75t_L g1661 ( 
.A1(n_1474),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.C1(n_283),
.C2(n_284),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1410),
.B(n_282),
.Y(n_1662)
);

AOI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1319),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.C(n_289),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1508),
.A2(n_287),
.B(n_289),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1515),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1517),
.A2(n_290),
.B(n_291),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1322),
.A2(n_292),
.B(n_293),
.Y(n_1667)
);

AO31x2_ASAP7_75t_L g1668 ( 
.A1(n_1458),
.A2(n_293),
.A3(n_294),
.B(n_295),
.Y(n_1668)
);

BUFx4f_ASAP7_75t_L g1669 ( 
.A(n_1464),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1320),
.B(n_295),
.Y(n_1670)
);

NAND2x1p5_ASAP7_75t_L g1671 ( 
.A(n_1354),
.B(n_297),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1307),
.B(n_1419),
.Y(n_1672)
);

AO31x2_ASAP7_75t_L g1673 ( 
.A1(n_1505),
.A2(n_298),
.A3(n_299),
.B(n_301),
.Y(n_1673)
);

A2O1A1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1465),
.A2(n_298),
.B(n_299),
.C(n_301),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1419),
.B(n_303),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1433),
.A2(n_305),
.B(n_306),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1494),
.A2(n_306),
.B(n_307),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1437),
.A2(n_307),
.B(n_308),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1341),
.B(n_309),
.Y(n_1679)
);

AOI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1459),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.C(n_313),
.Y(n_1680)
);

OAI21xp33_ASAP7_75t_L g1681 ( 
.A1(n_1306),
.A2(n_310),
.B(n_313),
.Y(n_1681)
);

INVx5_ASAP7_75t_L g1682 ( 
.A(n_1509),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1327),
.B(n_314),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1340),
.B(n_1343),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1494),
.A2(n_315),
.B(n_316),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1359),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1345),
.B(n_320),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1362),
.B(n_323),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1405),
.A2(n_324),
.B(n_325),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1406),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_1690)
);

A2O1A1Ixp33_ASAP7_75t_L g1691 ( 
.A1(n_1473),
.A2(n_327),
.B(n_328),
.C(n_329),
.Y(n_1691)
);

AO31x2_ASAP7_75t_L g1692 ( 
.A1(n_1490),
.A2(n_327),
.A3(n_329),
.B(n_330),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1477),
.B(n_330),
.Y(n_1693)
);

OAI21xp33_ASAP7_75t_L g1694 ( 
.A1(n_1355),
.A2(n_331),
.B(n_333),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1362),
.B(n_334),
.Y(n_1695)
);

AOI21xp33_ASAP7_75t_L g1696 ( 
.A1(n_1353),
.A2(n_335),
.B(n_336),
.Y(n_1696)
);

INVx5_ASAP7_75t_L g1697 ( 
.A(n_1519),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1418),
.B(n_338),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1444),
.A2(n_339),
.B(n_340),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1381),
.B(n_339),
.Y(n_1700)
);

AO31x2_ASAP7_75t_L g1701 ( 
.A1(n_1503),
.A2(n_340),
.A3(n_341),
.B(n_342),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1429),
.A2(n_1521),
.B(n_1370),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1484),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1368),
.A2(n_343),
.B(n_345),
.Y(n_1704)
);

OAI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1408),
.A2(n_346),
.B(n_347),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1477),
.B(n_349),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1422),
.B(n_349),
.Y(n_1707)
);

OAI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1386),
.A2(n_350),
.B(n_351),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1430),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1360),
.B(n_354),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1423),
.B(n_354),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1432),
.Y(n_1712)
);

AO21x1_ASAP7_75t_L g1713 ( 
.A1(n_1522),
.A2(n_355),
.B(n_357),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1367),
.B(n_1401),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1357),
.B(n_1468),
.Y(n_1715)
);

AO21x1_ASAP7_75t_L g1716 ( 
.A1(n_1524),
.A2(n_358),
.B(n_359),
.Y(n_1716)
);

NAND3xp33_ASAP7_75t_L g1717 ( 
.A(n_1443),
.B(n_358),
.C(n_359),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1462),
.Y(n_1718)
);

A2O1A1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1438),
.A2(n_360),
.B(n_361),
.C(n_362),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1471),
.A2(n_363),
.B(n_364),
.Y(n_1720)
);

A2O1A1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1438),
.A2(n_365),
.B(n_366),
.C(n_367),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1323),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1529),
.A2(n_365),
.B(n_368),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1385),
.B(n_369),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1514),
.A2(n_369),
.B(n_370),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1413),
.B(n_370),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1387),
.B(n_1332),
.Y(n_1727)
);

A2O1A1Ixp33_ASAP7_75t_L g1728 ( 
.A1(n_1449),
.A2(n_374),
.B(n_375),
.C(n_376),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1416),
.B(n_377),
.Y(n_1729)
);

BUFx12f_ASAP7_75t_L g1730 ( 
.A(n_1335),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1519),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1371),
.A2(n_378),
.B(n_379),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1488),
.A2(n_379),
.B(n_380),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1338),
.B(n_381),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1454),
.Y(n_1735)
);

NOR2x1_ASAP7_75t_L g1736 ( 
.A(n_1335),
.B(n_383),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1330),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1397),
.B(n_383),
.Y(n_1738)
);

A2O1A1Ixp33_ASAP7_75t_L g1739 ( 
.A1(n_1449),
.A2(n_384),
.B(n_385),
.C(n_386),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1409),
.A2(n_384),
.B(n_385),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1411),
.B(n_1369),
.Y(n_1741)
);

NAND2x1p5_ASAP7_75t_L g1742 ( 
.A(n_1375),
.B(n_389),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_1394),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1446),
.B(n_387),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1446),
.B(n_387),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1526),
.A2(n_388),
.B(n_1527),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1448),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1516),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1501),
.A2(n_1305),
.B(n_1463),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1486),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_SL g1751 ( 
.A1(n_1486),
.A2(n_1497),
.B(n_1454),
.Y(n_1751)
);

AOI21xp33_ASAP7_75t_L g1752 ( 
.A1(n_1301),
.A2(n_1346),
.B(n_1325),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1482),
.A2(n_1329),
.B(n_1344),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1431),
.A2(n_1445),
.B1(n_1366),
.B2(n_1440),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1479),
.B(n_1348),
.Y(n_1755)
);

AO31x2_ASAP7_75t_L g1756 ( 
.A1(n_1512),
.A2(n_1457),
.A3(n_1453),
.B(n_1528),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1479),
.B(n_1338),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1450),
.B(n_1321),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1511),
.B(n_1485),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1511),
.B(n_1396),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1464),
.B(n_1474),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1497),
.B(n_1396),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1464),
.B(n_1461),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1447),
.A2(n_1350),
.B(n_1094),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1317),
.B(n_1097),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1478),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1427),
.B(n_1439),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1337),
.Y(n_1768)
);

OAI22x1_ASAP7_75t_L g1769 ( 
.A1(n_1317),
.A2(n_1214),
.B1(n_1108),
.B2(n_1237),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1427),
.B(n_1439),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1337),
.Y(n_1771)
);

AO31x2_ASAP7_75t_L g1772 ( 
.A1(n_1480),
.A2(n_1232),
.A3(n_1240),
.B(n_1239),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1337),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1314),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1427),
.B(n_1439),
.Y(n_1775)
);

NOR2x1_ASAP7_75t_SL g1776 ( 
.A(n_1352),
.B(n_1299),
.Y(n_1776)
);

AOI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1415),
.A2(n_1191),
.B1(n_1015),
.B2(n_1211),
.C(n_1133),
.Y(n_1777)
);

BUFx6f_ASAP7_75t_L g1778 ( 
.A(n_1478),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1350),
.A2(n_1094),
.B(n_1185),
.Y(n_1779)
);

A2O1A1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1350),
.A2(n_1495),
.B(n_1388),
.C(n_1439),
.Y(n_1780)
);

AOI21xp33_ASAP7_75t_L g1781 ( 
.A1(n_1358),
.A2(n_1318),
.B(n_1009),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1427),
.A2(n_1452),
.B1(n_1460),
.B2(n_1439),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1333),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1350),
.A2(n_1094),
.B(n_1185),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1317),
.B(n_1097),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1317),
.B(n_1097),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1350),
.A2(n_1094),
.B(n_1185),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1317),
.B(n_1097),
.Y(n_1788)
);

NAND2x1p5_ASAP7_75t_L g1789 ( 
.A(n_1313),
.B(n_1299),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1427),
.B(n_1439),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1427),
.A2(n_1452),
.B1(n_1460),
.B2(n_1439),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1337),
.Y(n_1792)
);

AO31x2_ASAP7_75t_L g1793 ( 
.A1(n_1480),
.A2(n_1232),
.A3(n_1240),
.B(n_1239),
.Y(n_1793)
);

NAND2x1p5_ASAP7_75t_L g1794 ( 
.A(n_1313),
.B(n_1299),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1299),
.B(n_1303),
.Y(n_1795)
);

AO31x2_ASAP7_75t_L g1796 ( 
.A1(n_1480),
.A2(n_1232),
.A3(n_1240),
.B(n_1239),
.Y(n_1796)
);

AND2x6_ASAP7_75t_L g1797 ( 
.A(n_1299),
.B(n_1354),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1337),
.Y(n_1798)
);

A2O1A1Ixp33_ASAP7_75t_L g1799 ( 
.A1(n_1350),
.A2(n_1495),
.B(n_1388),
.C(n_1439),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1300),
.Y(n_1800)
);

NAND2xp33_ASAP7_75t_SL g1801 ( 
.A(n_1492),
.B(n_951),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1337),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1337),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1427),
.B(n_1439),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1337),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1299),
.B(n_1303),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1337),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1427),
.B(n_1439),
.Y(n_1808)
);

BUFx3_ASAP7_75t_L g1809 ( 
.A(n_1314),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1414),
.B(n_951),
.Y(n_1810)
);

INVx5_ASAP7_75t_L g1811 ( 
.A(n_1478),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1427),
.B(n_1439),
.Y(n_1812)
);

AOI21xp33_ASAP7_75t_L g1813 ( 
.A1(n_1358),
.A2(n_1318),
.B(n_1009),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1427),
.B(n_1439),
.Y(n_1814)
);

AO31x2_ASAP7_75t_L g1815 ( 
.A1(n_1480),
.A2(n_1232),
.A3(n_1240),
.B(n_1239),
.Y(n_1815)
);

A2O1A1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1350),
.A2(n_1495),
.B(n_1388),
.C(n_1439),
.Y(n_1816)
);

NOR2xp67_ASAP7_75t_L g1817 ( 
.A(n_1338),
.B(n_1335),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1427),
.B(n_1439),
.Y(n_1818)
);

AND2x2_ASAP7_75t_SL g1819 ( 
.A(n_1313),
.B(n_1272),
.Y(n_1819)
);

A2O1A1Ixp33_ASAP7_75t_L g1820 ( 
.A1(n_1350),
.A2(n_1495),
.B(n_1388),
.C(n_1439),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1337),
.Y(n_1821)
);

NAND2xp33_ASAP7_75t_L g1822 ( 
.A(n_1478),
.B(n_1138),
.Y(n_1822)
);

NAND2xp33_ASAP7_75t_SL g1823 ( 
.A(n_1492),
.B(n_951),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1478),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1299),
.B(n_1303),
.Y(n_1825)
);

A2O1A1Ixp33_ASAP7_75t_L g1826 ( 
.A1(n_1350),
.A2(n_1495),
.B(n_1388),
.C(n_1439),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1773),
.Y(n_1827)
);

INVx4_ASAP7_75t_L g1828 ( 
.A(n_1562),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1599),
.Y(n_1829)
);

INVx2_ASAP7_75t_SL g1830 ( 
.A(n_1562),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1582),
.B(n_1765),
.Y(n_1831)
);

CKINVDCx20_ASAP7_75t_R g1832 ( 
.A(n_1783),
.Y(n_1832)
);

OR2x6_ASAP7_75t_L g1833 ( 
.A(n_1561),
.B(n_1603),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1539),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_SL g1835 ( 
.A1(n_1653),
.A2(n_1669),
.B1(n_1565),
.B2(n_1604),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1616),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1562),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1626),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_1555),
.Y(n_1839)
);

OAI21x1_ASAP7_75t_L g1840 ( 
.A1(n_1779),
.A2(n_1787),
.B(n_1784),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1792),
.Y(n_1841)
);

BUFx3_ASAP7_75t_L g1842 ( 
.A(n_1562),
.Y(n_1842)
);

INVx3_ASAP7_75t_L g1843 ( 
.A(n_1811),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1798),
.Y(n_1844)
);

CKINVDCx6p67_ASAP7_75t_R g1845 ( 
.A(n_1730),
.Y(n_1845)
);

NAND2x1p5_ASAP7_75t_L g1846 ( 
.A(n_1811),
.B(n_1552),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1811),
.B(n_1534),
.Y(n_1847)
);

BUFx3_ASAP7_75t_L g1848 ( 
.A(n_1811),
.Y(n_1848)
);

INVx3_ASAP7_75t_L g1849 ( 
.A(n_1552),
.Y(n_1849)
);

INVx5_ASAP7_75t_SL g1850 ( 
.A(n_1552),
.Y(n_1850)
);

NAND2x1_ASAP7_75t_L g1851 ( 
.A(n_1797),
.B(n_1751),
.Y(n_1851)
);

O2A1O1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1691),
.A2(n_1538),
.B(n_1548),
.C(n_1643),
.Y(n_1852)
);

BUFx6f_ASAP7_75t_SL g1853 ( 
.A(n_1743),
.Y(n_1853)
);

OAI21x1_ASAP7_75t_SL g1854 ( 
.A1(n_1677),
.A2(n_1685),
.B(n_1776),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1777),
.B(n_1718),
.Y(n_1855)
);

OA21x2_ASAP7_75t_L g1856 ( 
.A1(n_1780),
.A2(n_1816),
.B(n_1799),
.Y(n_1856)
);

AOI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1780),
.A2(n_1816),
.B(n_1799),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1767),
.B(n_1770),
.Y(n_1858)
);

NAND2x1_ASAP7_75t_L g1859 ( 
.A(n_1797),
.B(n_1631),
.Y(n_1859)
);

AO21x2_ASAP7_75t_L g1860 ( 
.A1(n_1820),
.A2(n_1826),
.B(n_1636),
.Y(n_1860)
);

INVx4_ASAP7_75t_L g1861 ( 
.A(n_1552),
.Y(n_1861)
);

OA21x2_ASAP7_75t_L g1862 ( 
.A1(n_1820),
.A2(n_1826),
.B(n_1544),
.Y(n_1862)
);

CKINVDCx20_ASAP7_75t_R g1863 ( 
.A(n_1669),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1802),
.Y(n_1864)
);

NAND3xp33_ASAP7_75t_L g1865 ( 
.A(n_1538),
.B(n_1548),
.C(n_1530),
.Y(n_1865)
);

OR3x4_ASAP7_75t_SL g1866 ( 
.A(n_1574),
.B(n_1637),
.C(n_1644),
.Y(n_1866)
);

INVx8_ASAP7_75t_L g1867 ( 
.A(n_1797),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1672),
.B(n_1781),
.Y(n_1868)
);

CKINVDCx6p67_ASAP7_75t_R g1869 ( 
.A(n_1550),
.Y(n_1869)
);

BUFx2_ASAP7_75t_R g1870 ( 
.A(n_1545),
.Y(n_1870)
);

AOI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1785),
.A2(n_1788),
.B1(n_1786),
.B2(n_1777),
.Y(n_1871)
);

CKINVDCx20_ASAP7_75t_R g1872 ( 
.A(n_1576),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1782),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1791),
.B(n_1589),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1813),
.B(n_1727),
.Y(n_1875)
);

BUFx3_ASAP7_75t_L g1876 ( 
.A(n_1778),
.Y(n_1876)
);

BUFx3_ASAP7_75t_L g1877 ( 
.A(n_1778),
.Y(n_1877)
);

BUFx3_ASAP7_75t_L g1878 ( 
.A(n_1778),
.Y(n_1878)
);

BUFx12f_ASAP7_75t_L g1879 ( 
.A(n_1638),
.Y(n_1879)
);

BUFx2_ASAP7_75t_L g1880 ( 
.A(n_1800),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1805),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1807),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1656),
.B(n_1775),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1790),
.B(n_1804),
.Y(n_1884)
);

OA21x2_ASAP7_75t_L g1885 ( 
.A1(n_1624),
.A2(n_1627),
.B(n_1577),
.Y(n_1885)
);

OAI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1684),
.A2(n_1609),
.B(n_1714),
.Y(n_1886)
);

AO21x2_ASAP7_75t_L g1887 ( 
.A1(n_1702),
.A2(n_1720),
.B(n_1609),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1808),
.Y(n_1888)
);

INVx6_ASAP7_75t_L g1889 ( 
.A(n_1778),
.Y(n_1889)
);

BUFx8_ASAP7_75t_L g1890 ( 
.A(n_1824),
.Y(n_1890)
);

BUFx5_ASAP7_75t_L g1891 ( 
.A(n_1797),
.Y(n_1891)
);

CKINVDCx16_ASAP7_75t_R g1892 ( 
.A(n_1576),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1812),
.B(n_1814),
.Y(n_1893)
);

BUFx2_ASAP7_75t_L g1894 ( 
.A(n_1824),
.Y(n_1894)
);

BUFx2_ASAP7_75t_R g1895 ( 
.A(n_1774),
.Y(n_1895)
);

BUFx3_ASAP7_75t_L g1896 ( 
.A(n_1824),
.Y(n_1896)
);

BUFx2_ASAP7_75t_R g1897 ( 
.A(n_1809),
.Y(n_1897)
);

OAI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1746),
.A2(n_1700),
.B(n_1702),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1533),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1818),
.B(n_1556),
.Y(n_1900)
);

BUFx2_ASAP7_75t_SL g1901 ( 
.A(n_1817),
.Y(n_1901)
);

CKINVDCx6p67_ASAP7_75t_R g1902 ( 
.A(n_1620),
.Y(n_1902)
);

BUFx2_ASAP7_75t_L g1903 ( 
.A(n_1824),
.Y(n_1903)
);

INVx1_ASAP7_75t_SL g1904 ( 
.A(n_1722),
.Y(n_1904)
);

INVx1_ASAP7_75t_SL g1905 ( 
.A(n_1543),
.Y(n_1905)
);

BUFx8_ASAP7_75t_L g1906 ( 
.A(n_1761),
.Y(n_1906)
);

NAND2x1p5_ASAP7_75t_L g1907 ( 
.A(n_1642),
.B(n_1682),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1535),
.Y(n_1908)
);

OAI21x1_ASAP7_75t_SL g1909 ( 
.A1(n_1635),
.A2(n_1602),
.B(n_1573),
.Y(n_1909)
);

CKINVDCx11_ASAP7_75t_R g1910 ( 
.A(n_1543),
.Y(n_1910)
);

INVx2_ASAP7_75t_SL g1911 ( 
.A(n_1789),
.Y(n_1911)
);

AND2x6_ASAP7_75t_L g1912 ( 
.A(n_1646),
.B(n_1557),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1605),
.A2(n_1746),
.B(n_1753),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1768),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1536),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1771),
.Y(n_1916)
);

BUFx2_ASAP7_75t_SL g1917 ( 
.A(n_1606),
.Y(n_1917)
);

AO21x2_ASAP7_75t_L g1918 ( 
.A1(n_1570),
.A2(n_1581),
.B(n_1569),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1803),
.Y(n_1919)
);

BUFx2_ASAP7_75t_SL g1920 ( 
.A(n_1642),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1821),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1551),
.Y(n_1922)
);

HB1xp67_ASAP7_75t_L g1923 ( 
.A(n_1642),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1556),
.B(n_1540),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1553),
.Y(n_1925)
);

INVx8_ASAP7_75t_L g1926 ( 
.A(n_1682),
.Y(n_1926)
);

INVx2_ASAP7_75t_SL g1927 ( 
.A(n_1789),
.Y(n_1927)
);

INVx1_ASAP7_75t_SL g1928 ( 
.A(n_1654),
.Y(n_1928)
);

AO21x2_ASAP7_75t_L g1929 ( 
.A1(n_1650),
.A2(n_1723),
.B(n_1705),
.Y(n_1929)
);

AND2x4_ASAP7_75t_SL g1930 ( 
.A(n_1549),
.B(n_1766),
.Y(n_1930)
);

OA21x2_ASAP7_75t_L g1931 ( 
.A1(n_1591),
.A2(n_1721),
.B(n_1719),
.Y(n_1931)
);

BUFx6f_ASAP7_75t_L g1932 ( 
.A(n_1631),
.Y(n_1932)
);

OAI21x1_ASAP7_75t_L g1933 ( 
.A1(n_1762),
.A2(n_1749),
.B(n_1611),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1595),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1613),
.B(n_1670),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1540),
.B(n_1558),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1536),
.B(n_1698),
.Y(n_1937)
);

BUFx3_ASAP7_75t_L g1938 ( 
.A(n_1682),
.Y(n_1938)
);

INVx1_ASAP7_75t_SL g1939 ( 
.A(n_1654),
.Y(n_1939)
);

HB1xp67_ASAP7_75t_L g1940 ( 
.A(n_1697),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1810),
.B(n_1608),
.Y(n_1941)
);

OA21x2_ASAP7_75t_L g1942 ( 
.A1(n_1591),
.A2(n_1721),
.B(n_1719),
.Y(n_1942)
);

OAI21x1_ASAP7_75t_L g1943 ( 
.A1(n_1733),
.A2(n_1567),
.B(n_1651),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1801),
.Y(n_1944)
);

BUFx2_ASAP7_75t_SL g1945 ( 
.A(n_1697),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1686),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1607),
.Y(n_1947)
);

AND2x4_ASAP7_75t_L g1948 ( 
.A(n_1697),
.B(n_1549),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1697),
.B(n_1766),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1671),
.Y(n_1950)
);

OAI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1700),
.A2(n_1715),
.B(n_1687),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1810),
.B(n_1665),
.Y(n_1952)
);

OA21x2_ASAP7_75t_L g1953 ( 
.A1(n_1728),
.A2(n_1739),
.B(n_1689),
.Y(n_1953)
);

INVx1_ASAP7_75t_SL g1954 ( 
.A(n_1686),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1769),
.B(n_1639),
.Y(n_1955)
);

INVx2_ASAP7_75t_SL g1956 ( 
.A(n_1794),
.Y(n_1956)
);

OR2x6_ASAP7_75t_L g1957 ( 
.A(n_1546),
.B(n_1557),
.Y(n_1957)
);

BUFx4f_ASAP7_75t_L g1958 ( 
.A(n_1546),
.Y(n_1958)
);

OA21x2_ASAP7_75t_L g1959 ( 
.A1(n_1660),
.A2(n_1666),
.B(n_1664),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1687),
.B(n_1707),
.Y(n_1960)
);

OAI21x1_ASAP7_75t_L g1961 ( 
.A1(n_1560),
.A2(n_1647),
.B(n_1659),
.Y(n_1961)
);

OA21x2_ASAP7_75t_L g1962 ( 
.A1(n_1667),
.A2(n_1681),
.B(n_1674),
.Y(n_1962)
);

O2A1O1Ixp33_ASAP7_75t_L g1963 ( 
.A1(n_1691),
.A2(n_1643),
.B(n_1645),
.C(n_1590),
.Y(n_1963)
);

AO21x2_ASAP7_75t_L g1964 ( 
.A1(n_1740),
.A2(n_1596),
.B(n_1592),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1735),
.B(n_1675),
.Y(n_1965)
);

NAND2x1p5_ASAP7_75t_L g1966 ( 
.A(n_1819),
.B(n_1564),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1671),
.Y(n_1967)
);

OAI21x1_ASAP7_75t_L g1968 ( 
.A1(n_1647),
.A2(n_1659),
.B(n_1676),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1738),
.B(n_1724),
.Y(n_1969)
);

OA21x2_ASAP7_75t_L g1970 ( 
.A1(n_1694),
.A2(n_1587),
.B(n_1676),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1795),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1742),
.Y(n_1972)
);

AO22x2_ASAP7_75t_L g1973 ( 
.A1(n_1574),
.A2(n_1637),
.B1(n_1693),
.B2(n_1706),
.Y(n_1973)
);

OAI21xp5_ASAP7_75t_L g1974 ( 
.A1(n_1649),
.A2(n_1679),
.B(n_1625),
.Y(n_1974)
);

NAND3xp33_ASAP7_75t_L g1975 ( 
.A(n_1619),
.B(n_1663),
.C(n_1578),
.Y(n_1975)
);

BUFx2_ASAP7_75t_SL g1976 ( 
.A(n_1634),
.Y(n_1976)
);

AOI22xp33_ASAP7_75t_SL g1977 ( 
.A1(n_1531),
.A2(n_1641),
.B1(n_1571),
.B2(n_1633),
.Y(n_1977)
);

OAI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1658),
.A2(n_1662),
.B(n_1683),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1742),
.Y(n_1979)
);

OAI21x1_ASAP7_75t_SL g1980 ( 
.A1(n_1580),
.A2(n_1583),
.B(n_1708),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1588),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1610),
.B(n_1584),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1622),
.B(n_1703),
.Y(n_1983)
);

AOI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1693),
.A2(n_1706),
.B1(n_1579),
.B2(n_1648),
.Y(n_1984)
);

CKINVDCx11_ASAP7_75t_R g1985 ( 
.A(n_1634),
.Y(n_1985)
);

OAI21x1_ASAP7_75t_L g1986 ( 
.A1(n_1678),
.A2(n_1699),
.B(n_1704),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1758),
.B(n_1572),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1741),
.B(n_1541),
.Y(n_1988)
);

CKINVDCx14_ASAP7_75t_R g1989 ( 
.A(n_1823),
.Y(n_1989)
);

OAI322xp33_ASAP7_75t_L g1990 ( 
.A1(n_1655),
.A2(n_1531),
.A3(n_1615),
.B1(n_1618),
.B2(n_1593),
.C1(n_1648),
.C2(n_1640),
.Y(n_1990)
);

AO21x2_ASAP7_75t_L g1991 ( 
.A1(n_1710),
.A2(n_1744),
.B(n_1745),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1563),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1741),
.B(n_1754),
.Y(n_1993)
);

CKINVDCx11_ASAP7_75t_R g1994 ( 
.A(n_1734),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1575),
.Y(n_1995)
);

CKINVDCx20_ASAP7_75t_R g1996 ( 
.A(n_1579),
.Y(n_1996)
);

OA21x2_ASAP7_75t_L g1997 ( 
.A1(n_1725),
.A2(n_1716),
.B(n_1713),
.Y(n_1997)
);

AOI21x1_ASAP7_75t_L g1998 ( 
.A1(n_1628),
.A2(n_1632),
.B(n_1566),
.Y(n_1998)
);

AO21x2_ASAP7_75t_L g1999 ( 
.A1(n_1585),
.A2(n_1695),
.B(n_1688),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1594),
.Y(n_2000)
);

OAI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_1542),
.A2(n_1729),
.B(n_1726),
.Y(n_2001)
);

NAND2x1p5_ASAP7_75t_L g2002 ( 
.A(n_1819),
.B(n_1564),
.Y(n_2002)
);

OAI21x1_ASAP7_75t_SL g2003 ( 
.A1(n_1732),
.A2(n_1629),
.B(n_1630),
.Y(n_2003)
);

OAI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1598),
.A2(n_1717),
.B(n_1759),
.Y(n_2004)
);

OAI21x1_ASAP7_75t_SL g2005 ( 
.A1(n_1630),
.A2(n_1663),
.B(n_1736),
.Y(n_2005)
);

AO21x2_ASAP7_75t_L g2006 ( 
.A1(n_1537),
.A2(n_1696),
.B(n_1597),
.Y(n_2006)
);

OA21x2_ASAP7_75t_L g2007 ( 
.A1(n_1657),
.A2(n_1680),
.B(n_1568),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1734),
.Y(n_2008)
);

OAI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1640),
.A2(n_1657),
.B(n_1709),
.Y(n_2009)
);

CKINVDCx11_ASAP7_75t_R g2010 ( 
.A(n_1795),
.Y(n_2010)
);

BUFx3_ASAP7_75t_L g2011 ( 
.A(n_1731),
.Y(n_2011)
);

AO22x2_ASAP7_75t_L g2012 ( 
.A1(n_1644),
.A2(n_1652),
.B1(n_1600),
.B2(n_1763),
.Y(n_2012)
);

AO31x2_ASAP7_75t_L g2013 ( 
.A1(n_1586),
.A2(n_1532),
.A3(n_1617),
.B(n_1554),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1712),
.Y(n_2014)
);

AOI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1757),
.A2(n_1755),
.B(n_1737),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1806),
.B(n_1825),
.Y(n_2016)
);

OAI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1747),
.A2(n_1690),
.B(n_1619),
.Y(n_2017)
);

OA21x2_ASAP7_75t_L g2018 ( 
.A1(n_1680),
.A2(n_1614),
.B(n_1815),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1711),
.B(n_1748),
.Y(n_2019)
);

BUFx10_ASAP7_75t_L g2020 ( 
.A(n_1806),
.Y(n_2020)
);

OAI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1614),
.A2(n_1752),
.B(n_1748),
.Y(n_2021)
);

NAND2x1p5_ASAP7_75t_L g2022 ( 
.A(n_1601),
.B(n_1623),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1760),
.A2(n_1623),
.B(n_1571),
.Y(n_2023)
);

AO21x2_ASAP7_75t_L g2024 ( 
.A1(n_1772),
.A2(n_1815),
.B(n_1796),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1825),
.B(n_1661),
.Y(n_2025)
);

AND2x4_ASAP7_75t_L g2026 ( 
.A(n_1750),
.B(n_1756),
.Y(n_2026)
);

INVx1_ASAP7_75t_SL g2027 ( 
.A(n_1822),
.Y(n_2027)
);

OAI21x1_ASAP7_75t_L g2028 ( 
.A1(n_1612),
.A2(n_1633),
.B(n_1641),
.Y(n_2028)
);

AOI22x1_ASAP7_75t_L g2029 ( 
.A1(n_1612),
.A2(n_1750),
.B1(n_1815),
.B2(n_1796),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1692),
.Y(n_2030)
);

NOR2xp67_ASAP7_75t_L g2031 ( 
.A(n_1750),
.B(n_1701),
.Y(n_2031)
);

AO21x2_ASAP7_75t_L g2032 ( 
.A1(n_1772),
.A2(n_1815),
.B(n_1796),
.Y(n_2032)
);

OAI21x1_ASAP7_75t_L g2033 ( 
.A1(n_1772),
.A2(n_1796),
.B(n_1793),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_L g2034 ( 
.A(n_1756),
.B(n_1793),
.Y(n_2034)
);

OAI21x1_ASAP7_75t_L g2035 ( 
.A1(n_1772),
.A2(n_1793),
.B(n_1559),
.Y(n_2035)
);

AO21x2_ASAP7_75t_L g2036 ( 
.A1(n_1559),
.A2(n_1621),
.B(n_1668),
.Y(n_2036)
);

INVx2_ASAP7_75t_SL g2037 ( 
.A(n_1692),
.Y(n_2037)
);

BUFx12f_ASAP7_75t_L g2038 ( 
.A(n_1692),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1692),
.Y(n_2039)
);

OA21x2_ASAP7_75t_L g2040 ( 
.A1(n_1559),
.A2(n_1621),
.B(n_1668),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1756),
.B(n_1673),
.Y(n_2041)
);

CKINVDCx20_ASAP7_75t_R g2042 ( 
.A(n_1701),
.Y(n_2042)
);

INVx6_ASAP7_75t_L g2043 ( 
.A(n_1701),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1673),
.Y(n_2044)
);

INVx3_ASAP7_75t_L g2045 ( 
.A(n_1673),
.Y(n_2045)
);

OA21x2_ASAP7_75t_L g2046 ( 
.A1(n_1621),
.A2(n_1668),
.B(n_1673),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1653),
.B(n_1677),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1773),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1672),
.B(n_1414),
.Y(n_2049)
);

INVx3_ASAP7_75t_L g2050 ( 
.A(n_1562),
.Y(n_2050)
);

AOI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_1764),
.A2(n_1799),
.B(n_1780),
.Y(n_2051)
);

INVx3_ASAP7_75t_L g2052 ( 
.A(n_1562),
.Y(n_2052)
);

CKINVDCx16_ASAP7_75t_R g2053 ( 
.A(n_1582),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1773),
.Y(n_2054)
);

NAND2x1p5_ASAP7_75t_L g2055 ( 
.A(n_1562),
.B(n_1811),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_L g2056 ( 
.A(n_1672),
.B(n_1414),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1777),
.B(n_1718),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1773),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1777),
.B(n_1718),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1765),
.B(n_1785),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_1672),
.B(n_1414),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1773),
.Y(n_2062)
);

OAI21x1_ASAP7_75t_SL g2063 ( 
.A1(n_1677),
.A2(n_1685),
.B(n_1547),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_1562),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1777),
.B(n_1718),
.Y(n_2065)
);

OAI21x1_ASAP7_75t_SL g2066 ( 
.A1(n_1677),
.A2(n_1685),
.B(n_1547),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1599),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1773),
.Y(n_2068)
);

BUFx2_ASAP7_75t_L g2069 ( 
.A(n_1582),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1764),
.A2(n_1799),
.B(n_1780),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_1582),
.B(n_1428),
.Y(n_2071)
);

AO222x2_ASAP7_75t_L g2072 ( 
.A1(n_1761),
.A2(n_1392),
.B1(n_1176),
.B2(n_1763),
.C1(n_1320),
.C2(n_1565),
.Y(n_2072)
);

INVx6_ASAP7_75t_L g2073 ( 
.A(n_1562),
.Y(n_2073)
);

NOR2xp33_ASAP7_75t_SL g2074 ( 
.A(n_1783),
.B(n_1313),
.Y(n_2074)
);

BUFx3_ASAP7_75t_L g2075 ( 
.A(n_1562),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1562),
.Y(n_2076)
);

INVxp67_ASAP7_75t_SL g2077 ( 
.A(n_1782),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1773),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1773),
.Y(n_2079)
);

INVxp33_ASAP7_75t_L g2080 ( 
.A(n_2055),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_1890),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1840),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_1858),
.B(n_1884),
.Y(n_2083)
);

INVx4_ASAP7_75t_SL g2084 ( 
.A(n_1912),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1983),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1899),
.Y(n_2086)
);

OAI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_2025),
.A2(n_1884),
.B1(n_1858),
.B2(n_1957),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1908),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_1890),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1888),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1914),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1916),
.Y(n_2092)
);

INVx2_ASAP7_75t_SL g2093 ( 
.A(n_1890),
.Y(n_2093)
);

BUFx3_ASAP7_75t_L g2094 ( 
.A(n_1926),
.Y(n_2094)
);

BUFx2_ASAP7_75t_L g2095 ( 
.A(n_2055),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_2049),
.B(n_2056),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2060),
.B(n_1969),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1919),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1921),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1934),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1947),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1922),
.Y(n_2102)
);

INVx2_ASAP7_75t_SL g2103 ( 
.A(n_1926),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_2026),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1925),
.Y(n_2105)
);

INVxp67_ASAP7_75t_L g2106 ( 
.A(n_1912),
.Y(n_2106)
);

HB1xp67_ASAP7_75t_L g2107 ( 
.A(n_2026),
.Y(n_2107)
);

INVx3_ASAP7_75t_L g2108 ( 
.A(n_2064),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1827),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_1884),
.B(n_1935),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1841),
.Y(n_2111)
);

AOI222xp33_ASAP7_75t_L g2112 ( 
.A1(n_2049),
.A2(n_2056),
.B1(n_2061),
.B2(n_1875),
.C1(n_1924),
.C2(n_1910),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1844),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2061),
.B(n_1855),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1864),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1881),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1882),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2048),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2054),
.Y(n_2119)
);

INVxp67_ASAP7_75t_L g2120 ( 
.A(n_1912),
.Y(n_2120)
);

BUFx3_ASAP7_75t_L g2121 ( 
.A(n_1926),
.Y(n_2121)
);

AOI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_1912),
.A2(n_1875),
.B1(n_1973),
.B2(n_1952),
.Y(n_2122)
);

AO21x2_ASAP7_75t_L g2123 ( 
.A1(n_2031),
.A2(n_2070),
.B(n_2051),
.Y(n_2123)
);

INVxp67_ASAP7_75t_L g2124 ( 
.A(n_1912),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2058),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2062),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2068),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1937),
.B(n_1871),
.Y(n_2128)
);

AND2x4_ASAP7_75t_L g2129 ( 
.A(n_1847),
.B(n_1957),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2078),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2079),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1981),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_2026),
.Y(n_2133)
);

AND2x4_ASAP7_75t_L g2134 ( 
.A(n_1847),
.B(n_1957),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1992),
.Y(n_2135)
);

HB1xp67_ASAP7_75t_SL g2136 ( 
.A(n_1976),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1995),
.Y(n_2137)
);

AOI22xp33_ASAP7_75t_SL g2138 ( 
.A1(n_1973),
.A2(n_2012),
.B1(n_1958),
.B2(n_1989),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2000),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2014),
.Y(n_2140)
);

CKINVDCx12_ASAP7_75t_R g2141 ( 
.A(n_1833),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1829),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1883),
.B(n_1955),
.Y(n_2143)
);

BUFx2_ASAP7_75t_L g2144 ( 
.A(n_1907),
.Y(n_2144)
);

BUFx3_ASAP7_75t_L g2145 ( 
.A(n_1907),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1836),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_2064),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1838),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_1915),
.B(n_1893),
.Y(n_2149)
);

HB1xp67_ASAP7_75t_L g2150 ( 
.A(n_1873),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1838),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2067),
.Y(n_2152)
);

AOI22xp33_ASAP7_75t_L g2153 ( 
.A1(n_1973),
.A2(n_1868),
.B1(n_2012),
.B2(n_1993),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2016),
.B(n_1952),
.Y(n_2154)
);

AOI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_1868),
.A2(n_2012),
.B1(n_1993),
.B2(n_1951),
.Y(n_2155)
);

AOI21xp5_ASAP7_75t_L g2156 ( 
.A1(n_1913),
.A2(n_1857),
.B(n_1898),
.Y(n_2156)
);

AOI22xp33_ASAP7_75t_L g2157 ( 
.A1(n_1835),
.A2(n_1977),
.B1(n_1960),
.B2(n_1886),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1847),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2028),
.Y(n_2159)
);

INVx2_ASAP7_75t_SL g2160 ( 
.A(n_1902),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2057),
.B(n_2059),
.Y(n_2161)
);

HB1xp67_ASAP7_75t_L g2162 ( 
.A(n_1873),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1920),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1945),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1923),
.Y(n_2165)
);

BUFx3_ASAP7_75t_L g2166 ( 
.A(n_1846),
.Y(n_2166)
);

OR2x2_ASAP7_75t_L g2167 ( 
.A(n_1831),
.B(n_1928),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1856),
.Y(n_2168)
);

BUFx4f_ASAP7_75t_SL g2169 ( 
.A(n_1845),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1923),
.Y(n_2170)
);

NOR2xp33_ASAP7_75t_L g2171 ( 
.A(n_2072),
.B(n_1900),
.Y(n_2171)
);

INVx1_ASAP7_75t_SL g2172 ( 
.A(n_2010),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1940),
.Y(n_2173)
);

BUFx2_ASAP7_75t_L g2174 ( 
.A(n_1846),
.Y(n_2174)
);

CKINVDCx9p33_ASAP7_75t_R g2175 ( 
.A(n_2069),
.Y(n_2175)
);

BUFx3_ASAP7_75t_L g2176 ( 
.A(n_2076),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1940),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1834),
.Y(n_2178)
);

AND2x4_ASAP7_75t_L g2179 ( 
.A(n_1948),
.B(n_1949),
.Y(n_2179)
);

AOI22xp33_ASAP7_75t_L g2180 ( 
.A1(n_1835),
.A2(n_1977),
.B1(n_2005),
.B2(n_2065),
.Y(n_2180)
);

HB1xp67_ASAP7_75t_L g2181 ( 
.A(n_1932),
.Y(n_2181)
);

AND2x4_ASAP7_75t_L g2182 ( 
.A(n_1948),
.B(n_1949),
.Y(n_2182)
);

AO21x1_ASAP7_75t_SL g2183 ( 
.A1(n_1950),
.A2(n_1972),
.B(n_1967),
.Y(n_2183)
);

AOI22xp33_ASAP7_75t_L g2184 ( 
.A1(n_1936),
.A2(n_1910),
.B1(n_2047),
.B2(n_2042),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1979),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1911),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1927),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_1939),
.B(n_1946),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1941),
.B(n_1987),
.Y(n_2189)
);

INVx3_ASAP7_75t_L g2190 ( 
.A(n_1867),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1956),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_1954),
.B(n_1880),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2008),
.Y(n_2193)
);

AOI22xp5_ASAP7_75t_L g2194 ( 
.A1(n_1941),
.A2(n_1872),
.B1(n_1987),
.B2(n_1996),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1958),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1842),
.Y(n_2196)
);

BUFx12f_ASAP7_75t_L g2197 ( 
.A(n_1985),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_1832),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1848),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1848),
.Y(n_2200)
);

BUFx2_ASAP7_75t_L g2201 ( 
.A(n_2075),
.Y(n_2201)
);

OAI22xp33_ASAP7_75t_L g2202 ( 
.A1(n_2077),
.A2(n_1905),
.B1(n_1984),
.B2(n_1892),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2075),
.Y(n_2203)
);

INVx3_ASAP7_75t_L g2204 ( 
.A(n_1867),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1901),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1860),
.Y(n_2206)
);

INVx3_ASAP7_75t_L g2207 ( 
.A(n_1867),
.Y(n_2207)
);

INVx2_ASAP7_75t_SL g2208 ( 
.A(n_2073),
.Y(n_2208)
);

OAI21x1_ASAP7_75t_SL g2209 ( 
.A1(n_1854),
.A2(n_2066),
.B(n_2063),
.Y(n_2209)
);

AOI22xp33_ASAP7_75t_L g2210 ( 
.A1(n_2042),
.A2(n_1990),
.B1(n_1975),
.B2(n_1985),
.Y(n_2210)
);

AOI22xp33_ASAP7_75t_L g2211 ( 
.A1(n_1994),
.A2(n_2038),
.B1(n_1865),
.B2(n_1874),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1843),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2071),
.B(n_1965),
.Y(n_2213)
);

AOI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_1872),
.A2(n_1996),
.B1(n_1994),
.B2(n_1863),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1843),
.Y(n_2215)
);

INVx2_ASAP7_75t_SL g2216 ( 
.A(n_2073),
.Y(n_2216)
);

BUFx3_ASAP7_75t_L g2217 ( 
.A(n_2073),
.Y(n_2217)
);

CKINVDCx9p33_ASAP7_75t_R g2218 ( 
.A(n_1989),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2050),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2053),
.B(n_1904),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_1839),
.B(n_1971),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2050),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2052),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2034),
.B(n_1982),
.Y(n_2224)
);

BUFx2_ASAP7_75t_L g2225 ( 
.A(n_1828),
.Y(n_2225)
);

AOI21xp33_ASAP7_75t_SL g2226 ( 
.A1(n_1944),
.A2(n_1833),
.B(n_1830),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2020),
.B(n_2010),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2020),
.B(n_1894),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2052),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1837),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2013),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1885),
.Y(n_2232)
);

AOI22xp33_ASAP7_75t_L g2233 ( 
.A1(n_2038),
.A2(n_2077),
.B1(n_2003),
.B2(n_2034),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_1903),
.B(n_1850),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_1850),
.B(n_1861),
.Y(n_2235)
);

NOR2xp33_ASAP7_75t_R g2236 ( 
.A(n_1863),
.B(n_2074),
.Y(n_2236)
);

INVx3_ASAP7_75t_L g2237 ( 
.A(n_1828),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2013),
.Y(n_2238)
);

INVxp67_ASAP7_75t_SL g2239 ( 
.A(n_2037),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2013),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2030),
.Y(n_2241)
);

INVx6_ASAP7_75t_L g2242 ( 
.A(n_1861),
.Y(n_2242)
);

INVx1_ASAP7_75t_SL g2243 ( 
.A(n_1870),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2039),
.Y(n_2244)
);

AOI22xp33_ASAP7_75t_L g2245 ( 
.A1(n_1988),
.A2(n_2017),
.B1(n_2018),
.B2(n_1909),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2019),
.B(n_1850),
.Y(n_2246)
);

AOI21xp33_ASAP7_75t_L g2247 ( 
.A1(n_2006),
.A2(n_1980),
.B(n_1963),
.Y(n_2247)
);

INVx4_ASAP7_75t_L g2248 ( 
.A(n_1869),
.Y(n_2248)
);

INVx3_ASAP7_75t_L g2249 ( 
.A(n_1938),
.Y(n_2249)
);

AOI221xp5_ASAP7_75t_L g2250 ( 
.A1(n_1852),
.A2(n_1963),
.B1(n_2001),
.B2(n_1974),
.C(n_2041),
.Y(n_2250)
);

CKINVDCx8_ASAP7_75t_R g2251 ( 
.A(n_1866),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2041),
.B(n_1906),
.Y(n_2252)
);

INVx2_ASAP7_75t_SL g2253 ( 
.A(n_1889),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2023),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1917),
.Y(n_2255)
);

AOI22xp33_ASAP7_75t_SL g2256 ( 
.A1(n_1959),
.A2(n_1953),
.B1(n_1942),
.B2(n_1931),
.Y(n_2256)
);

INVx4_ASAP7_75t_L g2257 ( 
.A(n_1938),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_2169),
.Y(n_2258)
);

AOI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_2087),
.A2(n_2171),
.B1(n_2112),
.B2(n_2180),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2085),
.B(n_2041),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2232),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_L g2262 ( 
.A(n_2096),
.B(n_2072),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2143),
.B(n_2045),
.Y(n_2263)
);

BUFx3_ASAP7_75t_L g2264 ( 
.A(n_2094),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2097),
.B(n_1876),
.Y(n_2265)
);

AOI22xp33_ASAP7_75t_L g2266 ( 
.A1(n_2171),
.A2(n_2006),
.B1(n_1959),
.B2(n_2018),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2086),
.Y(n_2267)
);

BUFx2_ASAP7_75t_L g2268 ( 
.A(n_2257),
.Y(n_2268)
);

HB1xp67_ASAP7_75t_L g2269 ( 
.A(n_2239),
.Y(n_2269)
);

INVxp67_ASAP7_75t_L g2270 ( 
.A(n_2188),
.Y(n_2270)
);

AND2x4_ASAP7_75t_L g2271 ( 
.A(n_2084),
.B(n_2045),
.Y(n_2271)
);

BUFx2_ASAP7_75t_L g2272 ( 
.A(n_2257),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2088),
.Y(n_2273)
);

AND2x4_ASAP7_75t_L g2274 ( 
.A(n_2084),
.B(n_2044),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2110),
.B(n_1876),
.Y(n_2275)
);

HB1xp67_ASAP7_75t_L g2276 ( 
.A(n_2239),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2149),
.B(n_1877),
.Y(n_2277)
);

BUFx2_ASAP7_75t_L g2278 ( 
.A(n_2218),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_2167),
.B(n_1833),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2091),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2114),
.B(n_2009),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2128),
.B(n_2024),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2153),
.B(n_2036),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2153),
.B(n_2036),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2092),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2098),
.Y(n_2286)
);

AND2x4_ASAP7_75t_SL g2287 ( 
.A(n_2179),
.B(n_1948),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2099),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2089),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2100),
.Y(n_2290)
);

INVx2_ASAP7_75t_SL g2291 ( 
.A(n_2242),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2189),
.B(n_2024),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2154),
.B(n_1877),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2101),
.Y(n_2294)
);

AOI22xp33_ASAP7_75t_L g2295 ( 
.A1(n_2155),
.A2(n_1959),
.B1(n_2007),
.B2(n_1931),
.Y(n_2295)
);

INVx2_ASAP7_75t_SL g2296 ( 
.A(n_2242),
.Y(n_2296)
);

BUFx3_ASAP7_75t_L g2297 ( 
.A(n_2094),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2083),
.B(n_1878),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2213),
.B(n_2032),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_2083),
.B(n_2192),
.Y(n_2300)
);

BUFx3_ASAP7_75t_L g2301 ( 
.A(n_2121),
.Y(n_2301)
);

HB1xp67_ASAP7_75t_L g2302 ( 
.A(n_2159),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2102),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2105),
.Y(n_2304)
);

AOI22xp33_ASAP7_75t_L g2305 ( 
.A1(n_2155),
.A2(n_2007),
.B1(n_1931),
.B2(n_1942),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2132),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2224),
.B(n_2032),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2109),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2179),
.B(n_1878),
.Y(n_2309)
);

OR2x2_ASAP7_75t_L g2310 ( 
.A(n_2165),
.B(n_1896),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2231),
.B(n_2046),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2111),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2113),
.Y(n_2313)
);

BUFx3_ASAP7_75t_L g2314 ( 
.A(n_2121),
.Y(n_2314)
);

OR2x2_ASAP7_75t_L g2315 ( 
.A(n_2170),
.B(n_1896),
.Y(n_2315)
);

BUFx3_ASAP7_75t_L g2316 ( 
.A(n_2095),
.Y(n_2316)
);

BUFx2_ASAP7_75t_L g2317 ( 
.A(n_2218),
.Y(n_2317)
);

AOI22xp33_ASAP7_75t_L g2318 ( 
.A1(n_2138),
.A2(n_2007),
.B1(n_1942),
.B2(n_1991),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2115),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2116),
.Y(n_2320)
);

AOI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_2138),
.A2(n_1991),
.B1(n_2043),
.B2(n_1953),
.Y(n_2321)
);

AOI22xp33_ASAP7_75t_L g2322 ( 
.A1(n_2157),
.A2(n_1953),
.B1(n_1999),
.B2(n_2021),
.Y(n_2322)
);

AOI22xp33_ASAP7_75t_SL g2323 ( 
.A1(n_2129),
.A2(n_2029),
.B1(n_1866),
.B2(n_1944),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2117),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2238),
.B(n_2046),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2182),
.B(n_2194),
.Y(n_2326)
);

OAI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_2157),
.A2(n_2027),
.B1(n_1966),
.B2(n_2002),
.Y(n_2327)
);

AND2x2_ASAP7_75t_SL g2328 ( 
.A(n_2129),
.B(n_2044),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2182),
.B(n_1849),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2144),
.B(n_1849),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2227),
.B(n_1949),
.Y(n_2331)
);

INVx5_ASAP7_75t_L g2332 ( 
.A(n_2248),
.Y(n_2332)
);

OR2x2_ASAP7_75t_L g2333 ( 
.A(n_2173),
.B(n_2040),
.Y(n_2333)
);

HB1xp67_ASAP7_75t_L g2334 ( 
.A(n_2104),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2118),
.Y(n_2335)
);

INVx4_ASAP7_75t_L g2336 ( 
.A(n_2084),
.Y(n_2336)
);

OR2x2_ASAP7_75t_L g2337 ( 
.A(n_2177),
.B(n_2090),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2119),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2080),
.B(n_1889),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2125),
.Y(n_2340)
);

BUFx2_ASAP7_75t_L g2341 ( 
.A(n_2145),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2126),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2161),
.B(n_1999),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2127),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2080),
.B(n_1889),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2130),
.Y(n_2346)
);

OR2x2_ASAP7_75t_L g2347 ( 
.A(n_2252),
.B(n_2040),
.Y(n_2347)
);

AOI22xp33_ASAP7_75t_L g2348 ( 
.A1(n_2180),
.A2(n_1978),
.B1(n_2004),
.B2(n_1929),
.Y(n_2348)
);

BUFx2_ASAP7_75t_L g2349 ( 
.A(n_2145),
.Y(n_2349)
);

AOI22xp33_ASAP7_75t_L g2350 ( 
.A1(n_2210),
.A2(n_1929),
.B1(n_1962),
.B2(n_1964),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2240),
.B(n_2035),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2104),
.B(n_2033),
.Y(n_2352)
);

AOI22xp33_ASAP7_75t_L g2353 ( 
.A1(n_2210),
.A2(n_1962),
.B1(n_1964),
.B2(n_1918),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2131),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2135),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2137),
.Y(n_2356)
);

HB1xp67_ASAP7_75t_L g2357 ( 
.A(n_2107),
.Y(n_2357)
);

OAI21xp5_ASAP7_75t_SL g2358 ( 
.A1(n_2243),
.A2(n_1966),
.B(n_2002),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2139),
.Y(n_2359)
);

HB1xp67_ASAP7_75t_L g2360 ( 
.A(n_2107),
.Y(n_2360)
);

BUFx2_ASAP7_75t_L g2361 ( 
.A(n_2225),
.Y(n_2361)
);

AND2x4_ASAP7_75t_L g2362 ( 
.A(n_2241),
.B(n_1933),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2140),
.B(n_2178),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2193),
.Y(n_2364)
);

BUFx3_ASAP7_75t_L g2365 ( 
.A(n_2103),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2185),
.Y(n_2366)
);

HB1xp67_ASAP7_75t_L g2367 ( 
.A(n_2133),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2142),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2146),
.Y(n_2369)
);

OR2x2_ASAP7_75t_L g2370 ( 
.A(n_2220),
.B(n_2221),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2148),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2244),
.B(n_1887),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2201),
.B(n_2022),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2081),
.B(n_2022),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2093),
.B(n_1930),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2152),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2122),
.B(n_2250),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2134),
.B(n_1930),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_2134),
.B(n_2228),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2183),
.B(n_1968),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2245),
.B(n_1852),
.Y(n_2381)
);

INVx2_ASAP7_75t_SL g2382 ( 
.A(n_2242),
.Y(n_2382)
);

HB1xp67_ASAP7_75t_L g2383 ( 
.A(n_2181),
.Y(n_2383)
);

INVxp67_ASAP7_75t_L g2384 ( 
.A(n_2136),
.Y(n_2384)
);

OR2x2_ASAP7_75t_L g2385 ( 
.A(n_2184),
.B(n_2011),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2186),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2187),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_L g2388 ( 
.A(n_2251),
.B(n_1879),
.Y(n_2388)
);

OAI21xp33_ASAP7_75t_L g2389 ( 
.A1(n_2211),
.A2(n_1961),
.B(n_1986),
.Y(n_2389)
);

OR2x2_ASAP7_75t_L g2390 ( 
.A(n_2184),
.B(n_2011),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2233),
.B(n_1862),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2267),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2261),
.Y(n_2393)
);

OR2x2_ASAP7_75t_L g2394 ( 
.A(n_2270),
.B(n_2150),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_SL g2395 ( 
.A(n_2268),
.B(n_2272),
.Y(n_2395)
);

BUFx3_ASAP7_75t_L g2396 ( 
.A(n_2264),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2263),
.B(n_2233),
.Y(n_2397)
);

INVx3_ASAP7_75t_L g2398 ( 
.A(n_2271),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2261),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_2263),
.B(n_2168),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2273),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2280),
.Y(n_2402)
);

OR2x2_ASAP7_75t_L g2403 ( 
.A(n_2361),
.B(n_2150),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2285),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2286),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2352),
.B(n_2123),
.Y(n_2406)
);

OAI222xp33_ASAP7_75t_L g2407 ( 
.A1(n_2259),
.A2(n_2211),
.B1(n_2136),
.B2(n_2124),
.C1(n_2120),
.C2(n_2106),
.Y(n_2407)
);

OR2x2_ASAP7_75t_L g2408 ( 
.A(n_2282),
.B(n_2162),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2308),
.B(n_2245),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2312),
.B(n_2202),
.Y(n_2410)
);

BUFx2_ASAP7_75t_L g2411 ( 
.A(n_2278),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2288),
.Y(n_2412)
);

OR2x2_ASAP7_75t_L g2413 ( 
.A(n_2299),
.B(n_2162),
.Y(n_2413)
);

AOI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_2262),
.A2(n_2377),
.B1(n_2202),
.B2(n_2327),
.Y(n_2414)
);

HB1xp67_ASAP7_75t_L g2415 ( 
.A(n_2269),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2290),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2294),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2303),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2352),
.B(n_2123),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2300),
.B(n_2158),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2304),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2391),
.B(n_2256),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2306),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2313),
.Y(n_2424)
);

INVx1_ASAP7_75t_SL g2425 ( 
.A(n_2289),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2319),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2320),
.B(n_2254),
.Y(n_2427)
);

OR2x2_ASAP7_75t_L g2428 ( 
.A(n_2337),
.B(n_2172),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2324),
.B(n_2196),
.Y(n_2429)
);

BUFx2_ASAP7_75t_L g2430 ( 
.A(n_2317),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2335),
.Y(n_2431)
);

CKINVDCx16_ASAP7_75t_R g2432 ( 
.A(n_2264),
.Y(n_2432)
);

BUFx3_ASAP7_75t_L g2433 ( 
.A(n_2297),
.Y(n_2433)
);

INVxp67_ASAP7_75t_SL g2434 ( 
.A(n_2269),
.Y(n_2434)
);

AOI22xp33_ASAP7_75t_L g2435 ( 
.A1(n_2262),
.A2(n_2236),
.B1(n_2197),
.B2(n_1962),
.Y(n_2435)
);

OAI22xp5_ASAP7_75t_L g2436 ( 
.A1(n_2323),
.A2(n_2120),
.B1(n_2124),
.B2(n_2106),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2338),
.B(n_2199),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2265),
.B(n_2174),
.Y(n_2438)
);

INVx4_ASAP7_75t_R g2439 ( 
.A(n_2297),
.Y(n_2439)
);

HB1xp67_ASAP7_75t_L g2440 ( 
.A(n_2276),
.Y(n_2440)
);

INVxp67_ASAP7_75t_L g2441 ( 
.A(n_2365),
.Y(n_2441)
);

OR2x2_ASAP7_75t_L g2442 ( 
.A(n_2370),
.B(n_2151),
.Y(n_2442)
);

OR2x2_ASAP7_75t_L g2443 ( 
.A(n_2260),
.B(n_2249),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2340),
.B(n_2342),
.Y(n_2444)
);

INVx2_ASAP7_75t_SL g2445 ( 
.A(n_2276),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2391),
.B(n_2372),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2344),
.B(n_2200),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2372),
.B(n_2256),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2283),
.B(n_2284),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2346),
.B(n_2203),
.Y(n_2450)
);

OR2x2_ASAP7_75t_L g2451 ( 
.A(n_2292),
.B(n_2249),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2283),
.B(n_2206),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2284),
.B(n_2206),
.Y(n_2453)
);

AOI22xp33_ASAP7_75t_L g2454 ( 
.A1(n_2348),
.A2(n_2236),
.B1(n_2247),
.B2(n_1918),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2354),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2355),
.Y(n_2456)
);

OR2x2_ASAP7_75t_L g2457 ( 
.A(n_2363),
.B(n_2163),
.Y(n_2457)
);

AND2x4_ASAP7_75t_L g2458 ( 
.A(n_2380),
.B(n_2082),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2356),
.B(n_2230),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2359),
.B(n_2366),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2351),
.B(n_2082),
.Y(n_2461)
);

INVxp67_ASAP7_75t_L g2462 ( 
.A(n_2365),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2364),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2386),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2387),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2368),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2369),
.Y(n_2467)
);

OR2x2_ASAP7_75t_L g2468 ( 
.A(n_2279),
.B(n_2164),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2281),
.B(n_2212),
.Y(n_2469)
);

AND2x2_ASAP7_75t_SL g2470 ( 
.A(n_2328),
.B(n_2336),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2293),
.B(n_2191),
.Y(n_2471)
);

OR2x2_ASAP7_75t_L g2472 ( 
.A(n_2334),
.B(n_2237),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2266),
.B(n_2215),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2371),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2277),
.B(n_2166),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2376),
.Y(n_2476)
);

INVxp67_ASAP7_75t_L g2477 ( 
.A(n_2301),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2333),
.Y(n_2478)
);

AOI22xp5_ASAP7_75t_L g2479 ( 
.A1(n_2358),
.A2(n_2141),
.B1(n_2205),
.B2(n_2255),
.Y(n_2479)
);

OAI21xp33_ASAP7_75t_L g2480 ( 
.A1(n_2266),
.A2(n_2156),
.B(n_2214),
.Y(n_2480)
);

INVx3_ASAP7_75t_L g2481 ( 
.A(n_2271),
.Y(n_2481)
);

INVxp67_ASAP7_75t_L g2482 ( 
.A(n_2301),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2334),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2379),
.B(n_2166),
.Y(n_2484)
);

BUFx2_ASAP7_75t_SL g2485 ( 
.A(n_2396),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2446),
.B(n_2311),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2464),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2446),
.B(n_2325),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2409),
.B(n_2307),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2397),
.B(n_2326),
.Y(n_2490)
);

OR2x2_ASAP7_75t_L g2491 ( 
.A(n_2408),
.B(n_2403),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2478),
.B(n_2381),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2465),
.Y(n_2493)
);

OAI221xp5_ASAP7_75t_SL g2494 ( 
.A1(n_2414),
.A2(n_2348),
.B1(n_2321),
.B2(n_2322),
.C(n_2353),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2422),
.B(n_2325),
.Y(n_2495)
);

AND2x4_ASAP7_75t_L g2496 ( 
.A(n_2398),
.B(n_2271),
.Y(n_2496)
);

CKINVDCx5p33_ASAP7_75t_R g2497 ( 
.A(n_2432),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2393),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2392),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2401),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2422),
.B(n_2347),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2402),
.Y(n_2502)
);

AND2x2_ASAP7_75t_L g2503 ( 
.A(n_2406),
.B(n_2362),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2393),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2399),
.Y(n_2505)
);

OR2x2_ASAP7_75t_L g2506 ( 
.A(n_2442),
.B(n_2357),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2404),
.Y(n_2507)
);

AND2x4_ASAP7_75t_L g2508 ( 
.A(n_2398),
.B(n_2362),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2405),
.Y(n_2509)
);

BUFx2_ASAP7_75t_L g2510 ( 
.A(n_2396),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2397),
.B(n_2328),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2406),
.B(n_2419),
.Y(n_2512)
);

AND2x2_ASAP7_75t_L g2513 ( 
.A(n_2420),
.B(n_2357),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_2395),
.B(n_2316),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2419),
.B(n_2362),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2412),
.Y(n_2516)
);

AND2x4_ASAP7_75t_L g2517 ( 
.A(n_2398),
.B(n_2274),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2416),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2449),
.B(n_2322),
.Y(n_2519)
);

INVx6_ASAP7_75t_L g2520 ( 
.A(n_2433),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2417),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2418),
.Y(n_2522)
);

INVxp67_ASAP7_75t_L g2523 ( 
.A(n_2395),
.Y(n_2523)
);

NOR3xp33_ASAP7_75t_L g2524 ( 
.A(n_2480),
.B(n_2388),
.C(n_2226),
.Y(n_2524)
);

OR2x2_ASAP7_75t_L g2525 ( 
.A(n_2413),
.B(n_2360),
.Y(n_2525)
);

OR2x2_ASAP7_75t_L g2526 ( 
.A(n_2394),
.B(n_2360),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2448),
.B(n_2302),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2421),
.Y(n_2528)
);

AND2x4_ASAP7_75t_L g2529 ( 
.A(n_2481),
.B(n_2274),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2449),
.B(n_2343),
.Y(n_2530)
);

OR2x2_ASAP7_75t_L g2531 ( 
.A(n_2445),
.B(n_2434),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2423),
.B(n_2367),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2424),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2426),
.Y(n_2534)
);

NOR3xp33_ASAP7_75t_L g2535 ( 
.A(n_2407),
.B(n_2388),
.C(n_2248),
.Y(n_2535)
);

OAI21xp33_ASAP7_75t_L g2536 ( 
.A1(n_2435),
.A2(n_2321),
.B(n_2389),
.Y(n_2536)
);

AND2x2_ASAP7_75t_L g2537 ( 
.A(n_2448),
.B(n_2302),
.Y(n_2537)
);

OR2x2_ASAP7_75t_L g2538 ( 
.A(n_2445),
.B(n_2367),
.Y(n_2538)
);

AND2x4_ASAP7_75t_L g2539 ( 
.A(n_2481),
.B(n_2274),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2431),
.B(n_2305),
.Y(n_2540)
);

OR2x2_ASAP7_75t_L g2541 ( 
.A(n_2415),
.B(n_2383),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2498),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2498),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2487),
.Y(n_2544)
);

AND2x4_ASAP7_75t_SL g2545 ( 
.A(n_2496),
.B(n_2336),
.Y(n_2545)
);

INVxp67_ASAP7_75t_L g2546 ( 
.A(n_2485),
.Y(n_2546)
);

NAND3xp33_ASAP7_75t_L g2547 ( 
.A(n_2524),
.B(n_2536),
.C(n_2523),
.Y(n_2547)
);

INVxp67_ASAP7_75t_L g2548 ( 
.A(n_2510),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2512),
.B(n_2486),
.Y(n_2549)
);

INVx1_ASAP7_75t_SL g2550 ( 
.A(n_2497),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2504),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2512),
.B(n_2452),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2486),
.B(n_2452),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2495),
.B(n_2410),
.Y(n_2554)
);

OR2x2_ASAP7_75t_L g2555 ( 
.A(n_2491),
.B(n_2415),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2493),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2495),
.B(n_2483),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2488),
.B(n_2453),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2499),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2504),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_2488),
.B(n_2453),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2500),
.Y(n_2562)
);

INVxp67_ASAP7_75t_SL g2563 ( 
.A(n_2531),
.Y(n_2563)
);

NAND2x1p5_ASAP7_75t_L g2564 ( 
.A(n_2514),
.B(n_2470),
.Y(n_2564)
);

OR2x2_ASAP7_75t_L g2565 ( 
.A(n_2530),
.B(n_2440),
.Y(n_2565)
);

HB1xp67_ASAP7_75t_L g2566 ( 
.A(n_2541),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2501),
.B(n_2400),
.Y(n_2567)
);

OR2x2_ASAP7_75t_L g2568 ( 
.A(n_2525),
.B(n_2440),
.Y(n_2568)
);

NAND2x1p5_ASAP7_75t_L g2569 ( 
.A(n_2514),
.B(n_2470),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2501),
.B(n_2400),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2502),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2507),
.Y(n_2572)
);

AND2x4_ASAP7_75t_L g2573 ( 
.A(n_2508),
.B(n_2481),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2505),
.Y(n_2574)
);

AND2x4_ASAP7_75t_L g2575 ( 
.A(n_2508),
.B(n_2458),
.Y(n_2575)
);

OR2x2_ASAP7_75t_L g2576 ( 
.A(n_2506),
.B(n_2461),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2509),
.Y(n_2577)
);

OR2x6_ASAP7_75t_L g2578 ( 
.A(n_2520),
.B(n_2336),
.Y(n_2578)
);

NAND2x2_ASAP7_75t_L g2579 ( 
.A(n_2535),
.B(n_2314),
.Y(n_2579)
);

NAND2x1p5_ASAP7_75t_L g2580 ( 
.A(n_2496),
.B(n_2332),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2516),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2518),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2521),
.Y(n_2583)
);

AND2x4_ASAP7_75t_SL g2584 ( 
.A(n_2496),
.B(n_2475),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2503),
.B(n_2461),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2565),
.Y(n_2586)
);

OR2x2_ASAP7_75t_L g2587 ( 
.A(n_2565),
.B(n_2527),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2566),
.B(n_2527),
.Y(n_2588)
);

AOI22xp5_ASAP7_75t_L g2589 ( 
.A1(n_2547),
.A2(n_2524),
.B1(n_2535),
.B2(n_2435),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2555),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2555),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2581),
.Y(n_2592)
);

INVxp67_ASAP7_75t_L g2593 ( 
.A(n_2563),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2581),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2549),
.B(n_2554),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2542),
.Y(n_2596)
);

OR2x2_ASAP7_75t_L g2597 ( 
.A(n_2576),
.B(n_2537),
.Y(n_2597)
);

INVx1_ASAP7_75t_SL g2598 ( 
.A(n_2584),
.Y(n_2598)
);

NAND3xp33_ASAP7_75t_L g2599 ( 
.A(n_2546),
.B(n_2494),
.C(n_2332),
.Y(n_2599)
);

O2A1O1Ixp33_ASAP7_75t_SL g2600 ( 
.A1(n_2550),
.A2(n_2384),
.B(n_2425),
.C(n_2441),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2544),
.B(n_2537),
.Y(n_2601)
);

AND2x4_ASAP7_75t_L g2602 ( 
.A(n_2584),
.B(n_2508),
.Y(n_2602)
);

AOI32xp33_ASAP7_75t_L g2603 ( 
.A1(n_2549),
.A2(n_2430),
.A3(n_2411),
.B1(n_2497),
.B2(n_2436),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2568),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2552),
.B(n_2503),
.Y(n_2605)
);

AND2x4_ASAP7_75t_L g2606 ( 
.A(n_2545),
.B(n_2517),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2568),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2552),
.B(n_2515),
.Y(n_2608)
);

OAI33xp33_ASAP7_75t_L g2609 ( 
.A1(n_2548),
.A2(n_2428),
.A3(n_2492),
.B1(n_2519),
.B2(n_2457),
.B3(n_2489),
.Y(n_2609)
);

O2A1O1Ixp33_ASAP7_75t_L g2610 ( 
.A1(n_2564),
.A2(n_2462),
.B(n_2160),
.C(n_2459),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2576),
.Y(n_2611)
);

OR2x2_ASAP7_75t_L g2612 ( 
.A(n_2557),
.B(n_2526),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2542),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2556),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2559),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2562),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2571),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2543),
.Y(n_2618)
);

INVx3_ASAP7_75t_L g2619 ( 
.A(n_2580),
.Y(n_2619)
);

OAI22xp5_ASAP7_75t_L g2620 ( 
.A1(n_2579),
.A2(n_2520),
.B1(n_2482),
.B2(n_2477),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2572),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_SL g2622 ( 
.A(n_2580),
.B(n_2433),
.Y(n_2622)
);

CKINVDCx16_ASAP7_75t_R g2623 ( 
.A(n_2578),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2577),
.B(n_2522),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2582),
.Y(n_2625)
);

OR2x2_ASAP7_75t_L g2626 ( 
.A(n_2567),
.B(n_2513),
.Y(n_2626)
);

INVxp67_ASAP7_75t_SL g2627 ( 
.A(n_2580),
.Y(n_2627)
);

OAI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2598),
.A2(n_2623),
.B1(n_2579),
.B2(n_2627),
.Y(n_2628)
);

OAI21xp5_ASAP7_75t_L g2629 ( 
.A1(n_2589),
.A2(n_2569),
.B(n_2564),
.Y(n_2629)
);

AOI31xp33_ASAP7_75t_L g2630 ( 
.A1(n_2600),
.A2(n_2564),
.A3(n_2569),
.B(n_2258),
.Y(n_2630)
);

OAI21xp5_ASAP7_75t_L g2631 ( 
.A1(n_2599),
.A2(n_2569),
.B(n_2332),
.Y(n_2631)
);

AOI22xp5_ASAP7_75t_L g2632 ( 
.A1(n_2599),
.A2(n_2573),
.B1(n_2575),
.B2(n_2490),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2592),
.Y(n_2633)
);

OAI211xp5_ASAP7_75t_L g2634 ( 
.A1(n_2603),
.A2(n_2479),
.B(n_2332),
.C(n_2454),
.Y(n_2634)
);

NAND3xp33_ASAP7_75t_SL g2635 ( 
.A(n_2610),
.B(n_2258),
.C(n_2198),
.Y(n_2635)
);

INVx1_ASAP7_75t_SL g2636 ( 
.A(n_2598),
.Y(n_2636)
);

OAI22xp33_ASAP7_75t_L g2637 ( 
.A1(n_2622),
.A2(n_2578),
.B1(n_2520),
.B2(n_2573),
.Y(n_2637)
);

AOI21xp5_ASAP7_75t_L g2638 ( 
.A1(n_2622),
.A2(n_2578),
.B(n_2545),
.Y(n_2638)
);

OAI22xp5_ASAP7_75t_L g2639 ( 
.A1(n_2619),
.A2(n_2578),
.B1(n_2575),
.B2(n_2573),
.Y(n_2639)
);

AOI22xp33_ASAP7_75t_L g2640 ( 
.A1(n_2609),
.A2(n_2575),
.B1(n_2511),
.B2(n_2515),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2594),
.Y(n_2641)
);

INVxp67_ASAP7_75t_L g2642 ( 
.A(n_2624),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2586),
.B(n_2590),
.Y(n_2643)
);

OAI21xp5_ASAP7_75t_L g2644 ( 
.A1(n_2593),
.A2(n_2454),
.B(n_2318),
.Y(n_2644)
);

INVxp33_ASAP7_75t_L g2645 ( 
.A(n_2606),
.Y(n_2645)
);

AOI322xp5_ASAP7_75t_L g2646 ( 
.A1(n_2611),
.A2(n_2561),
.A3(n_2553),
.B1(n_2558),
.B2(n_2567),
.C1(n_2570),
.C2(n_2585),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2624),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2596),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2619),
.A2(n_2570),
.B1(n_2558),
.B2(n_2561),
.Y(n_2649)
);

OAI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2620),
.A2(n_2538),
.B1(n_2472),
.B2(n_2169),
.Y(n_2650)
);

AOI21xp5_ASAP7_75t_L g2651 ( 
.A1(n_2620),
.A2(n_2529),
.B(n_2517),
.Y(n_2651)
);

AOI21xp33_ASAP7_75t_L g2652 ( 
.A1(n_2614),
.A2(n_2540),
.B(n_2473),
.Y(n_2652)
);

INVxp67_ASAP7_75t_L g2653 ( 
.A(n_2615),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2587),
.Y(n_2654)
);

INVxp67_ASAP7_75t_L g2655 ( 
.A(n_2616),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2643),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2642),
.B(n_2647),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2636),
.Y(n_2658)
);

NAND4xp25_ASAP7_75t_L g2659 ( 
.A(n_2629),
.B(n_2353),
.C(n_2350),
.D(n_2318),
.Y(n_2659)
);

AOI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2634),
.A2(n_2607),
.B1(n_2604),
.B2(n_2591),
.Y(n_2660)
);

NOR2x1p5_ASAP7_75t_L g2661 ( 
.A(n_2635),
.B(n_2602),
.Y(n_2661)
);

AOI211xp5_ASAP7_75t_SL g2662 ( 
.A1(n_2630),
.A2(n_2628),
.B(n_2650),
.C(n_2637),
.Y(n_2662)
);

O2A1O1Ixp33_ASAP7_75t_L g2663 ( 
.A1(n_2631),
.A2(n_2621),
.B(n_2625),
.C(n_2617),
.Y(n_2663)
);

OAI211xp5_ASAP7_75t_L g2664 ( 
.A1(n_2638),
.A2(n_2314),
.B(n_2349),
.C(n_2341),
.Y(n_2664)
);

OAI211xp5_ASAP7_75t_SL g2665 ( 
.A1(n_2632),
.A2(n_2601),
.B(n_2350),
.C(n_2588),
.Y(n_2665)
);

AOI21xp5_ASAP7_75t_L g2666 ( 
.A1(n_2645),
.A2(n_2606),
.B(n_2602),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2642),
.B(n_2595),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_SL g2668 ( 
.A1(n_2639),
.A2(n_2517),
.B1(n_2539),
.B2(n_2529),
.Y(n_2668)
);

AOI221x1_ASAP7_75t_L g2669 ( 
.A1(n_2651),
.A2(n_2583),
.B1(n_2601),
.B2(n_2534),
.C(n_2533),
.Y(n_2669)
);

AO22x1_ASAP7_75t_L g2670 ( 
.A1(n_2649),
.A2(n_2439),
.B1(n_2316),
.B2(n_2605),
.Y(n_2670)
);

OAI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2640),
.A2(n_2626),
.B1(n_2597),
.B2(n_2612),
.Y(n_2671)
);

HB1xp67_ASAP7_75t_L g2672 ( 
.A(n_2653),
.Y(n_2672)
);

AOI22xp33_ASAP7_75t_SL g2673 ( 
.A1(n_2644),
.A2(n_2529),
.B1(n_2539),
.B2(n_2484),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2646),
.B(n_2608),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2648),
.Y(n_2675)
);

NOR4xp25_ASAP7_75t_L g2676 ( 
.A(n_2653),
.B(n_2460),
.C(n_2444),
.D(n_2528),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2655),
.B(n_2553),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_SL g2678 ( 
.A(n_2652),
.B(n_2613),
.Y(n_2678)
);

NOR3xp33_ASAP7_75t_L g2679 ( 
.A(n_2633),
.B(n_2195),
.C(n_2237),
.Y(n_2679)
);

OAI211xp5_ASAP7_75t_L g2680 ( 
.A1(n_2654),
.A2(n_1832),
.B(n_2375),
.C(n_2175),
.Y(n_2680)
);

AOI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2641),
.A2(n_2471),
.B1(n_2539),
.B2(n_2585),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2643),
.Y(n_2682)
);

OAI22xp5_ASAP7_75t_SL g2683 ( 
.A1(n_2645),
.A2(n_1879),
.B1(n_2175),
.B2(n_2291),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2636),
.Y(n_2684)
);

AOI21xp5_ASAP7_75t_SL g2685 ( 
.A1(n_2661),
.A2(n_1853),
.B(n_2291),
.Y(n_2685)
);

NAND4xp25_ASAP7_75t_SL g2686 ( 
.A(n_2666),
.B(n_2468),
.C(n_2331),
.D(n_2305),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2658),
.Y(n_2687)
);

O2A1O1Ixp5_ASAP7_75t_L g2688 ( 
.A1(n_2662),
.A2(n_2618),
.B(n_2532),
.C(n_2469),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2656),
.B(n_2682),
.Y(n_2689)
);

NOR2xp33_ASAP7_75t_SL g2690 ( 
.A(n_2683),
.B(n_1895),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2684),
.B(n_2455),
.Y(n_2691)
);

AOI211xp5_ASAP7_75t_L g2692 ( 
.A1(n_2680),
.A2(n_2385),
.B(n_2390),
.C(n_2378),
.Y(n_2692)
);

NOR3x1_ASAP7_75t_L g2693 ( 
.A(n_2680),
.B(n_2382),
.C(n_2296),
.Y(n_2693)
);

AND4x1_ASAP7_75t_L g2694 ( 
.A(n_2666),
.B(n_1897),
.C(n_1853),
.D(n_2374),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2672),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2675),
.Y(n_2696)
);

NOR3xp33_ASAP7_75t_L g2697 ( 
.A(n_2664),
.B(n_2216),
.C(n_2208),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2657),
.Y(n_2698)
);

NOR2xp67_ASAP7_75t_L g2699 ( 
.A(n_2664),
.B(n_2543),
.Y(n_2699)
);

OAI211xp5_ASAP7_75t_SL g2700 ( 
.A1(n_2660),
.A2(n_2295),
.B(n_2437),
.C(n_2429),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2667),
.Y(n_2701)
);

NAND3xp33_ASAP7_75t_L g2702 ( 
.A(n_2669),
.B(n_2295),
.C(n_2222),
.Y(n_2702)
);

NOR3x1_ASAP7_75t_L g2703 ( 
.A(n_2670),
.B(n_2382),
.C(n_2296),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2676),
.B(n_2456),
.Y(n_2704)
);

OA22x2_ASAP7_75t_L g2705 ( 
.A1(n_2671),
.A2(n_2463),
.B1(n_2287),
.B2(n_2209),
.Y(n_2705)
);

A2O1A1Ixp33_ASAP7_75t_L g2706 ( 
.A1(n_2663),
.A2(n_2287),
.B(n_2190),
.C(n_2207),
.Y(n_2706)
);

NOR2x1_ASAP7_75t_L g2707 ( 
.A(n_2685),
.B(n_2665),
.Y(n_2707)
);

INVx2_ASAP7_75t_SL g2708 ( 
.A(n_2687),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2698),
.B(n_2674),
.Y(n_2709)
);

NAND4xp75_ASAP7_75t_L g2710 ( 
.A(n_2688),
.B(n_2678),
.C(n_2681),
.D(n_2677),
.Y(n_2710)
);

NAND4xp75_ASAP7_75t_SL g2711 ( 
.A(n_2694),
.B(n_2668),
.C(n_2673),
.D(n_2659),
.Y(n_2711)
);

NOR2x1_ASAP7_75t_L g2712 ( 
.A(n_2695),
.B(n_2706),
.Y(n_2712)
);

INVx2_ASAP7_75t_SL g2713 ( 
.A(n_2696),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2701),
.B(n_2679),
.Y(n_2714)
);

AND2x4_ASAP7_75t_L g2715 ( 
.A(n_2693),
.B(n_2438),
.Y(n_2715)
);

HB1xp67_ASAP7_75t_L g2716 ( 
.A(n_2689),
.Y(n_2716)
);

NOR3x1_ASAP7_75t_L g2717 ( 
.A(n_2689),
.B(n_1851),
.C(n_2447),
.Y(n_2717)
);

NOR2x1_ASAP7_75t_L g2718 ( 
.A(n_2686),
.B(n_2217),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_SL g2719 ( 
.A(n_2690),
.B(n_1891),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2691),
.Y(n_2720)
);

NOR3xp33_ASAP7_75t_SL g2721 ( 
.A(n_2700),
.B(n_2702),
.C(n_2704),
.Y(n_2721)
);

AOI21xp5_ASAP7_75t_L g2722 ( 
.A1(n_2705),
.A2(n_2450),
.B(n_2427),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_SL g2723 ( 
.A(n_2699),
.B(n_1891),
.Y(n_2723)
);

NOR3x1_ASAP7_75t_L g2724 ( 
.A(n_2705),
.B(n_2246),
.C(n_2253),
.Y(n_2724)
);

NOR3x1_ASAP7_75t_L g2725 ( 
.A(n_2703),
.B(n_1943),
.C(n_2443),
.Y(n_2725)
);

NAND3xp33_ASAP7_75t_L g2726 ( 
.A(n_2716),
.B(n_2692),
.C(n_2697),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2708),
.B(n_2466),
.Y(n_2727)
);

NAND4xp25_ASAP7_75t_L g2728 ( 
.A(n_2709),
.B(n_2190),
.C(n_2207),
.D(n_2204),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_SL g2729 ( 
.A(n_2707),
.B(n_2713),
.Y(n_2729)
);

NOR2x1_ASAP7_75t_L g2730 ( 
.A(n_2711),
.B(n_2217),
.Y(n_2730)
);

NOR2xp33_ASAP7_75t_L g2731 ( 
.A(n_2710),
.B(n_2467),
.Y(n_2731)
);

NAND2x1_ASAP7_75t_L g2732 ( 
.A(n_2712),
.B(n_2204),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_2715),
.B(n_2551),
.Y(n_2733)
);

HB1xp67_ASAP7_75t_L g2734 ( 
.A(n_2720),
.Y(n_2734)
);

AOI21xp5_ASAP7_75t_L g2735 ( 
.A1(n_2719),
.A2(n_2476),
.B(n_2474),
.Y(n_2735)
);

AO22x2_ASAP7_75t_SL g2736 ( 
.A1(n_2724),
.A2(n_2721),
.B1(n_2725),
.B2(n_2714),
.Y(n_2736)
);

CKINVDCx6p67_ASAP7_75t_R g2737 ( 
.A(n_2715),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2722),
.B(n_2717),
.Y(n_2738)
);

NOR3xp33_ASAP7_75t_L g2739 ( 
.A(n_2718),
.B(n_1998),
.C(n_2235),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2723),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2708),
.B(n_2551),
.Y(n_2741)
);

OAI22xp5_ASAP7_75t_L g2742 ( 
.A1(n_2737),
.A2(n_2451),
.B1(n_2574),
.B2(n_2560),
.Y(n_2742)
);

XNOR2xp5_ASAP7_75t_L g2743 ( 
.A(n_2736),
.B(n_2339),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2734),
.Y(n_2744)
);

NAND4xp75_ASAP7_75t_L g2745 ( 
.A(n_2730),
.B(n_2234),
.C(n_2345),
.D(n_2015),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2733),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2731),
.B(n_2560),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2727),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2741),
.Y(n_2749)
);

NAND4xp75_ASAP7_75t_L g2750 ( 
.A(n_2729),
.B(n_1997),
.C(n_2229),
.D(n_2219),
.Y(n_2750)
);

NOR2xp67_ASAP7_75t_L g2751 ( 
.A(n_2726),
.B(n_2223),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2726),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2735),
.B(n_2574),
.Y(n_2753)
);

CKINVDCx5p33_ASAP7_75t_R g2754 ( 
.A(n_2752),
.Y(n_2754)
);

OAI22x1_ASAP7_75t_L g2755 ( 
.A1(n_2743),
.A2(n_2738),
.B1(n_2740),
.B2(n_2732),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2744),
.Y(n_2756)
);

AND2x4_ASAP7_75t_L g2757 ( 
.A(n_2746),
.B(n_2739),
.Y(n_2757)
);

AOI22xp5_ASAP7_75t_L g2758 ( 
.A1(n_2745),
.A2(n_2728),
.B1(n_1906),
.B2(n_2330),
.Y(n_2758)
);

NOR2x1_ASAP7_75t_L g2759 ( 
.A(n_2749),
.B(n_2176),
.Y(n_2759)
);

OAI22x1_ASAP7_75t_L g2760 ( 
.A1(n_2748),
.A2(n_1906),
.B1(n_1997),
.B2(n_1970),
.Y(n_2760)
);

HB1xp67_ASAP7_75t_L g2761 ( 
.A(n_2751),
.Y(n_2761)
);

NAND2xp33_ASAP7_75t_R g2762 ( 
.A(n_2747),
.B(n_2108),
.Y(n_2762)
);

NOR2xp33_ASAP7_75t_L g2763 ( 
.A(n_2742),
.B(n_2751),
.Y(n_2763)
);

XNOR2x1_ASAP7_75t_L g2764 ( 
.A(n_2750),
.B(n_2753),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2744),
.Y(n_2765)
);

BUFx3_ASAP7_75t_L g2766 ( 
.A(n_2744),
.Y(n_2766)
);

AOI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2754),
.A2(n_2329),
.B1(n_2373),
.B2(n_2309),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2766),
.Y(n_2768)
);

AOI22xp5_ASAP7_75t_L g2769 ( 
.A1(n_2755),
.A2(n_1891),
.B1(n_2298),
.B2(n_2275),
.Y(n_2769)
);

OAI22x1_ASAP7_75t_L g2770 ( 
.A1(n_2756),
.A2(n_1997),
.B1(n_1970),
.B2(n_2147),
.Y(n_2770)
);

XNOR2xp5_ASAP7_75t_L g2771 ( 
.A(n_2758),
.B(n_1968),
.Y(n_2771)
);

XNOR2x1_ASAP7_75t_L g2772 ( 
.A(n_2765),
.B(n_1859),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_SL g2773 ( 
.A(n_2757),
.B(n_1891),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2768),
.B(n_2763),
.Y(n_2774)
);

XNOR2x1_ASAP7_75t_L g2775 ( 
.A(n_2772),
.B(n_2764),
.Y(n_2775)
);

XNOR2x1_ASAP7_75t_L g2776 ( 
.A(n_2771),
.B(n_2759),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2770),
.Y(n_2777)
);

OA21x2_ASAP7_75t_L g2778 ( 
.A1(n_2773),
.A2(n_2761),
.B(n_2757),
.Y(n_2778)
);

AOI21x1_ASAP7_75t_L g2779 ( 
.A1(n_2774),
.A2(n_2769),
.B(n_2760),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2778),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2778),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2777),
.Y(n_2782)
);

AOI21xp5_ASAP7_75t_L g2783 ( 
.A1(n_2775),
.A2(n_2767),
.B(n_2762),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2780),
.Y(n_2784)
);

INVx3_ASAP7_75t_L g2785 ( 
.A(n_2782),
.Y(n_2785)
);

AOI22x1_ASAP7_75t_L g2786 ( 
.A1(n_2781),
.A2(n_2783),
.B1(n_2776),
.B2(n_2779),
.Y(n_2786)
);

AO21x1_ASAP7_75t_SL g2787 ( 
.A1(n_2784),
.A2(n_2315),
.B(n_2310),
.Y(n_2787)
);

NOR2xp33_ASAP7_75t_L g2788 ( 
.A(n_2787),
.B(n_2785),
.Y(n_2788)
);

OR2x6_ASAP7_75t_L g2789 ( 
.A(n_2788),
.B(n_2785),
.Y(n_2789)
);

AOI211xp5_ASAP7_75t_L g2790 ( 
.A1(n_2789),
.A2(n_2785),
.B(n_2786),
.C(n_2176),
.Y(n_2790)
);


endmodule