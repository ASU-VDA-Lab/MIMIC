module fake_jpeg_31958_n_314 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_22),
.B(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_44),
.B(n_16),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_21),
.A2(n_0),
.B(n_1),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_61),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_51),
.B(n_66),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_53),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

CKINVDCx9p33_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

INVx5_ASAP7_75t_SL g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_58),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_16),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_65),
.Y(n_73)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_24),
.B(n_3),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_69),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_27),
.Y(n_69)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_43),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_36),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_78),
.B(n_85),
.C(n_102),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_27),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_19),
.B1(n_35),
.B2(n_31),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_88),
.B1(n_103),
.B2(n_64),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_29),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_35),
.B1(n_31),
.B2(n_19),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_29),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_47),
.Y(n_97)
);

CKINVDCx12_ASAP7_75t_R g98 ( 
.A(n_47),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g148 ( 
.A(n_98),
.Y(n_148)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_44),
.B(n_32),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_57),
.A2(n_35),
.B1(n_19),
.B2(n_42),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_32),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_110),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_53),
.A2(n_25),
.B(n_39),
.C(n_38),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_149)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

CKINVDCx12_ASAP7_75t_R g111 ( 
.A(n_50),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_111),
.Y(n_144)
);

BUFx10_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_113),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_37),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_138),
.C(n_145),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_37),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_121),
.Y(n_151)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_117),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_74),
.B(n_38),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_131),
.B1(n_88),
.B2(n_105),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_129),
.Y(n_154)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_99),
.B1(n_109),
.B2(n_59),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_136),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_81),
.A2(n_41),
.B1(n_42),
.B2(n_45),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_141),
.B(n_147),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_73),
.B(n_36),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_82),
.B(n_26),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_96),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_113),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_72),
.Y(n_140)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_81),
.A2(n_41),
.B1(n_40),
.B2(n_68),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_26),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_93),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_108),
.A2(n_50),
.B(n_68),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_76),
.B(n_39),
.C(n_68),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_70),
.B(n_8),
.C(n_9),
.Y(n_158)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_153),
.A2(n_177),
.B1(n_179),
.B2(n_181),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_109),
.B1(n_99),
.B2(n_105),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_156),
.A2(n_173),
.B1(n_169),
.B2(n_164),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_158),
.A2(n_118),
.B(n_11),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_161),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_79),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_163),
.B(n_144),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_87),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_165),
.Y(n_200)
);

BUFx4f_ASAP7_75t_SL g166 ( 
.A(n_137),
.Y(n_166)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_86),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_184),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_122),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_182),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_72),
.B1(n_91),
.B2(n_86),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_131),
.A2(n_91),
.B1(n_95),
.B2(n_87),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_95),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_178),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_93),
.B1(n_8),
.B2(n_9),
.Y(n_179)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_138),
.B(n_7),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_146),
.C(n_117),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_115),
.B(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_114),
.B(n_124),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_153),
.A2(n_149),
.B1(n_140),
.B2(n_125),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_150),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_186),
.A2(n_191),
.B(n_196),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_194),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_135),
.B1(n_130),
.B2(n_133),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_190),
.A2(n_195),
.B1(n_204),
.B2(n_205),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_125),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_142),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_159),
.A2(n_118),
.B(n_144),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_206),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_174),
.B(n_137),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_211),
.C(n_179),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_154),
.B(n_181),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_203),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_156),
.A2(n_168),
.B1(n_161),
.B2(n_184),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_155),
.A2(n_128),
.B1(n_127),
.B2(n_132),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_167),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_170),
.C(n_157),
.Y(n_234)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_148),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_213),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_151),
.B(n_148),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_180),
.Y(n_217)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

XOR2x1_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_158),
.Y(n_219)
);

AOI21x1_ASAP7_75t_L g255 ( 
.A1(n_219),
.A2(n_238),
.B(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_183),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_223),
.B(n_231),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_208),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_232),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_159),
.C(n_175),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_234),
.C(n_209),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_166),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_229),
.B(n_237),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_190),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_175),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g235 ( 
.A1(n_196),
.A2(n_177),
.B(n_169),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_185),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_199),
.A2(n_166),
.B(n_170),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_236),
.A2(n_164),
.B(n_205),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_200),
.B(n_157),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_202),
.A2(n_167),
.B(n_164),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_245),
.C(n_246),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_220),
.B(n_224),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_248),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_255),
.B(n_219),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_191),
.C(n_201),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_192),
.C(n_197),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_237),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_221),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_249),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_188),
.B1(n_207),
.B2(n_197),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_250),
.A2(n_258),
.B1(n_230),
.B2(n_235),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_211),
.C(n_186),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_226),
.C(n_230),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_253),
.B(n_236),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_216),
.A2(n_204),
.B1(n_195),
.B2(n_207),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_257),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_216),
.A2(n_188),
.B1(n_186),
.B2(n_206),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_266),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_242),
.Y(n_281)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_217),
.A3(n_235),
.B1(n_208),
.B2(n_227),
.C1(n_232),
.C2(n_223),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_267),
.B(n_268),
.Y(n_277)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_235),
.A3(n_227),
.B1(n_215),
.B2(n_218),
.C1(n_222),
.C2(n_203),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_215),
.B(n_233),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_252),
.B(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_240),
.B(n_233),
.Y(n_273)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_239),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_276),
.C(n_280),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_256),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_256),
.Y(n_280)
);

XNOR2x1_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_273),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_272),
.B(n_270),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_269),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_245),
.C(n_251),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_285),
.B(n_246),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_271),
.B1(n_264),
.B2(n_258),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_286),
.A2(n_294),
.B1(n_295),
.B2(n_210),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_288),
.B(n_291),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_284),
.A2(n_262),
.B1(n_254),
.B2(n_247),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_292),
.B1(n_287),
.B2(n_162),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_265),
.B(n_266),
.Y(n_290)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_285),
.B(n_270),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_293),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_275),
.B(n_265),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g297 ( 
.A1(n_295),
.A2(n_261),
.B(n_274),
.C(n_279),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_297),
.A2(n_298),
.B1(n_300),
.B2(n_152),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_253),
.A3(n_274),
.B1(n_269),
.B2(n_276),
.C1(n_280),
.C2(n_198),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_198),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_289),
.B1(n_302),
.B2(n_299),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_304),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_302),
.B(n_287),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_152),
.C(n_162),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_297),
.C(n_116),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_307),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_306),
.C(n_10),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_312),
.B(n_14),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_10),
.B(n_14),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_309),
.Y(n_314)
);


endmodule