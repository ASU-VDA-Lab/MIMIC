module fake_jpeg_1695_n_575 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_575);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_575;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_13),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g143 ( 
.A(n_58),
.Y(n_143)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_60),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_61),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_63),
.Y(n_175)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_9),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_65),
.B(n_77),
.Y(n_134)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_71),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_73),
.Y(n_174)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_76),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_32),
.B(n_9),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_85),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_80),
.Y(n_187)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_81),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_82),
.Y(n_169)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_20),
.B(n_9),
.Y(n_85)
);

CKINVDCx9p33_ASAP7_75t_R g86 ( 
.A(n_44),
.Y(n_86)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_88),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_8),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_89),
.B(n_91),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_90),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_23),
.B(n_8),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

BUFx8_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_94),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_95),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_55),
.Y(n_96)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_99),
.Y(n_212)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_102),
.Y(n_177)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_52),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_104),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_24),
.B(n_10),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_16),
.Y(n_159)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_114),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_56),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_115),
.B(n_55),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_40),
.A2(n_7),
.B1(n_17),
.B2(n_2),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_43),
.B1(n_38),
.B2(n_48),
.Y(n_168)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_37),
.B(n_7),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_120),
.B(n_124),
.Y(n_211)
);

BUFx24_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

INVx6_ASAP7_75t_SL g154 ( 
.A(n_121),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

BUFx2_ASAP7_75t_R g126 ( 
.A(n_123),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_37),
.B(n_11),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_94),
.A2(n_55),
.B1(n_56),
.B2(n_43),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g267 ( 
.A1(n_135),
.A2(n_151),
.B1(n_158),
.B2(n_172),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_65),
.B(n_55),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_150),
.B(n_156),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_104),
.A2(n_25),
.B1(n_41),
.B2(n_22),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_77),
.B(n_96),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_82),
.B(n_25),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_157),
.B(n_159),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_100),
.A2(n_22),
.B1(n_42),
.B2(n_33),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_163),
.B(n_183),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_92),
.B(n_24),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_164),
.B(n_171),
.Y(n_264)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_168),
.A2(n_186),
.B1(n_205),
.B2(n_66),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_58),
.B(n_47),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_114),
.A2(n_56),
.B1(n_58),
.B2(n_78),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_95),
.B(n_33),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_176),
.B(n_178),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_61),
.B(n_42),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_67),
.Y(n_181)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_123),
.B(n_38),
.C(n_34),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_99),
.A2(n_56),
.B1(n_47),
.B2(n_49),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_88),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_93),
.Y(n_189)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_105),
.B(n_49),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_191),
.B(n_0),
.Y(n_249)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_81),
.Y(n_192)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_73),
.Y(n_194)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_80),
.Y(n_198)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_78),
.A2(n_56),
.B1(n_48),
.B2(n_41),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_213),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_137),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_214),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_SL g312 ( 
.A(n_215),
.B(n_247),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_149),
.Y(n_216)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_216),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_217),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_154),
.A2(n_34),
.B1(n_75),
.B2(n_72),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_220),
.A2(n_224),
.B1(n_226),
.B2(n_231),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_L g223 ( 
.A1(n_135),
.A2(n_90),
.B1(n_70),
.B2(n_76),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_223),
.A2(n_233),
.B1(n_244),
.B2(n_132),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_156),
.A2(n_87),
.B1(n_121),
.B2(n_68),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_161),
.Y(n_225)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_225),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_180),
.A2(n_87),
.B1(n_121),
.B2(n_50),
.Y(n_226)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_139),
.Y(n_229)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_229),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_127),
.Y(n_230)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_230),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_129),
.A2(n_50),
.B1(n_45),
.B2(n_125),
.Y(n_231)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_126),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_232),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_186),
.A2(n_119),
.B1(n_106),
.B2(n_122),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_150),
.A2(n_13),
.B(n_18),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_234),
.B(n_249),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_129),
.Y(n_235)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_235),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_140),
.A2(n_50),
.B1(n_45),
.B2(n_60),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_237),
.A2(n_260),
.B(n_268),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_161),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_239),
.B(n_240),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_143),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_195),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_241),
.B(n_250),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_242),
.B(n_271),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_205),
.A2(n_50),
.B1(n_45),
.B2(n_54),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_195),
.Y(n_245)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_245),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_175),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_211),
.A2(n_50),
.B1(n_45),
.B2(n_54),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_248),
.A2(n_252),
.B1(n_258),
.B2(n_269),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_128),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_199),
.A2(n_50),
.B1(n_45),
.B2(n_2),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_146),
.Y(n_253)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_253),
.Y(n_325)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_130),
.Y(n_254)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_203),
.A2(n_6),
.B1(n_17),
.B2(n_2),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_255),
.A2(n_282),
.B1(n_283),
.B2(n_209),
.Y(n_294)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_148),
.Y(n_256)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_256),
.Y(n_306)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_257),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_134),
.A2(n_5),
.B1(n_14),
.B2(n_3),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_259),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_134),
.A2(n_183),
.B(n_193),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_204),
.Y(n_261)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_261),
.Y(n_328)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_160),
.Y(n_262)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_262),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_127),
.Y(n_263)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_141),
.Y(n_265)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_265),
.Y(n_338)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_190),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_270),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_140),
.A2(n_0),
.B(n_1),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_211),
.A2(n_12),
.B1(n_3),
.B2(n_4),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_145),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_152),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_272),
.B(n_274),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_147),
.A2(n_5),
.B1(n_12),
.B2(n_13),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_273),
.A2(n_212),
.B1(n_210),
.B2(n_184),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_200),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_200),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_277),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_149),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_276),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_143),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_162),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_278),
.B(n_279),
.Y(n_332)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_133),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_209),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_280),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_196),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_281),
.Y(n_331)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_197),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_196),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_193),
.A2(n_5),
.B1(n_13),
.B2(n_14),
.Y(n_284)
);

O2A1O1Ixp33_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_144),
.B(n_155),
.C(n_169),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_236),
.A2(n_136),
.B(n_131),
.C(n_138),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_289),
.A2(n_242),
.B(n_274),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_173),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_291),
.B(n_297),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_292),
.A2(n_315),
.B1(n_213),
.B2(n_214),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_222),
.A2(n_170),
.B1(n_206),
.B2(n_187),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_293),
.A2(n_319),
.B1(n_333),
.B2(n_235),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_249),
.B(n_285),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_182),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_300),
.B(n_303),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_190),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_177),
.C(n_165),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_304),
.B(n_314),
.C(n_326),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_305),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_308),
.B(n_283),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_238),
.B(n_243),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_339),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_268),
.B(n_174),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_313),
.B(n_337),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_237),
.B(n_172),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_243),
.A2(n_212),
.B1(n_210),
.B2(n_174),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_234),
.A2(n_206),
.B1(n_187),
.B2(n_184),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_243),
.B(n_142),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_233),
.A2(n_185),
.B1(n_153),
.B2(n_142),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_258),
.B(n_1),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_269),
.B(n_1),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_338),
.Y(n_340)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_340),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_308),
.A2(n_267),
.B1(n_223),
.B2(n_284),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_341),
.A2(n_355),
.B1(n_364),
.B2(n_367),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_295),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_342),
.B(n_380),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_314),
.A2(n_244),
.B(n_267),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_343),
.A2(n_346),
.B(n_353),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_267),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_344),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_313),
.A2(n_312),
.B1(n_287),
.B2(n_307),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_345),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_307),
.A2(n_267),
.B(n_277),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_338),
.Y(n_348)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_348),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_304),
.B(n_275),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_350),
.A2(n_351),
.B1(n_375),
.B2(n_376),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_296),
.A2(n_245),
.B1(n_225),
.B2(n_261),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_SL g353 ( 
.A(n_323),
.B(n_247),
.Y(n_353)
);

NAND2xp33_ASAP7_75t_R g394 ( 
.A(n_354),
.B(n_371),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_246),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_374),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_305),
.A2(n_282),
.B(n_270),
.Y(n_358)
);

BUFx5_ASAP7_75t_L g385 ( 
.A(n_358),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_323),
.Y(n_359)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_359),
.Y(n_413)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_298),
.Y(n_360)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_360),
.Y(n_381)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_329),
.Y(n_363)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_363),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_303),
.A2(n_266),
.B1(n_253),
.B2(n_229),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_330),
.A2(n_218),
.B1(n_227),
.B2(n_221),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_365),
.A2(n_366),
.B1(n_379),
.B2(n_355),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_300),
.A2(n_262),
.B1(n_227),
.B2(n_221),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_297),
.A2(n_228),
.B1(n_276),
.B2(n_216),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_SL g368 ( 
.A(n_287),
.B(n_251),
.C(n_219),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_378),
.C(n_287),
.Y(n_386)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_298),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_369),
.B(n_373),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_R g371 ( 
.A(n_291),
.B(n_232),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_323),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_329),
.Y(n_374)
);

BUFx8_ASAP7_75t_L g376 ( 
.A(n_288),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_327),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_377),
.A2(n_334),
.B1(n_321),
.B2(n_327),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_289),
.B(n_228),
.C(n_281),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_292),
.A2(n_279),
.B1(n_263),
.B2(n_230),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_311),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_386),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_370),
.B(n_322),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_393),
.C(n_402),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_339),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_414),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_390),
.A2(n_395),
.B1(n_412),
.B2(n_403),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_343),
.A2(n_372),
.B1(n_356),
.B2(n_344),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_391),
.A2(n_399),
.B1(n_407),
.B2(n_358),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_317),
.C(n_306),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_342),
.B(n_317),
.Y(n_397)
);

NAND3xp33_ASAP7_75t_L g443 ( 
.A(n_397),
.B(n_376),
.C(n_332),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_352),
.B(n_347),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_353),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_372),
.A2(n_290),
.B1(n_337),
.B2(n_302),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_306),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_344),
.A2(n_302),
.B1(n_315),
.B2(n_334),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_403),
.A2(n_375),
.B1(n_367),
.B2(n_360),
.Y(n_415)
);

AOI32xp33_ASAP7_75t_L g404 ( 
.A1(n_346),
.A2(n_318),
.A3(n_331),
.B1(n_309),
.B2(n_336),
.Y(n_404)
);

NOR2x1_ASAP7_75t_SL g444 ( 
.A(n_404),
.B(n_332),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_357),
.B(n_324),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_406),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_362),
.A2(n_309),
.B1(n_336),
.B2(n_321),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_345),
.B(n_320),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_410),
.B(n_411),
.C(n_373),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_349),
.B(n_320),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_347),
.B(n_298),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_415),
.A2(n_422),
.B1(n_429),
.B2(n_445),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_399),
.A2(n_341),
.B1(n_375),
.B2(n_349),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_418),
.A2(n_425),
.B1(n_426),
.B2(n_427),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_401),
.A2(n_409),
.B1(n_361),
.B2(n_391),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_419),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_383),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_420),
.B(n_414),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_423),
.B(n_437),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_387),
.B(n_368),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_435),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_408),
.A2(n_375),
.B1(n_365),
.B2(n_354),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_408),
.A2(n_378),
.B1(n_364),
.B2(n_379),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_382),
.A2(n_369),
.B1(n_359),
.B2(n_340),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_389),
.Y(n_430)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_430),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_384),
.A2(n_359),
.B1(n_366),
.B2(n_371),
.Y(n_431)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_431),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_388),
.A2(n_348),
.B1(n_376),
.B2(n_377),
.Y(n_432)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_432),
.Y(n_470)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_389),
.Y(n_433)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_433),
.Y(n_455)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_405),
.Y(n_434)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_434),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_398),
.B(n_402),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_405),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_439),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_393),
.B(n_410),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_441),
.C(n_386),
.Y(n_448)
);

OA22x2_ASAP7_75t_L g439 ( 
.A1(n_409),
.A2(n_404),
.B1(n_401),
.B2(n_382),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_394),
.A2(n_376),
.B(n_374),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_442),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_332),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_381),
.B(n_383),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_443),
.B(n_444),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_412),
.A2(n_363),
.B1(n_328),
.B2(n_301),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_448),
.B(n_452),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_449),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_421),
.B(n_417),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_450),
.B(n_459),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_438),
.B(n_396),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_418),
.A2(n_390),
.B1(n_381),
.B2(n_413),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_453),
.A2(n_469),
.B1(n_427),
.B2(n_415),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_437),
.B(n_413),
.Y(n_456)
);

AO21x1_ASAP7_75t_L g485 ( 
.A1(n_456),
.A2(n_440),
.B(n_430),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_421),
.B(n_392),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_458),
.C(n_465),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_428),
.B(n_299),
.C(n_328),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_417),
.B(n_400),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_442),
.Y(n_460)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_423),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_464),
.B(n_445),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_424),
.B(n_324),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_428),
.B(n_286),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_473),
.C(n_436),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_425),
.A2(n_385),
.B1(n_400),
.B2(n_299),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_441),
.B(n_286),
.C(n_335),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_433),
.Y(n_474)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_474),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_454),
.A2(n_439),
.B(n_416),
.Y(n_475)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_475),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_472),
.A2(n_444),
.B1(n_439),
.B2(n_419),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_478),
.A2(n_484),
.B1(n_493),
.B2(n_495),
.Y(n_505)
);

FAx1_ASAP7_75t_SL g479 ( 
.A(n_456),
.B(n_439),
.CI(n_429),
.CON(n_479),
.SN(n_479)
);

A2O1A1Ixp33_ASAP7_75t_L g501 ( 
.A1(n_479),
.A2(n_468),
.B(n_467),
.C(n_458),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_480),
.A2(n_468),
.B1(n_497),
.B2(n_446),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_481),
.B(n_486),
.Y(n_506)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_455),
.Y(n_483)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_483),
.Y(n_510)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_447),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_485),
.B(n_469),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_385),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_487),
.B(n_463),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_461),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_489),
.B(n_494),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_472),
.A2(n_301),
.B(n_325),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_490),
.A2(n_492),
.B(n_473),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_325),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_461),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_471),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_462),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_497),
.Y(n_516)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_453),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_448),
.C(n_466),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_498),
.B(n_511),
.C(n_476),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_477),
.B(n_491),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_504),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_501),
.A2(n_508),
.B(n_485),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_502),
.A2(n_478),
.B1(n_480),
.B2(n_487),
.Y(n_519)
);

XNOR2x1_ASAP7_75t_L g529 ( 
.A(n_503),
.B(n_512),
.Y(n_529)
);

BUFx24_ASAP7_75t_SL g504 ( 
.A(n_491),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_496),
.A2(n_446),
.B1(n_457),
.B2(n_452),
.Y(n_509)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_509),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_488),
.B(n_464),
.C(n_451),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_476),
.B(n_451),
.Y(n_512)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_513),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_484),
.B(n_463),
.Y(n_515)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_515),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_518),
.B(n_524),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g534 ( 
.A1(n_519),
.A2(n_505),
.B1(n_500),
.B2(n_492),
.Y(n_534)
);

FAx1_ASAP7_75t_SL g522 ( 
.A(n_509),
.B(n_479),
.CI(n_501),
.CON(n_522),
.SN(n_522)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_522),
.B(n_528),
.Y(n_540)
);

A2O1A1Ixp33_ASAP7_75t_SL g523 ( 
.A1(n_516),
.A2(n_503),
.B(n_507),
.C(n_479),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_523),
.A2(n_482),
.B1(n_502),
.B2(n_495),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_506),
.B(n_481),
.C(n_486),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_474),
.Y(n_525)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_525),
.Y(n_535)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_510),
.Y(n_527)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_527),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_513),
.B(n_465),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_530),
.B(n_511),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_506),
.B(n_492),
.C(n_483),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_531),
.B(n_508),
.C(n_490),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_498),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_533),
.B(n_537),
.Y(n_545)
);

OAI21xp33_ASAP7_75t_L g549 ( 
.A1(n_534),
.A2(n_526),
.B(n_523),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_542),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_530),
.B(n_512),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_539),
.B(n_518),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_541),
.B(n_520),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_524),
.B(n_482),
.C(n_493),
.Y(n_542)
);

MAJx2_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_335),
.C(n_230),
.Y(n_543)
);

NOR2x1_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_528),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_544),
.B(n_552),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_540),
.A2(n_526),
.B1(n_519),
.B2(n_522),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_547),
.B(n_549),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_548),
.B(n_539),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_550),
.B(n_535),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_542),
.B(n_521),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_551),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_517),
.C(n_529),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_525),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_553),
.B(n_523),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_557),
.B(n_558),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_546),
.B(n_538),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_545),
.B(n_537),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_559),
.A2(n_560),
.B(n_549),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_561),
.Y(n_566)
);

NOR3x1_ASAP7_75t_SL g562 ( 
.A(n_554),
.B(n_540),
.C(n_523),
.Y(n_562)
);

OAI21xp33_ASAP7_75t_SL g567 ( 
.A1(n_562),
.A2(n_564),
.B(n_565),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_556),
.A2(n_555),
.B(n_561),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_563),
.B(n_547),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_568),
.B(n_569),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_566),
.B(n_552),
.Y(n_569)
);

O2A1O1Ixp33_ASAP7_75t_SL g571 ( 
.A1(n_567),
.A2(n_522),
.B(n_544),
.C(n_536),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_571),
.A2(n_543),
.B(n_207),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_572),
.B(n_207),
.Y(n_573)
);

AO21x1_ASAP7_75t_L g574 ( 
.A1(n_573),
.A2(n_570),
.B(n_14),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_574),
.A2(n_14),
.B(n_18),
.Y(n_575)
);


endmodule