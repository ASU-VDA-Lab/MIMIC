module fake_netlist_5_712_n_1769 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1769);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1769;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1587;
wire n_1473;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_77),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_87),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_98),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_21),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_46),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_32),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_23),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_130),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_45),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_9),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_1),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_76),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_24),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_44),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_47),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_59),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_64),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_20),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_25),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_14),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_75),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_124),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_90),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_62),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_22),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_55),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_10),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_131),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_13),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_32),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_95),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_107),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_71),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_112),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_109),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_33),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_8),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_24),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_86),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_34),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_47),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_137),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_23),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_101),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_113),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_92),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_38),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_158),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_38),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_74),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_133),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_94),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_28),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_96),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_16),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_39),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_0),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_43),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_41),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_121),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_100),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_52),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_27),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_97),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_111),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_34),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_154),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_27),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_48),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_57),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_160),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_37),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_149),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_28),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_65),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_114),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_29),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_35),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_16),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_20),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_128),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_69),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_70),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_63),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_30),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_119),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_83),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_12),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_7),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_143),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_3),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_46),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_54),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_142),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_25),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_39),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_33),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_12),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_105),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_88),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_4),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_115),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_15),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_118),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_99),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_84),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_68),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_56),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_135),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_134),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_35),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_79),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_72),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_122),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_48),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_141),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_18),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_125),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_80),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_78),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_31),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_37),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_139),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_41),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_9),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_153),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_161),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_147),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_44),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_10),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_7),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_123),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_73),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_104),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_5),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_42),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_53),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_4),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_81),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_67),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_146),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_108),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_120),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_132),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_51),
.Y(n_318)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_145),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_45),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_18),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_3),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_36),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_182),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_250),
.Y(n_325)
);

INVxp33_ASAP7_75t_SL g326 ( 
.A(n_274),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_163),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_166),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_182),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_165),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_182),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_172),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_182),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_188),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_304),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_314),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_250),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_250),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_179),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_314),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_165),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_168),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_190),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_204),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_204),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_206),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_232),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_238),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_238),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_192),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_245),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_245),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_314),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_296),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_322),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_232),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_195),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_322),
.Y(n_361)
);

INVxp33_ASAP7_75t_SL g362 ( 
.A(n_179),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_202),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_218),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_233),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_218),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_323),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_175),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_184),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_191),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_194),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_196),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_209),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_211),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_167),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_225),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_231),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_212),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_214),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_206),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_215),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_233),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_219),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_176),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_247),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_314),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_251),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_223),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_224),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_236),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_261),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_314),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_254),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_320),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_239),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_288),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_319),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_254),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_264),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_270),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_301),
.Y(n_401)
);

OAI21x1_ASAP7_75t_L g402 ( 
.A1(n_337),
.A2(n_280),
.B(n_237),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_325),
.B(n_277),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_324),
.Y(n_404)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_337),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_325),
.B(n_280),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_337),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_324),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_331),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_329),
.B(n_277),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_348),
.B(n_280),
.Y(n_411)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_329),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_348),
.B(n_256),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_336),
.Y(n_415)
);

NAND2xp33_ASAP7_75t_L g416 ( 
.A(n_375),
.B(n_288),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_396),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_396),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_348),
.B(n_256),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_332),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_208),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_338),
.B(n_305),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_341),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_341),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_334),
.B(n_305),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_338),
.B(n_171),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_334),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_342),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_380),
.B(n_171),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_339),
.B(n_237),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_342),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_339),
.B(n_180),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_367),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_355),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_327),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_L g440 ( 
.A(n_375),
.B(n_308),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_330),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_384),
.B(n_176),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_326),
.B(n_210),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_343),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_355),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_367),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_355),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_356),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_328),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_356),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_369),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_356),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_380),
.B(n_180),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_386),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_364),
.B(n_266),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_375),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_362),
.B(n_333),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_349),
.A2(n_252),
.B1(n_170),
.B2(n_295),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_386),
.B(n_266),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_394),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_392),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_364),
.B(n_267),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_359),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_392),
.B(n_267),
.Y(n_465)
);

NAND2xp33_ASAP7_75t_R g466 ( 
.A(n_335),
.B(n_308),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_345),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_369),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_R g469 ( 
.A(n_352),
.B(n_321),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_366),
.B(n_282),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_370),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_371),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_366),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_405),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_405),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_414),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_414),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_466),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_404),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_456),
.B(n_357),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_405),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_407),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_406),
.B(n_360),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_405),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_409),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_414),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_407),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_404),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_405),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_460),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_406),
.B(n_363),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_406),
.B(n_378),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_411),
.B(n_433),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_408),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_456),
.B(n_357),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_408),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_460),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_408),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_403),
.A2(n_387),
.B1(n_368),
.B2(n_284),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_443),
.B(n_384),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_443),
.B(n_379),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_411),
.B(n_381),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_428),
.B(n_383),
.Y(n_506)
);

OR2x6_ASAP7_75t_L g507 ( 
.A(n_403),
.B(n_282),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_420),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_420),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_461),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_460),
.Y(n_511)
);

CKINVDCx11_ASAP7_75t_R g512 ( 
.A(n_444),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_432),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_465),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_465),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_465),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_432),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_428),
.B(n_388),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_465),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_432),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_438),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_438),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_465),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_461),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_420),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_425),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_425),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_425),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_441),
.A2(n_395),
.B1(n_389),
.B2(n_390),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_411),
.B(n_201),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_441),
.B(n_301),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_425),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_407),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_438),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_448),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_407),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_466),
.A2(n_306),
.B1(n_290),
.B2(n_295),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_472),
.B(n_306),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_448),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_448),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_472),
.B(n_176),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_426),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_454),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_412),
.Y(n_544)
);

AO22x2_ASAP7_75t_L g545 ( 
.A1(n_442),
.A2(n_294),
.B1(n_276),
.B2(n_309),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_453),
.B(n_234),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_426),
.Y(n_547)
);

BUFx6f_ASAP7_75t_SL g548 ( 
.A(n_424),
.Y(n_548)
);

BUFx4f_ASAP7_75t_L g549 ( 
.A(n_430),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_469),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_457),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_422),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_453),
.B(n_242),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_433),
.B(n_246),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_454),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_433),
.B(n_257),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_407),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_457),
.B(n_439),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_454),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_469),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_422),
.B(n_259),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_426),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_426),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_422),
.B(n_263),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_424),
.B(n_272),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_452),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_452),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_407),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_452),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_449),
.B(n_189),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_452),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_467),
.B(n_189),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_407),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_436),
.B(n_387),
.C(n_368),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_423),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_467),
.B(n_189),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_435),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_435),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_412),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_424),
.A2(n_297),
.B1(n_347),
.B2(n_207),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_416),
.B(n_344),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_423),
.B(n_193),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_435),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_427),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_435),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_427),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_415),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_458),
.A2(n_290),
.B1(n_170),
.B2(n_213),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_435),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_413),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_455),
.B(n_347),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_440),
.B(n_365),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_427),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_415),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_436),
.B(n_193),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_424),
.B(n_273),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_475),
.B(n_382),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_417),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_459),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_424),
.B(n_275),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_475),
.B(n_393),
.Y(n_601)
);

INVxp33_ASAP7_75t_L g602 ( 
.A(n_417),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_459),
.Y(n_603)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_427),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_418),
.B(n_398),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_427),
.B(n_278),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_459),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_418),
.B(n_401),
.Y(n_608)
);

AO22x2_ASAP7_75t_L g609 ( 
.A1(n_430),
.A2(n_302),
.B1(n_300),
.B2(n_293),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_464),
.Y(n_610)
);

OAI21xp33_ASAP7_75t_SL g611 ( 
.A1(n_402),
.A2(n_372),
.B(n_371),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_458),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_427),
.B(n_281),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_459),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_413),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_427),
.B(n_283),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_455),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_419),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_445),
.B(n_447),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_459),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_430),
.A2(n_207),
.B1(n_310),
.B2(n_391),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_462),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_419),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_462),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_493),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_496),
.B(n_445),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_563),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_486),
.A2(n_199),
.B1(n_164),
.B2(n_292),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_524),
.B(n_455),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_494),
.B(n_207),
.Y(n_630)
);

NOR2x1p5_ASAP7_75t_L g631 ( 
.A(n_550),
.B(n_311),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_563),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_495),
.B(n_207),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_594),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_504),
.B(n_181),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_489),
.B(n_437),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_493),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_476),
.B(n_310),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_566),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_566),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_496),
.B(n_445),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_507),
.A2(n_434),
.B1(n_430),
.B2(n_471),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_489),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_476),
.B(n_477),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_591),
.B(n_463),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_480),
.B(n_546),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_617),
.B(n_445),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_617),
.B(n_445),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_594),
.Y(n_649)
);

AO22x2_ASAP7_75t_L g650 ( 
.A1(n_531),
.A2(n_186),
.B1(n_185),
.B2(n_287),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_478),
.A2(n_463),
.B1(n_471),
.B2(n_317),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_500),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_581),
.B(n_181),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_478),
.B(n_479),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_511),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_477),
.B(n_484),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_575),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_SL g658 ( 
.A(n_550),
.B(n_213),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_484),
.B(n_310),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_505),
.B(n_187),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_487),
.B(n_310),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_591),
.B(n_463),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_479),
.B(n_445),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_509),
.B(n_445),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_509),
.B(n_447),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_508),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_525),
.B(n_447),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_577),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_508),
.B(n_437),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_525),
.B(n_447),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_487),
.B(n_447),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_575),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_492),
.B(n_447),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_492),
.B(n_447),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_503),
.B(n_187),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_552),
.A2(n_198),
.B1(n_200),
.B2(n_216),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_560),
.B(n_319),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_514),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_514),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_515),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_552),
.B(n_450),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_515),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_577),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_548),
.A2(n_471),
.B1(n_289),
.B2(n_286),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_553),
.B(n_450),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_SL g686 ( 
.A(n_560),
.B(n_252),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_510),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_548),
.A2(n_307),
.B1(n_299),
.B2(n_291),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_516),
.B(n_450),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_524),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_516),
.B(n_450),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_519),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_574),
.B(n_313),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_519),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_523),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_523),
.B(n_450),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_549),
.B(n_450),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_578),
.Y(n_698)
);

O2A1O1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_611),
.A2(n_410),
.B(n_429),
.C(n_474),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_530),
.B(n_450),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_578),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_554),
.B(n_430),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_506),
.B(n_313),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_587),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_556),
.B(n_434),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_590),
.B(n_434),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_513),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_590),
.B(n_434),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_615),
.B(n_434),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_549),
.B(n_319),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_605),
.B(n_205),
.C(n_473),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_513),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_615),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_618),
.Y(n_714)
);

A2O1A1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_611),
.A2(n_402),
.B(n_473),
.C(n_470),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_618),
.B(n_462),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_518),
.B(n_169),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_608),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_517),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_623),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_623),
.B(n_462),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_587),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_598),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_561),
.B(n_462),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_526),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_565),
.B(n_319),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_SL g727 ( 
.A1(n_588),
.A2(n_253),
.B1(n_262),
.B2(n_311),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_564),
.B(n_421),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_507),
.A2(n_596),
.B1(n_600),
.B2(n_548),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_619),
.B(n_319),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_529),
.B(n_319),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_583),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_597),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_481),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_601),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_526),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_507),
.A2(n_402),
.B1(n_262),
.B2(n_253),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_541),
.B(n_173),
.Y(n_738)
);

BUFx8_ASAP7_75t_L g739 ( 
.A(n_512),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_545),
.Y(n_740)
);

BUFx5_ASAP7_75t_L g741 ( 
.A(n_527),
.Y(n_741)
);

AND2x6_ASAP7_75t_L g742 ( 
.A(n_536),
.B(n_217),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_527),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_507),
.B(n_421),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_507),
.B(n_431),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_528),
.B(n_319),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_609),
.A2(n_222),
.B1(n_315),
.B2(n_279),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_533),
.B(n_431),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_L g749 ( 
.A(n_621),
.B(n_221),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_517),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_573),
.B(n_604),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_610),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_528),
.B(n_226),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_583),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_609),
.A2(n_243),
.B1(n_260),
.B2(n_255),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_585),
.Y(n_756)
);

INVx8_ASAP7_75t_L g757 ( 
.A(n_488),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_532),
.B(n_410),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_532),
.B(n_248),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_542),
.B(n_429),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_542),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_547),
.B(n_562),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_547),
.B(n_249),
.Y(n_763)
);

NAND3x1_ASAP7_75t_L g764 ( 
.A(n_537),
.B(n_376),
.C(n_372),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_481),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_520),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_562),
.B(n_412),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_567),
.B(n_412),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_585),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_606),
.B(n_174),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_567),
.B(n_446),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_569),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_483),
.B(n_177),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_595),
.B(n_446),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_610),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_569),
.B(n_412),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_609),
.A2(n_502),
.B1(n_580),
.B2(n_545),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_571),
.B(n_451),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_545),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_602),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_571),
.B(n_451),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_536),
.B(n_468),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_545),
.A2(n_474),
.B1(n_470),
.B2(n_468),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_520),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_584),
.B(n_412),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_482),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_558),
.B(n_167),
.Y(n_787)
);

BUFx12f_ASAP7_75t_L g788 ( 
.A(n_612),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_L g789 ( 
.A(n_592),
.B(n_498),
.C(n_538),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_609),
.A2(n_321),
.B1(n_167),
.B2(n_183),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_643),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_646),
.A2(n_576),
.B1(n_572),
.B2(n_551),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_657),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_757),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_672),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_646),
.B(n_521),
.Y(n_796)
);

NOR2x1p5_ASAP7_75t_L g797 ( 
.A(n_789),
.B(n_612),
.Y(n_797)
);

AO22x1_ASAP7_75t_L g798 ( 
.A1(n_635),
.A2(n_271),
.B1(n_228),
.B2(n_227),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_643),
.Y(n_799)
);

OAI22x1_ASAP7_75t_SL g800 ( 
.A1(n_775),
.A2(n_318),
.B1(n_197),
.B2(n_203),
.Y(n_800)
);

AND2x6_ASAP7_75t_SL g801 ( 
.A(n_717),
.B(n_373),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_739),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_715),
.A2(n_613),
.B(n_616),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_625),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_682),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_645),
.B(n_521),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_662),
.B(n_551),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_625),
.Y(n_808)
);

INVxp33_ASAP7_75t_L g809 ( 
.A(n_686),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_693),
.A2(n_537),
.B1(n_582),
.B2(n_620),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_626),
.B(n_522),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_652),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_641),
.B(n_522),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_652),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_757),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_636),
.B(n_570),
.Y(n_816)
);

AOI211xp5_ASAP7_75t_L g817 ( 
.A1(n_727),
.A2(n_265),
.B(n_220),
.C(n_229),
.Y(n_817)
);

CKINVDCx8_ASAP7_75t_R g818 ( 
.A(n_757),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_666),
.Y(n_819)
);

AND2x6_ASAP7_75t_SL g820 ( 
.A(n_717),
.B(n_373),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_695),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_704),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_695),
.B(n_534),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_713),
.B(n_534),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_682),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_707),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_636),
.B(n_374),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_637),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_690),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_722),
.Y(n_830)
);

BUFx8_ASAP7_75t_L g831 ( 
.A(n_788),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_733),
.B(n_551),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_780),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_635),
.B(n_551),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_707),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_653),
.A2(n_536),
.B(n_568),
.C(n_593),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_712),
.Y(n_837)
);

INVxp67_ASAP7_75t_SL g838 ( 
.A(n_644),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_655),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_714),
.B(n_535),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_629),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_669),
.B(n_374),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_687),
.B(n_376),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_723),
.B(n_377),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_658),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_634),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_740),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_649),
.B(n_584),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_678),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_735),
.B(n_718),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_739),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_666),
.Y(n_852)
);

BUFx12f_ASAP7_75t_SL g853 ( 
.A(n_787),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_679),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_680),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_669),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_752),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_720),
.B(n_535),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_774),
.B(n_377),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_654),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_719),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_653),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_779),
.A2(n_622),
.B1(n_614),
.B2(n_607),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_631),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_750),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_774),
.B(n_385),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_692),
.B(n_539),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_702),
.A2(n_485),
.B(n_490),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_734),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_766),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_694),
.B(n_539),
.Y(n_871)
);

INVx5_ASAP7_75t_L g872 ( 
.A(n_742),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_703),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_SL g874 ( 
.A(n_675),
.B(n_178),
.C(n_230),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_725),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_675),
.B(n_385),
.Y(n_876)
);

AO21x2_ASAP7_75t_L g877 ( 
.A1(n_710),
.A2(n_491),
.B(n_482),
.Y(n_877)
);

OAI22xp33_ASAP7_75t_L g878 ( 
.A1(n_783),
.A2(n_235),
.B1(n_240),
.B2(n_241),
.Y(n_878)
);

NAND2x1p5_ASAP7_75t_L g879 ( 
.A(n_644),
.B(n_485),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_766),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_736),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_703),
.B(n_183),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_656),
.B(n_540),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_734),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_681),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_656),
.B(n_540),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_743),
.Y(n_887)
);

AND2x6_ASAP7_75t_SL g888 ( 
.A(n_773),
.B(n_738),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_761),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_772),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_660),
.B(n_584),
.Y(n_891)
);

NOR2xp67_ASAP7_75t_L g892 ( 
.A(n_660),
.B(n_391),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_677),
.A2(n_557),
.B1(n_485),
.B2(n_603),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_777),
.B(n_584),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_782),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_742),
.Y(n_896)
);

BUFx5_ASAP7_75t_L g897 ( 
.A(n_742),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_773),
.B(n_557),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_628),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_771),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_738),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_777),
.B(n_584),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_778),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_731),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_728),
.B(n_543),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_784),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_705),
.B(n_758),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_737),
.B(n_193),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_729),
.A2(n_557),
.B1(n_614),
.B2(n_603),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_781),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_715),
.A2(n_499),
.B(n_491),
.C(n_497),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_737),
.B(n_285),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_765),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_711),
.B(n_399),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_684),
.B(n_399),
.Y(n_915)
);

NAND2xp33_ASAP7_75t_L g916 ( 
.A(n_742),
.B(n_741),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_742),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_760),
.B(n_543),
.Y(n_918)
);

INVxp67_ASAP7_75t_SL g919 ( 
.A(n_647),
.Y(n_919)
);

AND2x4_ASAP7_75t_SL g920 ( 
.A(n_651),
.B(n_285),
.Y(n_920)
);

INVx3_ASAP7_75t_SL g921 ( 
.A(n_650),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_762),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_744),
.B(n_400),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_762),
.Y(n_924)
);

INVx5_ASAP7_75t_L g925 ( 
.A(n_765),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_745),
.B(n_400),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_731),
.B(n_244),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_784),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_688),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_642),
.B(n_285),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_699),
.A2(n_624),
.B(n_599),
.C(n_589),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_700),
.B(n_555),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_724),
.B(n_555),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_650),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_747),
.A2(n_497),
.B1(n_499),
.B2(n_501),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_648),
.B(n_559),
.Y(n_936)
);

BUFx4f_ASAP7_75t_L g937 ( 
.A(n_786),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_697),
.B(n_767),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_706),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_770),
.A2(n_624),
.B1(n_599),
.B2(n_589),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_790),
.B(n_183),
.Y(n_941)
);

INVxp67_ASAP7_75t_SL g942 ( 
.A(n_751),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_708),
.B(n_709),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_650),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_764),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_663),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_786),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_642),
.B(n_312),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_741),
.B(n_559),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_627),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_632),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_747),
.B(n_312),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_639),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_755),
.A2(n_258),
.B1(n_268),
.B2(n_269),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_755),
.B(n_312),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_630),
.B(n_298),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_790),
.A2(n_303),
.B1(n_354),
.B2(n_353),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_630),
.B(n_316),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_633),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_640),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_633),
.A2(n_501),
.B1(n_316),
.B2(n_397),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_741),
.B(n_316),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_668),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_664),
.B(n_0),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_683),
.Y(n_965)
);

NOR2x1p5_ASAP7_75t_L g966 ( 
.A(n_665),
.B(n_346),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_698),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_741),
.B(n_586),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_667),
.B(n_346),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_701),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_907),
.B(n_900),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_812),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_804),
.Y(n_973)
);

OR2x6_ASAP7_75t_L g974 ( 
.A(n_833),
.B(n_746),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_907),
.B(n_670),
.Y(n_975)
);

NAND3xp33_ASAP7_75t_SL g976 ( 
.A(n_873),
.B(n_676),
.C(n_726),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_943),
.A2(n_942),
.B(n_916),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_850),
.B(n_767),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_808),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_901),
.B(n_741),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_821),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_862),
.A2(n_921),
.B1(n_792),
.B2(n_902),
.Y(n_982)
);

AND3x2_ASAP7_75t_L g983 ( 
.A(n_941),
.B(n_350),
.C(n_351),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_814),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_847),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_826),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_927),
.A2(n_726),
.B(n_696),
.C(n_691),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_793),
.B(n_746),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_943),
.A2(n_697),
.B(n_685),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_874),
.A2(n_753),
.B(n_759),
.C(n_763),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_860),
.B(n_741),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_874),
.A2(n_753),
.B(n_759),
.C(n_763),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_847),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_835),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_942),
.A2(n_671),
.B(n_673),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_908),
.A2(n_638),
.B(n_661),
.C(n_659),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_860),
.B(n_716),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_832),
.B(n_768),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_919),
.A2(n_868),
.B(n_813),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_903),
.B(n_748),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_841),
.B(n_768),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_841),
.B(n_809),
.Y(n_1002)
);

BUFx4f_ASAP7_75t_SL g1003 ( 
.A(n_851),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_912),
.A2(n_661),
.B(n_638),
.C(n_659),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_818),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_856),
.B(n_721),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_882),
.A2(n_689),
.B(n_754),
.C(n_769),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_828),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_919),
.A2(n_674),
.B(n_785),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_R g1010 ( 
.A(n_857),
.B(n_749),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_852),
.B(n_756),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_852),
.B(n_732),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_910),
.B(n_674),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_921),
.A2(n_776),
.B1(n_785),
.B2(n_730),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_837),
.Y(n_1015)
);

INVx1_ASAP7_75t_SL g1016 ( 
.A(n_829),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_868),
.A2(n_730),
.B(n_776),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_892),
.B(n_586),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_853),
.B(n_1),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_944),
.A2(n_397),
.B1(n_350),
.B2(n_358),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_811),
.A2(n_586),
.B(n_412),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_791),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_811),
.A2(n_586),
.B(n_412),
.Y(n_1023)
);

CKINVDCx8_ASAP7_75t_R g1024 ( 
.A(n_802),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_816),
.B(n_351),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_797),
.A2(n_361),
.B1(n_358),
.B2(n_354),
.Y(n_1026)
);

NOR2x1_ASAP7_75t_L g1027 ( 
.A(n_819),
.B(n_353),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_861),
.Y(n_1028)
);

NAND2x1p5_ASAP7_75t_L g1029 ( 
.A(n_852),
.B(n_819),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_956),
.A2(n_361),
.B(n_586),
.C(n_8),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_865),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_923),
.B(n_2),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_894),
.A2(n_2),
.B1(n_6),
.B2(n_11),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_923),
.B(n_6),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_816),
.B(n_795),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_876),
.B(n_11),
.Y(n_1036)
);

NOR2x1_ASAP7_75t_SL g1037 ( 
.A(n_872),
.B(n_579),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_904),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_878),
.A2(n_17),
.B(n_19),
.C(n_21),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_843),
.B(n_17),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_810),
.B(n_579),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_899),
.B(n_579),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_926),
.B(n_19),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_791),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_926),
.B(n_22),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_813),
.A2(n_579),
.B(n_544),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_791),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_834),
.B(n_544),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_839),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_L g1050 ( 
.A(n_798),
.B(n_544),
.C(n_29),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_799),
.B(n_544),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_878),
.A2(n_26),
.B(n_30),
.C(n_31),
.Y(n_1052)
);

INVx8_ASAP7_75t_L g1053 ( 
.A(n_799),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_831),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_870),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_888),
.B(n_36),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_939),
.B(n_40),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_799),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_880),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_906),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_952),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_838),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_859),
.B(n_49),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_929),
.A2(n_103),
.B1(n_58),
.B2(n_60),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_849),
.Y(n_1065)
);

BUFx8_ASAP7_75t_L g1066 ( 
.A(n_864),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_854),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_794),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_822),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_949),
.A2(n_110),
.B(n_61),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_859),
.B(n_116),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_866),
.B(n_50),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_955),
.A2(n_66),
.B(n_82),
.C(n_85),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_945),
.B(n_89),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_949),
.A2(n_91),
.B(n_93),
.Y(n_1075)
);

CKINVDCx14_ASAP7_75t_R g1076 ( 
.A(n_815),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_932),
.A2(n_102),
.B(n_126),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_959),
.A2(n_958),
.B1(n_807),
.B2(n_945),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_845),
.B(n_127),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_855),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_898),
.B(n_129),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_911),
.A2(n_136),
.B(n_138),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_830),
.B(n_144),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_838),
.A2(n_148),
.B1(n_150),
.B2(n_934),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_937),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_796),
.A2(n_817),
.B1(n_905),
.B2(n_805),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_896),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_895),
.B(n_796),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_930),
.A2(n_948),
.B(n_954),
.C(n_957),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_928),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_801),
.B(n_820),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_827),
.B(n_842),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_915),
.A2(n_866),
.B1(n_842),
.B2(n_827),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_846),
.B(n_915),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_905),
.B(n_875),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_932),
.A2(n_933),
.B(n_891),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_922),
.A2(n_924),
.B(n_964),
.C(n_920),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_967),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_881),
.B(n_887),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_967),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_805),
.A2(n_825),
.B1(n_918),
.B2(n_935),
.Y(n_1101)
);

AO32x2_ASAP7_75t_L g1102 ( 
.A1(n_957),
.A2(n_954),
.A3(n_913),
.B1(n_869),
.B2(n_803),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_937),
.Y(n_1103)
);

INVxp67_ASAP7_75t_SL g1104 ( 
.A(n_825),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_918),
.A2(n_935),
.B1(n_806),
.B2(n_890),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_896),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_889),
.Y(n_1107)
);

OAI21xp33_ASAP7_75t_L g1108 ( 
.A1(n_844),
.A2(n_914),
.B(n_806),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_SL g1109 ( 
.A(n_800),
.B(n_848),
.C(n_962),
.Y(n_1109)
);

AO21x1_ASAP7_75t_L g1110 ( 
.A1(n_938),
.A2(n_803),
.B(n_911),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_966),
.A2(n_836),
.B(n_965),
.C(n_960),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_933),
.A2(n_936),
.B(n_823),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_969),
.A2(n_885),
.B1(n_946),
.B2(n_950),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_885),
.B(n_946),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_885),
.B(n_969),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_863),
.A2(n_872),
.B1(n_938),
.B2(n_824),
.Y(n_1116)
);

AO21x2_ASAP7_75t_L g1117 ( 
.A1(n_999),
.A2(n_909),
.B(n_931),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_971),
.A2(n_872),
.B1(n_869),
.B2(n_913),
.Y(n_1118)
);

AOI21x1_ASAP7_75t_SL g1119 ( 
.A1(n_1081),
.A2(n_824),
.B(n_840),
.Y(n_1119)
);

O2A1O1Ixp5_ASAP7_75t_L g1120 ( 
.A1(n_1097),
.A2(n_968),
.B(n_936),
.C(n_871),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1092),
.B(n_1063),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_971),
.B(n_840),
.Y(n_1122)
);

AO31x2_ASAP7_75t_L g1123 ( 
.A1(n_1110),
.A2(n_871),
.A3(n_867),
.B(n_823),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_1085),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1017),
.A2(n_867),
.B(n_883),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1092),
.B(n_970),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1088),
.B(n_858),
.Y(n_1127)
);

NAND2x1_ASAP7_75t_L g1128 ( 
.A(n_1106),
.B(n_884),
.Y(n_1128)
);

CKINVDCx11_ASAP7_75t_R g1129 ( 
.A(n_1024),
.Y(n_1129)
);

BUFx10_ASAP7_75t_L g1130 ( 
.A(n_1002),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1095),
.A2(n_858),
.B1(n_884),
.B2(n_879),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_975),
.B(n_886),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1089),
.A2(n_951),
.B(n_953),
.C(n_940),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_995),
.A2(n_877),
.B(n_925),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1096),
.A2(n_877),
.B(n_925),
.Y(n_1135)
);

CKINVDCx12_ASAP7_75t_R g1136 ( 
.A(n_1040),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_987),
.A2(n_925),
.B(n_893),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1000),
.B(n_1105),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_990),
.A2(n_961),
.B(n_963),
.C(n_947),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1105),
.B(n_925),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1116),
.A2(n_917),
.B(n_897),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1108),
.A2(n_831),
.B1(n_917),
.B2(n_897),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1049),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_992),
.A2(n_897),
.B(n_917),
.C(n_978),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1013),
.B(n_897),
.Y(n_1145)
);

O2A1O1Ixp5_ASAP7_75t_L g1146 ( 
.A1(n_1086),
.A2(n_897),
.B(n_980),
.C(n_1057),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1086),
.B(n_897),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1041),
.A2(n_1009),
.B(n_1007),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1016),
.B(n_1078),
.Y(n_1149)
);

BUFx8_ASAP7_75t_L g1150 ( 
.A(n_1054),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1082),
.A2(n_1021),
.B(n_1023),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_996),
.A2(n_1004),
.B(n_1101),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1101),
.A2(n_1046),
.B(n_1042),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_997),
.A2(n_991),
.B(n_1006),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1014),
.A2(n_1048),
.B(n_1077),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1014),
.A2(n_1070),
.B(n_1075),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1072),
.B(n_1025),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1090),
.A2(n_1012),
.B(n_1011),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_998),
.B(n_1114),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1115),
.B(n_973),
.Y(n_1160)
);

INVx3_ASAP7_75t_SL g1161 ( 
.A(n_1005),
.Y(n_1161)
);

AO21x2_ASAP7_75t_L g1162 ( 
.A1(n_1111),
.A2(n_1030),
.B(n_976),
.Y(n_1162)
);

AOI21x1_ASAP7_75t_SL g1163 ( 
.A1(n_1032),
.A2(n_1045),
.B(n_1043),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1085),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_979),
.B(n_981),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_982),
.A2(n_1084),
.B(n_1034),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_1016),
.Y(n_1167)
);

AO21x1_ASAP7_75t_L g1168 ( 
.A1(n_1084),
.A2(n_1033),
.B(n_982),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1099),
.B(n_1065),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_SL g1170 ( 
.A1(n_1073),
.A2(n_1052),
.B(n_1039),
.Y(n_1170)
);

NOR4xp25_ASAP7_75t_L g1171 ( 
.A(n_1062),
.B(n_1061),
.C(n_1038),
.D(n_1056),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_1050),
.B(n_1091),
.C(n_1109),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1018),
.A2(n_1051),
.B(n_972),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1094),
.B(n_1085),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1069),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1058),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_984),
.A2(n_1031),
.B(n_1060),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1067),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1094),
.B(n_1103),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_986),
.A2(n_994),
.B(n_1059),
.Y(n_1180)
);

BUFx8_ASAP7_75t_L g1181 ( 
.A(n_1103),
.Y(n_1181)
);

NAND3x1_ASAP7_75t_L g1182 ( 
.A(n_1074),
.B(n_1019),
.C(n_1093),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1015),
.A2(n_1028),
.B(n_1055),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1080),
.B(n_1107),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1037),
.A2(n_1104),
.B(n_1113),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1058),
.Y(n_1186)
);

AO22x2_ASAP7_75t_L g1187 ( 
.A1(n_1062),
.A2(n_1036),
.B1(n_1102),
.B2(n_985),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1103),
.B(n_1010),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1027),
.A2(n_1029),
.B(n_1047),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_L g1190 ( 
.A(n_1026),
.B(n_1079),
.C(n_983),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1025),
.B(n_1001),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1020),
.A2(n_1071),
.B(n_1083),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1064),
.A2(n_1098),
.B(n_1100),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_1035),
.B(n_993),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_988),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_974),
.A2(n_988),
.B(n_1102),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1029),
.A2(n_1022),
.B(n_1047),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1022),
.A2(n_1102),
.B(n_1087),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_974),
.A2(n_988),
.A3(n_1087),
.B(n_1106),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_974),
.A2(n_1087),
.B(n_1076),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1044),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_1068),
.B(n_1053),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1053),
.A2(n_1106),
.B(n_1044),
.C(n_1066),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1053),
.A2(n_1044),
.B(n_1066),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1003),
.B(n_971),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1008),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_982),
.A2(n_635),
.B(n_718),
.C(n_733),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1092),
.B(n_841),
.Y(n_1208)
);

AOI21x1_ASAP7_75t_L g1209 ( 
.A1(n_977),
.A2(n_999),
.B(n_989),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1017),
.A2(n_911),
.B(n_999),
.Y(n_1210)
);

NOR2xp67_ASAP7_75t_L g1211 ( 
.A(n_1069),
.B(n_657),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1090),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1002),
.B(n_733),
.Y(n_1213)
);

NOR4xp25_ASAP7_75t_L g1214 ( 
.A(n_1039),
.B(n_1052),
.C(n_874),
.D(n_1089),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1002),
.B(n_733),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1089),
.A2(n_635),
.B(n_653),
.C(n_792),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1068),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1058),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1092),
.B(n_841),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1017),
.A2(n_911),
.B(n_999),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1008),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_989),
.A2(n_977),
.B(n_1112),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1089),
.A2(n_635),
.B(n_653),
.C(n_792),
.Y(n_1223)
);

NAND2xp33_ASAP7_75t_L g1224 ( 
.A(n_971),
.B(n_873),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_1005),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1090),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1002),
.B(n_733),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1017),
.A2(n_911),
.B(n_999),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_971),
.B(n_1088),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1008),
.Y(n_1230)
);

OA21x2_ASAP7_75t_L g1231 ( 
.A1(n_999),
.A2(n_1110),
.B(n_803),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1008),
.Y(n_1232)
);

CKINVDCx11_ASAP7_75t_R g1233 ( 
.A(n_1024),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1092),
.B(n_841),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1090),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1017),
.A2(n_911),
.B(n_999),
.Y(n_1236)
);

AOI221xp5_ASAP7_75t_SL g1237 ( 
.A1(n_1039),
.A2(n_878),
.B1(n_727),
.B2(n_1052),
.C(n_817),
.Y(n_1237)
);

BUFx8_ASAP7_75t_L g1238 ( 
.A(n_1054),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_989),
.A2(n_977),
.B(n_1112),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_L g1240 ( 
.A(n_1069),
.B(n_657),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_989),
.A2(n_977),
.B(n_1112),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1089),
.A2(n_635),
.B(n_653),
.C(n_792),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_971),
.A2(n_873),
.B1(n_901),
.B2(n_862),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1017),
.A2(n_911),
.B(n_999),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1094),
.B(n_1092),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_971),
.B(n_1088),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_971),
.B(n_1088),
.Y(n_1247)
);

INVxp67_ASAP7_75t_SL g1248 ( 
.A(n_971),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1017),
.A2(n_911),
.B(n_999),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1089),
.A2(n_635),
.B(n_653),
.C(n_792),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1068),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1092),
.B(n_841),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_971),
.B(n_1088),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1017),
.A2(n_911),
.B(n_999),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1017),
.A2(n_911),
.B(n_999),
.Y(n_1255)
);

NAND2x1p5_ASAP7_75t_L g1256 ( 
.A(n_1087),
.B(n_852),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1151),
.A2(n_1134),
.B(n_1135),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1216),
.A2(n_1242),
.B(n_1223),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1177),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1134),
.A2(n_1135),
.B(n_1209),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_1124),
.Y(n_1261)
);

BUFx2_ASAP7_75t_SL g1262 ( 
.A(n_1225),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1213),
.A2(n_1227),
.B1(n_1215),
.B2(n_1243),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1210),
.A2(n_1228),
.B(n_1220),
.Y(n_1264)
);

AO21x2_ASAP7_75t_L g1265 ( 
.A1(n_1222),
.A2(n_1241),
.B(n_1239),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_SL g1266 ( 
.A1(n_1168),
.A2(n_1166),
.B(n_1170),
.Y(n_1266)
);

INVx5_ASAP7_75t_L g1267 ( 
.A(n_1124),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1180),
.Y(n_1268)
);

NAND2x1p5_ASAP7_75t_L g1269 ( 
.A(n_1204),
.B(n_1176),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1236),
.A2(n_1249),
.B(n_1244),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1243),
.B(n_1207),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1254),
.A2(n_1255),
.B(n_1125),
.Y(n_1272)
);

INVxp33_ASAP7_75t_L g1273 ( 
.A(n_1191),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1208),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1250),
.A2(n_1214),
.B(n_1166),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1224),
.A2(n_1149),
.B(n_1171),
.C(n_1192),
.Y(n_1276)
);

OAI221xp5_ASAP7_75t_L g1277 ( 
.A1(n_1237),
.A2(n_1172),
.B1(n_1190),
.B2(n_1205),
.C(n_1142),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1248),
.A2(n_1247),
.B1(n_1253),
.B2(n_1246),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1195),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1222),
.A2(n_1239),
.B(n_1241),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1183),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1181),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1159),
.B(n_1138),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1144),
.A2(n_1148),
.B(n_1137),
.Y(n_1284)
);

AO32x2_ASAP7_75t_L g1285 ( 
.A1(n_1131),
.A2(n_1118),
.A3(n_1187),
.B1(n_1196),
.B2(n_1123),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1157),
.B(n_1121),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1137),
.A2(n_1141),
.B(n_1147),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1219),
.B(n_1234),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1152),
.A2(n_1153),
.A3(n_1147),
.B(n_1140),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1217),
.Y(n_1290)
);

AO31x2_ASAP7_75t_L g1291 ( 
.A1(n_1152),
.A2(n_1140),
.A3(n_1131),
.B(n_1133),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1252),
.Y(n_1292)
);

INVx6_ASAP7_75t_L g1293 ( 
.A(n_1181),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1229),
.A2(n_1246),
.B(n_1247),
.C(n_1253),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1141),
.A2(n_1173),
.B(n_1119),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1124),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1229),
.B(n_1159),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1156),
.A2(n_1155),
.B(n_1154),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1200),
.B(n_1185),
.Y(n_1299)
);

OAI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1169),
.A2(n_1122),
.B1(n_1127),
.B2(n_1138),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1143),
.Y(n_1301)
);

AOI22x1_ASAP7_75t_L g1302 ( 
.A1(n_1187),
.A2(n_1200),
.B1(n_1193),
.B2(n_1178),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1251),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1146),
.A2(n_1120),
.B(n_1139),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1199),
.B(n_1174),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1199),
.B(n_1174),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1206),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1221),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1196),
.A2(n_1117),
.B(n_1118),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1199),
.B(n_1179),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1158),
.A2(n_1163),
.B(n_1145),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1202),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1230),
.Y(n_1313)
);

AND2x2_ASAP7_75t_SL g1314 ( 
.A(n_1231),
.B(n_1122),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1232),
.Y(n_1315)
);

CKINVDCx6p67_ASAP7_75t_R g1316 ( 
.A(n_1129),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1127),
.A2(n_1169),
.B(n_1132),
.C(n_1160),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1205),
.A2(n_1167),
.B1(n_1194),
.B2(n_1160),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1126),
.B(n_1245),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1165),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1165),
.Y(n_1321)
);

BUFx2_ASAP7_75t_R g1322 ( 
.A(n_1161),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1193),
.A2(n_1189),
.B(n_1235),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1212),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1188),
.B(n_1175),
.Y(n_1325)
);

NAND3xp33_ASAP7_75t_SL g1326 ( 
.A(n_1203),
.B(n_1226),
.C(n_1256),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1197),
.A2(n_1128),
.B(n_1256),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1211),
.A2(n_1240),
.B(n_1201),
.Y(n_1328)
);

BUFx12f_ASAP7_75t_L g1329 ( 
.A(n_1233),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1176),
.A2(n_1218),
.B(n_1186),
.Y(n_1330)
);

INVx4_ASAP7_75t_L g1331 ( 
.A(n_1164),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1186),
.A2(n_1117),
.B(n_1123),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1136),
.B(n_1130),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1162),
.A2(n_873),
.B1(n_862),
.B2(n_901),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1150),
.A2(n_1238),
.B(n_1151),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1150),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_SL g1337 ( 
.A(n_1238),
.B(n_775),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1243),
.B(n_873),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1184),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1168),
.A2(n_1166),
.B1(n_941),
.B2(n_873),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1216),
.A2(n_1242),
.B(n_1223),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1184),
.Y(n_1342)
);

AOI221xp5_ASAP7_75t_L g1343 ( 
.A1(n_1214),
.A2(n_727),
.B1(n_443),
.B2(n_873),
.C(n_901),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1177),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1129),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1182),
.A2(n_862),
.B1(n_901),
.B2(n_873),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1248),
.A2(n_873),
.B1(n_901),
.B2(n_537),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1191),
.B(n_1159),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1216),
.A2(n_1242),
.B(n_1223),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1151),
.A2(n_1134),
.B(n_1135),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1198),
.Y(n_1351)
);

OA21x2_ASAP7_75t_L g1352 ( 
.A1(n_1222),
.A2(n_1241),
.B(n_1239),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1168),
.A2(n_1166),
.B1(n_941),
.B2(n_873),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1216),
.A2(n_1242),
.B(n_1223),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1129),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1248),
.B(n_1229),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1151),
.A2(n_1134),
.B(n_1135),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1191),
.B(n_1157),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_SL g1359 ( 
.A1(n_1216),
.A2(n_1242),
.B(n_1250),
.C(n_1223),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1177),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1195),
.B(n_1199),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1184),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1184),
.Y(n_1363)
);

BUFx2_ASAP7_75t_R g1364 ( 
.A(n_1161),
.Y(n_1364)
);

OAI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1248),
.A2(n_873),
.B1(n_901),
.B2(n_537),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1184),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1184),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1177),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1213),
.A2(n_873),
.B1(n_862),
.B2(n_901),
.Y(n_1369)
);

INVx4_ASAP7_75t_L g1370 ( 
.A(n_1124),
.Y(n_1370)
);

AOI21xp33_ASAP7_75t_L g1371 ( 
.A1(n_1207),
.A2(n_635),
.B(n_873),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1151),
.A2(n_1134),
.B(n_1135),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1124),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1151),
.A2(n_1134),
.B(n_1135),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1174),
.B(n_1179),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1243),
.B(n_873),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1216),
.B(n_635),
.C(n_901),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1184),
.Y(n_1378)
);

O2A1O1Ixp33_ASAP7_75t_SL g1379 ( 
.A1(n_1216),
.A2(n_1242),
.B(n_1250),
.C(n_1223),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1177),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1168),
.A2(n_1166),
.B1(n_941),
.B2(n_873),
.Y(n_1381)
);

INVxp33_ASAP7_75t_L g1382 ( 
.A(n_1213),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1304),
.A2(n_1260),
.B(n_1258),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1288),
.B(n_1273),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1348),
.B(n_1294),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1273),
.B(n_1274),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1278),
.B(n_1300),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1292),
.B(n_1358),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1319),
.B(n_1286),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1340),
.A2(n_1381),
.B1(n_1353),
.B2(n_1343),
.Y(n_1390)
);

AND2x6_ASAP7_75t_L g1391 ( 
.A(n_1305),
.B(n_1306),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1279),
.B(n_1318),
.Y(n_1392)
);

O2A1O1Ixp5_ASAP7_75t_L g1393 ( 
.A1(n_1275),
.A2(n_1354),
.B(n_1349),
.C(n_1341),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1340),
.A2(n_1381),
.B1(n_1353),
.B2(n_1263),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1294),
.A2(n_1317),
.B(n_1377),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1271),
.B(n_1382),
.Y(n_1396)
);

AND2x6_ASAP7_75t_L g1397 ( 
.A(n_1305),
.B(n_1306),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1300),
.B(n_1283),
.Y(n_1398)
);

AOI221xp5_ASAP7_75t_L g1399 ( 
.A1(n_1359),
.A2(n_1379),
.B1(n_1365),
.B2(n_1347),
.C(n_1266),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1334),
.A2(n_1347),
.B(n_1365),
.C(n_1359),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1329),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1382),
.B(n_1375),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1265),
.A2(n_1352),
.B(n_1280),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1320),
.B(n_1321),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1339),
.B(n_1342),
.Y(n_1405)
);

BUFx4f_ASAP7_75t_L g1406 ( 
.A(n_1329),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1283),
.B(n_1317),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1284),
.A2(n_1257),
.B(n_1374),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1379),
.A2(n_1277),
.B(n_1338),
.C(n_1376),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1345),
.Y(n_1410)
);

NOR2xp67_ASAP7_75t_L g1411 ( 
.A(n_1312),
.B(n_1324),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_SL g1412 ( 
.A(n_1322),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1338),
.A2(n_1376),
.B1(n_1346),
.B2(n_1363),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1299),
.A2(n_1282),
.B(n_1326),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1303),
.Y(n_1415)
);

NOR2xp67_ASAP7_75t_L g1416 ( 
.A(n_1290),
.B(n_1325),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1362),
.B(n_1366),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1303),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1369),
.A2(n_1326),
.B(n_1299),
.C(n_1328),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1367),
.Y(n_1420)
);

O2A1O1Ixp5_ASAP7_75t_L g1421 ( 
.A1(n_1287),
.A2(n_1330),
.B(n_1361),
.C(n_1310),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1299),
.A2(n_1378),
.B(n_1333),
.C(n_1313),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1301),
.A2(n_1315),
.B1(n_1308),
.B2(n_1293),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1293),
.A2(n_1307),
.B1(n_1333),
.B2(n_1302),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1350),
.A2(n_1372),
.B(n_1357),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1282),
.A2(n_1352),
.B(n_1280),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1262),
.B(n_1314),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1293),
.A2(n_1314),
.B1(n_1352),
.B2(n_1280),
.Y(n_1428)
);

O2A1O1Ixp5_ASAP7_75t_L g1429 ( 
.A1(n_1259),
.A2(n_1380),
.B(n_1368),
.C(n_1360),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1289),
.B(n_1291),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1335),
.A2(n_1311),
.B(n_1295),
.C(n_1332),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1323),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1364),
.A2(n_1267),
.B1(n_1316),
.B2(n_1351),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1345),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1272),
.A2(n_1270),
.B(n_1264),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1336),
.A2(n_1337),
.B(n_1269),
.C(n_1309),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1355),
.A2(n_1269),
.B1(n_1370),
.B2(n_1261),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1373),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1373),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1298),
.A2(n_1268),
.B(n_1281),
.Y(n_1440)
);

NOR2xp67_ASAP7_75t_L g1441 ( 
.A(n_1296),
.B(n_1370),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1331),
.B(n_1285),
.Y(n_1442)
);

O2A1O1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1344),
.A2(n_1360),
.B(n_1368),
.C(n_1285),
.Y(n_1443)
);

CKINVDCx12_ASAP7_75t_R g1444 ( 
.A(n_1344),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1327),
.B(n_1285),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1329),
.Y(n_1446)
);

O2A1O1Ixp5_ASAP7_75t_L g1447 ( 
.A1(n_1275),
.A2(n_1258),
.B(n_1349),
.C(n_1341),
.Y(n_1447)
);

O2A1O1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1371),
.A2(n_1223),
.B(n_1242),
.C(n_1216),
.Y(n_1448)
);

O2A1O1Ixp5_ASAP7_75t_L g1449 ( 
.A1(n_1275),
.A2(n_1258),
.B(n_1349),
.C(n_1341),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1288),
.B(n_1273),
.Y(n_1450)
);

OA21x2_ASAP7_75t_L g1451 ( 
.A1(n_1304),
.A2(n_1260),
.B(n_1258),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1340),
.A2(n_1381),
.B1(n_1353),
.B2(n_873),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1340),
.A2(n_1381),
.B1(n_1353),
.B2(n_873),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1340),
.A2(n_1381),
.B1(n_1353),
.B2(n_873),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1278),
.B(n_1356),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1316),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1348),
.B(n_1274),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1288),
.B(n_1273),
.Y(n_1458)
);

A2O1A1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1371),
.A2(n_1207),
.B(n_1276),
.C(n_1271),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1297),
.B(n_1348),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1297),
.B(n_1348),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1393),
.A2(n_1449),
.B(n_1447),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1445),
.B(n_1442),
.Y(n_1463)
);

BUFx4f_ASAP7_75t_L g1464 ( 
.A(n_1391),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1432),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1445),
.B(n_1430),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1431),
.B(n_1403),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1443),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1440),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1429),
.A2(n_1425),
.B(n_1408),
.Y(n_1470)
);

INVx5_ASAP7_75t_L g1471 ( 
.A(n_1391),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1383),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1391),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1451),
.B(n_1428),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1426),
.B(n_1396),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1397),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1387),
.A2(n_1398),
.B(n_1407),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1425),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1392),
.B(n_1398),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1459),
.A2(n_1387),
.B(n_1448),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1455),
.B(n_1427),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1421),
.B(n_1384),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1435),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1420),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1435),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1395),
.A2(n_1390),
.B(n_1394),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1455),
.B(n_1385),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1404),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1405),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1444),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1417),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1423),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1460),
.B(n_1461),
.Y(n_1493)
);

AO21x2_ASAP7_75t_L g1494 ( 
.A1(n_1390),
.A2(n_1394),
.B(n_1436),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1422),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1450),
.B(n_1458),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1386),
.B(n_1399),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1424),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1424),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1467),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1463),
.B(n_1414),
.Y(n_1501)
);

AO21x2_ASAP7_75t_L g1502 ( 
.A1(n_1470),
.A2(n_1453),
.B(n_1452),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1477),
.B(n_1457),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1463),
.B(n_1402),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1469),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1463),
.B(n_1388),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1477),
.B(n_1487),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1465),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1466),
.B(n_1389),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1466),
.B(n_1438),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1465),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1477),
.B(n_1413),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1477),
.B(n_1413),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1477),
.B(n_1437),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1474),
.B(n_1439),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1467),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1483),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1474),
.B(n_1400),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1483),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1474),
.B(n_1419),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1486),
.A2(n_1454),
.B1(n_1452),
.B2(n_1453),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1487),
.B(n_1409),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1485),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1517),
.A2(n_1470),
.B(n_1472),
.Y(n_1524)
);

AOI33xp33_ASAP7_75t_L g1525 ( 
.A1(n_1521),
.A2(n_1482),
.A3(n_1497),
.B1(n_1498),
.B2(n_1499),
.B3(n_1495),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1515),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1515),
.Y(n_1527)
);

OAI21xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1513),
.A2(n_1476),
.B(n_1495),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1521),
.A2(n_1486),
.B1(n_1480),
.B2(n_1494),
.Y(n_1529)
);

AOI221xp5_ASAP7_75t_L g1530 ( 
.A1(n_1522),
.A2(n_1462),
.B1(n_1454),
.B2(n_1486),
.C(n_1480),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1502),
.A2(n_1486),
.B1(n_1480),
.B2(n_1494),
.Y(n_1531)
);

INVx4_ASAP7_75t_L g1532 ( 
.A(n_1500),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1522),
.B(n_1493),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1503),
.B(n_1482),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1512),
.A2(n_1464),
.B1(n_1495),
.B2(n_1433),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1500),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1501),
.B(n_1475),
.Y(n_1537)
);

NOR3xp33_ASAP7_75t_SL g1538 ( 
.A(n_1513),
.B(n_1446),
.C(n_1401),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1507),
.B(n_1481),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1515),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1500),
.B(n_1471),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1508),
.Y(n_1542)
);

OA222x2_ASAP7_75t_L g1543 ( 
.A1(n_1513),
.A2(n_1499),
.B1(n_1498),
.B2(n_1479),
.C1(n_1492),
.C2(n_1481),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1512),
.A2(n_1464),
.B1(n_1433),
.B2(n_1479),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1502),
.A2(n_1486),
.B1(n_1480),
.B2(n_1494),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1508),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1504),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1502),
.A2(n_1480),
.B1(n_1494),
.B2(n_1475),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1508),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1510),
.Y(n_1550)
);

OR2x6_ASAP7_75t_L g1551 ( 
.A(n_1500),
.B(n_1476),
.Y(n_1551)
);

OAI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1500),
.A2(n_1462),
.B1(n_1481),
.B2(n_1493),
.C(n_1416),
.Y(n_1552)
);

OAI33xp33_ASAP7_75t_L g1553 ( 
.A1(n_1507),
.A2(n_1468),
.A3(n_1479),
.B1(n_1484),
.B2(n_1488),
.B3(n_1491),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_1504),
.Y(n_1554)
);

OAI33xp33_ASAP7_75t_L g1555 ( 
.A1(n_1503),
.A2(n_1468),
.A3(n_1484),
.B1(n_1489),
.B2(n_1491),
.B3(n_1488),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1500),
.B(n_1471),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1505),
.A2(n_1478),
.B(n_1472),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1511),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1503),
.B(n_1482),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1501),
.B(n_1475),
.Y(n_1560)
);

NAND4xp25_ASAP7_75t_L g1561 ( 
.A(n_1518),
.B(n_1411),
.C(n_1499),
.D(n_1498),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1533),
.B(n_1520),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1539),
.B(n_1503),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1534),
.B(n_1514),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1557),
.A2(n_1523),
.B(n_1519),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1524),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1524),
.Y(n_1567)
);

INVxp67_ASAP7_75t_L g1568 ( 
.A(n_1561),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1542),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1542),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1552),
.B(n_1406),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1546),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1534),
.B(n_1559),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1546),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_L g1575 ( 
.A(n_1530),
.B(n_1520),
.C(n_1518),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1549),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1551),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1537),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1537),
.B(n_1501),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1559),
.B(n_1514),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1549),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1558),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1551),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1551),
.Y(n_1584)
);

INVx4_ASAP7_75t_SL g1585 ( 
.A(n_1551),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1525),
.B(n_1520),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1535),
.B(n_1464),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1560),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1544),
.B(n_1464),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1560),
.B(n_1526),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1547),
.B(n_1514),
.Y(n_1591)
);

AOI211xp5_ASAP7_75t_L g1592 ( 
.A1(n_1575),
.A2(n_1568),
.B(n_1571),
.C(n_1587),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1585),
.B(n_1543),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1565),
.Y(n_1594)
);

NAND4xp25_ASAP7_75t_SL g1595 ( 
.A(n_1586),
.B(n_1531),
.C(n_1545),
.D(n_1529),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1585),
.B(n_1543),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1591),
.B(n_1573),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1585),
.B(n_1532),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1591),
.B(n_1554),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1585),
.B(n_1532),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1562),
.B(n_1527),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1585),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1579),
.B(n_1532),
.Y(n_1603)
);

NAND2xp33_ASAP7_75t_R g1604 ( 
.A(n_1577),
.B(n_1410),
.Y(n_1604)
);

CKINVDCx16_ASAP7_75t_R g1605 ( 
.A(n_1577),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1579),
.B(n_1536),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1569),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1565),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1569),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1589),
.B(n_1406),
.Y(n_1610)
);

NAND2x1p5_ASAP7_75t_L g1611 ( 
.A(n_1583),
.B(n_1471),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1583),
.B(n_1536),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1570),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1570),
.B(n_1572),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1572),
.B(n_1540),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1584),
.B(n_1536),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1574),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1584),
.B(n_1541),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1565),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1574),
.B(n_1541),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1576),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1576),
.B(n_1541),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1578),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1590),
.B(n_1556),
.Y(n_1624)
);

NAND4xp25_ASAP7_75t_L g1625 ( 
.A(n_1564),
.B(n_1548),
.C(n_1561),
.D(n_1520),
.Y(n_1625)
);

NAND5xp2_ASAP7_75t_L g1626 ( 
.A(n_1590),
.B(n_1538),
.C(n_1518),
.D(n_1497),
.E(n_1412),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1588),
.B(n_1556),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1565),
.Y(n_1628)
);

AND2x2_ASAP7_75t_SL g1629 ( 
.A(n_1573),
.B(n_1464),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1581),
.B(n_1556),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1580),
.B(n_1528),
.C(n_1518),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1581),
.B(n_1500),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1582),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1633),
.Y(n_1634)
);

XOR2x2_ASAP7_75t_L g1635 ( 
.A(n_1592),
.B(n_1494),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1633),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1629),
.B(n_1580),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1592),
.B(n_1509),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_SL g1639 ( 
.A(n_1593),
.B(n_1514),
.C(n_1490),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1605),
.B(n_1509),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1607),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1629),
.B(n_1563),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1607),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1604),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1623),
.B(n_1563),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1609),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1595),
.B(n_1434),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1609),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1613),
.Y(n_1649)
);

NOR2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1625),
.B(n_1473),
.Y(n_1650)
);

O2A1O1Ixp33_ASAP7_75t_L g1651 ( 
.A1(n_1625),
.A2(n_1528),
.B(n_1553),
.C(n_1555),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1605),
.B(n_1509),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1623),
.B(n_1509),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1620),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1601),
.B(n_1550),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1613),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1618),
.B(n_1506),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1618),
.B(n_1506),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1617),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1617),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1602),
.B(n_1506),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1593),
.A2(n_1490),
.B(n_1501),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1602),
.B(n_1506),
.Y(n_1663)
);

NAND2x1p5_ASAP7_75t_L g1664 ( 
.A(n_1629),
.B(n_1471),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1621),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1596),
.B(n_1496),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1621),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1610),
.B(n_1456),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1598),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1654),
.B(n_1596),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1644),
.B(n_1631),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1669),
.B(n_1598),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1635),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1635),
.B(n_1634),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1636),
.B(n_1601),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1656),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1669),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1654),
.B(n_1600),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1647),
.A2(n_1626),
.B1(n_1502),
.B2(n_1631),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1656),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1666),
.B(n_1597),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1647),
.B(n_1620),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1637),
.B(n_1600),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1668),
.B(n_1626),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1668),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1637),
.B(n_1642),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1664),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1642),
.B(n_1624),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1638),
.B(n_1614),
.Y(n_1689)
);

CKINVDCx14_ASAP7_75t_R g1690 ( 
.A(n_1639),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1650),
.B(n_1624),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1640),
.B(n_1620),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_1645),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1657),
.B(n_1597),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1662),
.B(n_1612),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1693),
.B(n_1652),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1690),
.A2(n_1651),
.B1(n_1664),
.B2(n_1661),
.Y(n_1697)
);

OAI31xp33_ASAP7_75t_L g1698 ( 
.A1(n_1673),
.A2(n_1611),
.A3(n_1616),
.B(n_1612),
.Y(n_1698)
);

OAI21xp33_ASAP7_75t_L g1699 ( 
.A1(n_1673),
.A2(n_1663),
.B(n_1653),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1680),
.Y(n_1700)
);

NOR2xp67_ASAP7_75t_SL g1701 ( 
.A(n_1685),
.B(n_1415),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_SL g1702 ( 
.A(n_1673),
.B(n_1611),
.C(n_1616),
.Y(n_1702)
);

AOI21xp33_ASAP7_75t_L g1703 ( 
.A1(n_1693),
.A2(n_1643),
.B(n_1641),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1671),
.A2(n_1627),
.B1(n_1658),
.B2(n_1502),
.Y(n_1704)
);

OAI21xp5_ASAP7_75t_SL g1705 ( 
.A1(n_1679),
.A2(n_1611),
.B(n_1627),
.Y(n_1705)
);

AOI21xp33_ASAP7_75t_L g1706 ( 
.A1(n_1674),
.A2(n_1685),
.B(n_1684),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1686),
.B(n_1603),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1672),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1674),
.A2(n_1667),
.B1(n_1665),
.B2(n_1646),
.C(n_1648),
.Y(n_1709)
);

AOI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1677),
.A2(n_1660),
.B1(n_1659),
.B2(n_1649),
.C(n_1632),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1686),
.Y(n_1711)
);

NOR2x1_ASAP7_75t_L g1712 ( 
.A(n_1685),
.B(n_1614),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1688),
.A2(n_1502),
.B1(n_1516),
.B2(n_1500),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1682),
.B(n_1655),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1688),
.A2(n_1516),
.B1(n_1500),
.B2(n_1622),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1680),
.Y(n_1716)
);

AND2x2_ASAP7_75t_SL g1717 ( 
.A(n_1714),
.B(n_1696),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1708),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1706),
.A2(n_1695),
.B1(n_1683),
.B2(n_1675),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1711),
.B(n_1683),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1712),
.B(n_1676),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1707),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1700),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1716),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1697),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1699),
.B(n_1675),
.Y(n_1726)
);

OAI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1719),
.A2(n_1721),
.B1(n_1726),
.B2(n_1725),
.C(n_1709),
.Y(n_1727)
);

OAI211xp5_ASAP7_75t_L g1728 ( 
.A1(n_1719),
.A2(n_1703),
.B(n_1705),
.C(n_1698),
.Y(n_1728)
);

OAI21xp5_ASAP7_75t_SL g1729 ( 
.A1(n_1720),
.A2(n_1702),
.B(n_1698),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1721),
.Y(n_1730)
);

OAI211xp5_ASAP7_75t_L g1731 ( 
.A1(n_1720),
.A2(n_1710),
.B(n_1704),
.C(n_1676),
.Y(n_1731)
);

AND5x1_ASAP7_75t_L g1732 ( 
.A(n_1717),
.B(n_1683),
.C(n_1670),
.D(n_1678),
.E(n_1672),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1722),
.B(n_1683),
.Y(n_1733)
);

O2A1O1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1718),
.A2(n_1680),
.B(n_1689),
.C(n_1695),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1723),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1727),
.A2(n_1728),
.B1(n_1729),
.B2(n_1681),
.Y(n_1736)
);

NOR4xp25_ASAP7_75t_L g1737 ( 
.A(n_1727),
.B(n_1724),
.C(n_1670),
.D(n_1689),
.Y(n_1737)
);

A2O1A1Ixp33_ASAP7_75t_L g1738 ( 
.A1(n_1734),
.A2(n_1701),
.B(n_1672),
.C(n_1687),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1733),
.Y(n_1739)
);

AND5x1_ASAP7_75t_L g1740 ( 
.A(n_1732),
.B(n_1672),
.C(n_1678),
.D(n_1687),
.E(n_1715),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1739),
.B(n_1730),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_SL g1742 ( 
.A(n_1738),
.B(n_1735),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1737),
.B(n_1691),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1736),
.A2(n_1731),
.B1(n_1678),
.B2(n_1713),
.C(n_1691),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1740),
.B(n_1678),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1739),
.B(n_1692),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1746),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1742),
.A2(n_1681),
.B1(n_1694),
.B2(n_1620),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1745),
.A2(n_1694),
.B1(n_1630),
.B2(n_1622),
.Y(n_1749)
);

CKINVDCx20_ASAP7_75t_R g1750 ( 
.A(n_1741),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1743),
.A2(n_1630),
.B(n_1622),
.Y(n_1751)
);

AND4x2_ASAP7_75t_L g1752 ( 
.A(n_1751),
.B(n_1744),
.C(n_1594),
.D(n_1622),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1747),
.B(n_1750),
.Y(n_1753)
);

BUFx4f_ASAP7_75t_SL g1754 ( 
.A(n_1749),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1753),
.B(n_1748),
.Y(n_1755)
);

OAI322xp33_ASAP7_75t_L g1756 ( 
.A1(n_1755),
.A2(n_1752),
.A3(n_1754),
.B1(n_1594),
.B2(n_1608),
.C1(n_1619),
.C2(n_1628),
.Y(n_1756)
);

OA22x2_ASAP7_75t_L g1757 ( 
.A1(n_1756),
.A2(n_1608),
.B1(n_1619),
.B2(n_1628),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1756),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1758),
.B(n_1630),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1757),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1759),
.Y(n_1761)
);

CKINVDCx20_ASAP7_75t_R g1762 ( 
.A(n_1760),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_SL g1763 ( 
.A1(n_1761),
.A2(n_1418),
.B(n_1415),
.Y(n_1763)
);

AOI222xp33_ASAP7_75t_L g1764 ( 
.A1(n_1762),
.A2(n_1594),
.B1(n_1608),
.B2(n_1628),
.C1(n_1619),
.C2(n_1630),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1763),
.A2(n_1764),
.B(n_1594),
.Y(n_1765)
);

OAI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1603),
.B(n_1606),
.Y(n_1766)
);

AOI22x1_ASAP7_75t_L g1767 ( 
.A1(n_1766),
.A2(n_1415),
.B1(n_1599),
.B2(n_1606),
.Y(n_1767)
);

AOI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1767),
.A2(n_1632),
.B1(n_1615),
.B2(n_1566),
.C(n_1567),
.Y(n_1768)
);

AOI211xp5_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1441),
.B(n_1599),
.C(n_1632),
.Y(n_1769)
);


endmodule