module real_jpeg_17833_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_475),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_0),
.B(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_1),
.Y(n_476)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_2),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_2),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_2),
.B(n_141),
.Y(n_140)
);

NAND2x1p5_ASAP7_75t_L g189 ( 
.A(n_2),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_2),
.B(n_137),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_2),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_2),
.B(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_3),
.Y(n_165)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_3),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_4),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g391 ( 
.A(n_4),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_5),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_5),
.A2(n_11),
.B1(n_115),
.B2(n_119),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_5),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_5),
.B(n_55),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_5),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_5),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_5),
.B(n_456),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_6),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_6),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_6),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_6),
.B(n_90),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_6),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_6),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_6),
.B(n_459),
.Y(n_458)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_7),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_7),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_7),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_8),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_8),
.Y(n_168)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_8),
.Y(n_268)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_8),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_9),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_9),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_9),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_9),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_9),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_9),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_9),
.B(n_372),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_10),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_10),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_10),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_10),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_10),
.B(n_345),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_10),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_10),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_10),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_11),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_11),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_11),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_11),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_11),
.B(n_406),
.Y(n_405)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_12),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_12),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_13),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_13),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_13),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_13),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_13),
.B(n_90),
.Y(n_264)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_13),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_14),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_15),
.Y(n_87)
);

BUFx4f_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_15),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_16),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_16),
.B(n_76),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_16),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_16),
.B(n_350),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_SL g387 ( 
.A(n_16),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_16),
.B(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_16),
.B(n_420),
.Y(n_419)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_17),
.Y(n_103)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_17),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_17),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_442),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2x1_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_436),
.Y(n_21)
);

NAND4xp25_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_224),
.C(n_307),
.D(n_312),
.Y(n_22)
);

NOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_173),
.Y(n_23)
);

NOR2xp67_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_147),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_25),
.B(n_147),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_98),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_26),
.B(n_99),
.C(n_124),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_66),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_46),
.Y(n_27)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_28),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_31),
.B(n_40),
.C(n_41),
.Y(n_223)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_41),
.A2(n_42),
.B1(n_294),
.B2(n_298),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_42),
.B(n_291),
.C(n_298),
.Y(n_470)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_46),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_57),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B1(n_52),
.B2(n_56),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_48),
.A2(n_52),
.B(n_57),
.C(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_50),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_51),
.B(n_56),
.Y(n_199)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_54),
.Y(n_416)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.C(n_62),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_58),
.A2(n_62),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_58),
.A2(n_95),
.B1(n_127),
.B2(n_158),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_60),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_62),
.B(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_65),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_66),
.B(n_177),
.C(n_178),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_79),
.C(n_88),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_67),
.B(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_71),
.C(n_75),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_79),
.A2(n_80),
.B1(n_88),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g429 ( 
.A(n_83),
.Y(n_429)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_84),
.A2(n_160),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_86),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_87),
.Y(n_425)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.C(n_95),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_89),
.A2(n_95),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_89),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_91),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_92),
.B(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_94),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_95),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_95),
.A2(n_140),
.B1(n_158),
.B2(n_258),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_95),
.B(n_258),
.C(n_301),
.Y(n_471)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_97),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_124),
.Y(n_98)
);

XOR2x2_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_114),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_113),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_101),
.B(n_183),
.C(n_184),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_102),
.B(n_106),
.C(n_109),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_112),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_109),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

XNOR2x1_ASAP7_75t_SL g321 ( 
.A(n_112),
.B(n_140),
.Y(n_321)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_130),
.B(n_133),
.Y(n_129)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g407 ( 
.A(n_117),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_122),
.Y(n_457)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_123),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.C(n_138),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_129),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_128),
.B(n_263),
.C(n_269),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_131),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.C(n_145),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_139),
.B(n_319),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_140),
.A2(n_221),
.B1(n_222),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_140),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_140),
.B(n_222),
.C(n_253),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_319)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_154),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_148),
.B(n_335),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_154),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.C(n_161),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_155),
.B(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_159),
.B(n_161),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_160),
.B(n_215),
.C(n_222),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.C(n_169),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_162),
.B(n_169),
.Y(n_359)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_166),
.B(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21x1_ASAP7_75t_SL g437 ( 
.A1(n_173),
.A2(n_438),
.B(n_439),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_174),
.B(n_175),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_176),
.B(n_180),
.C(n_203),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_202),
.B2(n_203),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_196),
.B2(n_197),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_188)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_195),
.C(n_197),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_196),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_249),
.C(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_213),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_223),
.C(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_208),
.C(n_212),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_212),
.Y(n_207)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_210),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_211),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_212),
.A2(n_453),
.B1(n_454),
.B2(n_455),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_212),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_223),
.Y(n_213)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_217),
.Y(n_459)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_221),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_221),
.B(n_329),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_222),
.B(n_329),
.Y(n_328)
);

A2O1A1O1Ixp25_ASAP7_75t_L g436 ( 
.A1(n_224),
.A2(n_307),
.B(n_437),
.C(n_440),
.D(n_441),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_270),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_225),
.B(n_270),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_247),
.C(n_251),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_226),
.A2(n_227),
.B1(n_251),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_246),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_232),
.C(n_245),
.Y(n_271)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_245),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_234),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_244),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_240),
.B2(n_241),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_240),
.C(n_244),
.Y(n_277)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_241),
.B(n_285),
.C(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_248),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_251),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_259),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_260),
.C(n_261),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_269),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_271),
.B(n_273),
.C(n_473),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_287),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_286),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_274),
.B(n_277),
.C(n_278),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_276),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

AO22x1_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_278)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_280),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_283),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_287),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_299),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_289),
.B(n_290),
.C(n_299),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_294),
.Y(n_298)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_302),
.B(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_308),
.B(n_309),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_337),
.B(n_435),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_334),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_314),
.B(n_334),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.C(n_320),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_315),
.A2(n_316),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_318),
.B(n_320),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.C(n_328),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_328),
.B(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_333),
.Y(n_404)
);

AOI21x1_ASAP7_75t_SL g337 ( 
.A1(n_338),
.A2(n_363),
.B(n_434),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_360),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_339),
.B(n_360),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.C(n_358),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_358),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_349),
.C(n_355),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_368),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_355),
.Y(n_368)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

OAI21x1_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_382),
.B(n_433),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_380),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_365),
.B(n_380),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_369),
.C(n_378),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_366),
.A2(n_367),
.B1(n_393),
.B2(n_395),
.Y(n_392)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_369),
.A2(n_378),
.B1(n_379),
.B2(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_369),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_375),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_370),
.A2(n_371),
.B1(n_375),
.B2(n_376),
.Y(n_385)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_396),
.B(n_432),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_392),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_384),
.B(n_392),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.C(n_390),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_409),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_386),
.A2(n_387),
.B1(n_390),
.B2(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_390),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_393),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_397),
.A2(n_411),
.B(n_431),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_408),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_398),
.B(n_408),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_405),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_405),
.Y(n_417)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_418),
.B(n_430),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_417),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_413),
.B(n_417),
.Y(n_430)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_426),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_474),
.Y(n_442)
);

OR2x2_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_472),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_472),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_463),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_461),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_452),
.B1(n_458),
.B2(n_460),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx8_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_458),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_469),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);


endmodule