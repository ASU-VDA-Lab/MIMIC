module fake_jpeg_16463_n_116 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_116);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

AOI21xp33_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_0),
.B(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_26),
.B(n_15),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_16),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_20),
.B1(n_14),
.B2(n_25),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_13),
.B1(n_18),
.B2(n_19),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_16),
.B1(n_14),
.B2(n_25),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_23),
.B1(n_22),
.B2(n_21),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_54),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_34),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_16),
.B(n_19),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_56),
.C(n_12),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_17),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_13),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_58),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_27),
.C(n_31),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_43),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_71),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_55),
.B1(n_53),
.B2(n_30),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_0),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_57),
.B(n_50),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_54),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_60),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_83),
.B(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_56),
.B1(n_51),
.B2(n_46),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_84),
.B1(n_65),
.B2(n_61),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_48),
.C(n_49),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_80),
.C(n_81),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_64),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_73),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_27),
.C(n_59),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_39),
.B(n_59),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_76),
.B1(n_87),
.B2(n_77),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_92),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_65),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_93),
.C(n_82),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_73),
.B1(n_63),
.B2(n_70),
.C(n_62),
.Y(n_91)
);

A2O1A1O1Ixp25_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_81),
.B(n_84),
.C(n_83),
.D(n_72),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_63),
.C(n_18),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_72),
.C(n_27),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_99),
.Y(n_101)
);

AOI321xp33_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_90),
.A3(n_39),
.B1(n_24),
.B2(n_27),
.C(n_28),
.Y(n_103)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_93),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_28),
.C(n_39),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_21),
.B1(n_22),
.B2(n_29),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_104),
.Y(n_106)
);

AOI221xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_99),
.B1(n_98),
.B2(n_24),
.C(n_4),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_39),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_100),
.A3(n_101),
.B1(n_96),
.B2(n_94),
.C1(n_104),
.C2(n_95),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_24),
.C(n_3),
.Y(n_111)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_109),
.C(n_0),
.Y(n_112)
);

AOI322xp5_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_10),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_10),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_6),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_114),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_7),
.Y(n_116)
);


endmodule