module fake_jpeg_31980_n_540 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_540);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_540;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_58),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_19),
.B(n_10),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_63),
.Y(n_107)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_62),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_64),
.B(n_75),
.Y(n_116)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_27),
.B(n_18),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_76),
.B(n_77),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_27),
.B(n_9),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_19),
.B(n_9),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_39),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

CKINVDCx6p67_ASAP7_75t_R g109 ( 
.A(n_83),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_87),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_31),
.B(n_9),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_31),
.B(n_17),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_89),
.B(n_91),
.Y(n_147)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_42),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_35),
.B(n_7),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_92),
.B(n_93),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_42),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_35),
.B(n_7),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_95),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_101),
.Y(n_138)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_102),
.B(n_51),
.Y(n_150)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_103),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_104),
.B(n_145),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_86),
.A2(n_88),
.B1(n_90),
.B2(n_59),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_111),
.A2(n_118),
.B1(n_37),
.B2(n_40),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_39),
.B1(n_50),
.B2(n_49),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_119),
.B(n_120),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_83),
.B(n_23),
.Y(n_120)
);

BUFx16f_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

CKINVDCx6p67_ASAP7_75t_R g213 ( 
.A(n_125),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

CKINVDCx6p67_ASAP7_75t_R g226 ( 
.A(n_127),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_79),
.A2(n_23),
.B(n_50),
.C(n_49),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_131),
.B(n_132),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_74),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_55),
.B(n_51),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_150),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

NAND2x1p5_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_36),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_84),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_164),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx3_ASAP7_75t_SL g189 ( 
.A(n_155),
.Y(n_189)
);

BUFx12_ASAP7_75t_L g160 ( 
.A(n_53),
.Y(n_160)
);

CKINVDCx12_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_56),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_162),
.Y(n_224)
);

BUFx12_ASAP7_75t_L g163 ( 
.A(n_58),
.Y(n_163)
);

CKINVDCx12_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_62),
.B(n_33),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_168),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_124),
.A2(n_78),
.B1(n_73),
.B2(n_97),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_171),
.A2(n_151),
.B1(n_110),
.B2(n_139),
.Y(n_247)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_172),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_173),
.A2(n_176),
.B1(n_199),
.B2(n_223),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_116),
.B(n_33),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_174),
.B(n_179),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_38),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_175),
.B(n_202),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_70),
.B1(n_69),
.B2(n_66),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_177),
.Y(n_261)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_116),
.B(n_38),
.Y(n_179)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_182),
.Y(n_259)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_183),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_20),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_185),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_43),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_186),
.Y(n_244)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_112),
.B(n_68),
.C(n_65),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_193),
.Y(n_239)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_108),
.Y(n_191)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_191),
.Y(n_269)
);

BUFx12_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_194),
.Y(n_268)
);

CKINVDCx12_ASAP7_75t_R g195 ( 
.A(n_109),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_109),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_197),
.B(n_204),
.Y(n_258)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_198),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_107),
.A2(n_71),
.B1(n_57),
.B2(n_37),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_43),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_142),
.B(n_41),
.C(n_40),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_109),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_205),
.B(n_212),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_142),
.B(n_41),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_210),
.Y(n_242)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_208),
.Y(n_274)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_209),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_136),
.B(n_29),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_211),
.Y(n_240)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_216),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_136),
.B(n_29),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_138),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_115),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_115),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_217),
.B(n_218),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_137),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_111),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_148),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_225),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_152),
.B(n_36),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_221),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_222),
.A2(n_129),
.B1(n_127),
.B2(n_155),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_107),
.A2(n_26),
.B1(n_36),
.B2(n_11),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_137),
.Y(n_225)
);

NAND2xp33_ASAP7_75t_SL g227 ( 
.A(n_145),
.B(n_36),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_227),
.B(n_45),
.Y(n_275)
);

AO22x1_ASAP7_75t_SL g229 ( 
.A1(n_227),
.A2(n_161),
.B1(n_156),
.B2(n_154),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_229),
.B(n_249),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_231),
.A2(n_276),
.B1(n_189),
.B2(n_226),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_213),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_237),
.B(n_245),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_170),
.A2(n_161),
.B1(n_130),
.B2(n_152),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_243),
.A2(n_247),
.B1(n_252),
.B2(n_257),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_213),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_248),
.B(n_263),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_162),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_L g252 ( 
.A1(n_190),
.A2(n_144),
.B1(n_158),
.B2(n_114),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_169),
.A2(n_134),
.B1(n_141),
.B2(n_114),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_256),
.A2(n_167),
.B1(n_182),
.B2(n_45),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_200),
.A2(n_138),
.B1(n_139),
.B2(n_36),
.Y(n_257)
);

AO22x2_ASAP7_75t_L g260 ( 
.A1(n_206),
.A2(n_26),
.B1(n_160),
.B2(n_163),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_260),
.B(n_267),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_213),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_171),
.A2(n_198),
.B1(n_201),
.B2(n_211),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_265),
.A2(n_266),
.B1(n_12),
.B2(n_16),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_196),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_204),
.B(n_0),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_224),
.B(n_187),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_270),
.A2(n_271),
.B(n_275),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_224),
.B(n_0),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_214),
.A2(n_177),
.B1(n_194),
.B2(n_178),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_172),
.B(n_0),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_1),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_239),
.A2(n_226),
.B(n_168),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_282),
.A2(n_314),
.B(n_290),
.Y(n_344)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_283),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_284),
.B(n_325),
.Y(n_347)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_238),
.B(n_193),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_286),
.B(n_287),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_193),
.Y(n_287)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_230),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_192),
.C(n_226),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_289),
.B(n_297),
.Y(n_328)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_249),
.A2(n_181),
.B(n_191),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_293),
.A2(n_271),
.B(n_267),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_235),
.A2(n_222),
.B1(n_212),
.B2(n_209),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_294),
.A2(n_316),
.B1(n_252),
.B2(n_265),
.Y(n_330)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_295),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_296),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_232),
.B(n_188),
.C(n_180),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_255),
.Y(n_299)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_299),
.Y(n_358)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_244),
.Y(n_300)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_300),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_301),
.Y(n_362)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_244),
.Y(n_302)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_302),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_279),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_303),
.B(n_306),
.Y(n_345)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_274),
.Y(n_304)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_304),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_246),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_232),
.B(n_188),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_307),
.B(n_309),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_248),
.B(n_180),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_274),
.Y(n_310)
);

NAND2xp33_ASAP7_75t_SL g361 ( 
.A(n_310),
.B(n_313),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_246),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_312),
.Y(n_333)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_264),
.Y(n_313)
);

AND2x6_ASAP7_75t_L g314 ( 
.A(n_260),
.B(n_189),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_315),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_235),
.A2(n_229),
.B1(n_243),
.B2(n_260),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_242),
.B(n_45),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_317),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_242),
.B(n_45),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_318),
.Y(n_351)
);

BUFx12_ASAP7_75t_L g320 ( 
.A(n_259),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_320),
.Y(n_365)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_253),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_321),
.Y(n_348)
);

OAI21xp33_ASAP7_75t_SL g360 ( 
.A1(n_322),
.A2(n_324),
.B(n_269),
.Y(n_360)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_253),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_323),
.Y(n_352)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_237),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_240),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_327),
.A2(n_273),
.B1(n_262),
.B2(n_278),
.Y(n_346)
);

AO21x1_ASAP7_75t_L g392 ( 
.A1(n_329),
.A2(n_336),
.B(n_344),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_330),
.A2(n_346),
.B1(n_360),
.B2(n_297),
.Y(n_370)
);

XNOR2x2_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_260),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_281),
.A2(n_228),
.B1(n_229),
.B2(n_260),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_337),
.A2(n_354),
.B1(n_293),
.B2(n_319),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_289),
.B(n_236),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_338),
.B(n_273),
.C(n_310),
.Y(n_381)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_236),
.C(n_258),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_341),
.B(n_311),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_290),
.A2(n_228),
.B1(n_277),
.B2(n_278),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_357),
.Y(n_375)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_353),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_298),
.A2(n_259),
.B1(n_234),
.B2(n_250),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_298),
.A2(n_241),
.B1(n_250),
.B2(n_230),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_308),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_364),
.B(n_282),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_370),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_371),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_372),
.B(n_338),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_345),
.B(n_302),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_374),
.B(n_386),
.Y(n_406)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_353),
.Y(n_376)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_335),
.Y(n_377)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_377),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_334),
.A2(n_327),
.B1(n_311),
.B2(n_314),
.Y(n_378)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_378),
.Y(n_418)
);

OA22x2_ASAP7_75t_L g379 ( 
.A1(n_337),
.A2(n_324),
.B1(n_300),
.B2(n_283),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_379),
.B(n_383),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_332),
.B(n_285),
.Y(n_380)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_380),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_381),
.B(n_385),
.C(n_396),
.Y(n_421)
);

INVx13_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_387),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_334),
.A2(n_304),
.B1(n_299),
.B2(n_291),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_331),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_384),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_292),
.C(n_295),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_333),
.B(n_326),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_362),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_336),
.A2(n_325),
.B(n_288),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_388),
.Y(n_422)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_335),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_389),
.Y(n_405)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_339),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_390),
.Y(n_423)
);

NOR2x1p5_ASAP7_75t_L g391 ( 
.A(n_342),
.B(n_332),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_391),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_320),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_393),
.B(n_394),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_363),
.B(n_11),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_330),
.A2(n_301),
.B1(n_315),
.B2(n_296),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_395),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_328),
.B(n_269),
.C(n_251),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_339),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_398),
.Y(n_409)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_359),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_341),
.B(n_15),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_399),
.B(n_401),
.Y(n_428)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_400),
.B(n_402),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_347),
.B(n_320),
.Y(n_401)
);

INVx8_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_347),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_367),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_375),
.A2(n_344),
.B(n_350),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_412),
.A2(n_392),
.B(n_393),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g414 ( 
.A1(n_384),
.A2(n_340),
.B1(n_362),
.B2(n_366),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_414),
.A2(n_343),
.B1(n_387),
.B2(n_367),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_429),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_351),
.C(n_350),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_381),
.C(n_380),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_373),
.B(n_351),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_427),
.B(n_431),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_372),
.B(n_329),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_385),
.B(n_361),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_432),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_373),
.B(n_366),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_392),
.B(n_354),
.Y(n_432)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_433),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_391),
.A2(n_357),
.B1(n_349),
.B2(n_358),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_434),
.A2(n_369),
.B1(n_376),
.B2(n_391),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_427),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_435),
.B(n_446),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_437),
.B(n_445),
.Y(n_467)
);

OAI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_419),
.A2(n_402),
.B1(n_400),
.B2(n_398),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_438),
.A2(n_448),
.B1(n_450),
.B2(n_453),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_456),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_422),
.A2(n_388),
.B(n_375),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_440),
.Y(n_480)
);

AO22x1_ASAP7_75t_SL g441 ( 
.A1(n_426),
.A2(n_379),
.B1(n_388),
.B2(n_389),
.Y(n_441)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_441),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_442),
.B(n_425),
.C(n_430),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_379),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_451),
.Y(n_474)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_431),
.Y(n_444)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_444),
.Y(n_468)
);

BUFx24_ASAP7_75t_SL g445 ( 
.A(n_410),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_416),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_410),
.A2(n_397),
.B1(n_390),
.B2(n_377),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_406),
.B(n_382),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_449),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_421),
.B(n_379),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_409),
.Y(n_452)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_452),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_418),
.A2(n_358),
.B1(n_356),
.B2(n_355),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_418),
.A2(n_356),
.B1(n_355),
.B2(n_349),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_455),
.Y(n_475)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_426),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_419),
.A2(n_365),
.B1(n_352),
.B2(n_348),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_411),
.A2(n_323),
.B1(n_321),
.B2(n_251),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_434),
.Y(n_469)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_413),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_459),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_458),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_463),
.B(n_473),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_460),
.Y(n_464)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_464),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_469),
.A2(n_465),
.B1(n_461),
.B2(n_475),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_415),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_476),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_436),
.B(n_429),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_442),
.B(n_412),
.C(n_411),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_478),
.B(n_447),
.C(n_432),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_443),
.B(n_428),
.C(n_420),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_454),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_447),
.B(n_451),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_481),
.B(n_472),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_480),
.A2(n_422),
.B1(n_437),
.B2(n_440),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_482),
.A2(n_495),
.B1(n_498),
.B2(n_469),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_483),
.B(n_487),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_471),
.B(n_446),
.Y(n_484)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_484),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_480),
.A2(n_424),
.B(n_417),
.Y(n_485)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_485),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_468),
.B(n_404),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_488),
.B(n_497),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_462),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_491),
.Y(n_507)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_470),
.Y(n_490)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_490),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_478),
.B(n_456),
.C(n_417),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_492),
.B(n_474),
.C(n_473),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_477),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_461),
.A2(n_457),
.B1(n_404),
.B2(n_441),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_496),
.B(n_441),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_466),
.A2(n_424),
.B1(n_405),
.B2(n_423),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_499),
.B(n_512),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_488),
.Y(n_518)
);

NOR2x1_ASAP7_75t_SL g503 ( 
.A(n_493),
.B(n_467),
.Y(n_503)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_503),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_481),
.C(n_476),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_494),
.C(n_497),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_508),
.B(n_492),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_484),
.A2(n_407),
.B(n_408),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_509),
.A2(n_485),
.B(n_496),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_SL g510 ( 
.A1(n_495),
.A2(n_413),
.B1(n_407),
.B2(n_423),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_510),
.A2(n_12),
.B1(n_13),
.B2(n_5),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_482),
.B(n_405),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_507),
.B(n_486),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_514),
.B(n_520),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_517),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_516),
.B(n_518),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_500),
.B(n_494),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_45),
.C(n_6),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_521),
.A2(n_510),
.B(n_502),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_506),
.B(n_512),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_523),
.B(n_526),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_519),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_513),
.A2(n_505),
.B(n_504),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_530),
.B(n_532),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_516),
.C(n_511),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_531),
.B(n_527),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_527),
.A2(n_518),
.B1(n_501),
.B2(n_511),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_534),
.A2(n_529),
.B(n_531),
.Y(n_535)
);

A2O1A1Ixp33_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_533),
.B(n_528),
.C(n_521),
.Y(n_536)
);

AO21x1_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_12),
.B(n_4),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_537),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_3),
.B(n_5),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_3),
.Y(n_540)
);


endmodule