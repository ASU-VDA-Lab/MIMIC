module fake_jpeg_13033_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx2_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVxp67_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx24_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx2_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_18),
.Y(n_26)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_11),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_21),
.B1(n_22),
.B2(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_23),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_8),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_9),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_9),
.B1(n_12),
.B2(n_15),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_18),
.B1(n_23),
.B2(n_10),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_29),
.B1(n_14),
.B2(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_22),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_21),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_22),
.A2(n_15),
.B1(n_12),
.B2(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_27),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_14),
.B1(n_10),
.B2(n_4),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_45),
.C(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_29),
.B1(n_25),
.B2(n_28),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_44),
.Y(n_46)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_41),
.C(n_43),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

BUFx24_ASAP7_75t_SL g54 ( 
.A(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_50),
.Y(n_55)
);


endmodule