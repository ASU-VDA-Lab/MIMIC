module fake_jpeg_2421_n_440 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_440);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_440;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_46),
.B(n_48),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_47),
.B(n_71),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_56),
.B(n_63),
.Y(n_136)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_59),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_16),
.B(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_68),
.B(n_70),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_1),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_75),
.B(n_80),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_78),
.B(n_88),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_36),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_35),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_86),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_35),
.B1(n_24),
.B2(n_33),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_89),
.A2(n_98),
.B1(n_99),
.B2(n_102),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_37),
.B1(n_15),
.B2(n_25),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_93),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_33),
.B1(n_26),
.B2(n_37),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_37),
.B1(n_15),
.B2(n_25),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_33),
.B1(n_26),
.B2(n_15),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_54),
.A2(n_35),
.B1(n_33),
.B2(n_42),
.Y(n_109)
);

AO22x1_ASAP7_75t_L g175 ( 
.A1(n_109),
.A2(n_129),
.B1(n_138),
.B2(n_58),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_49),
.A2(n_41),
.B(n_29),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_122),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_66),
.Y(n_122)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_67),
.A2(n_42),
.B1(n_39),
.B2(n_26),
.Y(n_127)
);

BUFx24_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_74),
.A2(n_41),
.B1(n_29),
.B2(n_39),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_57),
.B(n_42),
.C(n_18),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_81),
.C(n_72),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_67),
.A2(n_18),
.B1(n_38),
.B2(n_34),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_66),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_140),
.Y(n_218)
);

OR2x4_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_85),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_141),
.A2(n_154),
.B(n_156),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_97),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_142),
.Y(n_209)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_132),
.B(n_88),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_147),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_59),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_150),
.Y(n_196)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_133),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_174),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_97),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_151),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_78),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_134),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_152),
.Y(n_217)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_153),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_87),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_112),
.B(n_83),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_155),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_91),
.B(n_84),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_103),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_157),
.Y(n_212)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_98),
.A3(n_102),
.B1(n_118),
.B2(n_129),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_158),
.A2(n_163),
.B(n_176),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_108),
.B(n_123),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_166),
.Y(n_203)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_38),
.B(n_31),
.C(n_34),
.Y(n_163)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_165),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_73),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_113),
.B(n_31),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_177),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_114),
.B(n_21),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_114),
.B(n_21),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_169),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_40),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_170),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_172),
.Y(n_219)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_92),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_175),
.A2(n_184),
.B1(n_115),
.B2(n_124),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_95),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_127),
.A2(n_40),
.B(n_32),
.C(n_30),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_100),
.B(n_61),
.Y(n_178)
);

AND2x4_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_126),
.Y(n_186)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_94),
.B(n_79),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_69),
.C(n_64),
.Y(n_213)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_94),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_100),
.Y(n_183)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_101),
.B(n_77),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_186),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_190),
.A2(n_192),
.B1(n_197),
.B2(n_218),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_139),
.A2(n_125),
.B1(n_101),
.B2(n_106),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_191),
.A2(n_194),
.B1(n_198),
.B2(n_205),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_93),
.B(n_99),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_192),
.A2(n_191),
.B(n_176),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_124),
.B1(n_121),
.B2(n_116),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_106),
.B1(n_116),
.B2(n_115),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_182),
.A2(n_121),
.B1(n_111),
.B2(n_105),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_204),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_145),
.A2(n_111),
.B1(n_105),
.B2(n_76),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_154),
.Y(n_211)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_178),
.Y(n_230)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_150),
.Y(n_214)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_146),
.Y(n_216)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_223),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_247),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_224),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_227),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_141),
.B(n_140),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_228),
.A2(n_234),
.B(n_236),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_167),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_243),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_230),
.B(n_251),
.Y(n_286)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_231),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_196),
.B(n_214),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_232),
.B(n_238),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_140),
.C(n_155),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_233),
.B(n_241),
.C(n_250),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_215),
.A2(n_171),
.B(n_174),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_202),
.A2(n_171),
.B(n_163),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_237),
.A2(n_257),
.B1(n_161),
.B2(n_181),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_188),
.B(n_193),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_155),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_158),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_186),
.B(n_157),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_245),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_209),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_189),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_249),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_157),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_156),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_156),
.C(n_178),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_203),
.B(n_183),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_207),
.Y(n_273)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_185),
.Y(n_254)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_186),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_255),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_210),
.A2(n_175),
.B(n_171),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_256),
.A2(n_259),
.B(n_187),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_212),
.A2(n_164),
.B1(n_180),
.B2(n_175),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_198),
.B(n_164),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_199),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_243),
.A2(n_205),
.B1(n_208),
.B2(n_185),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_264),
.A2(n_268),
.B1(n_282),
.B2(n_235),
.Y(n_304)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_225),
.Y(n_265)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

OAI22x1_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_186),
.B1(n_160),
.B2(n_165),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_269),
.B(n_275),
.Y(n_323)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_225),
.Y(n_270)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_245),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_251),
.Y(n_299)
);

NAND3xp33_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_248),
.C(n_232),
.Y(n_295)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_244),
.Y(n_275)
);

BUFx8_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_276),
.Y(n_307)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_259),
.A2(n_207),
.B1(n_219),
.B2(n_201),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_242),
.A2(n_213),
.B1(n_186),
.B2(n_219),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_292),
.B1(n_233),
.B2(n_245),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_284),
.A2(n_285),
.B(n_287),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_236),
.A2(n_206),
.B(n_187),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_228),
.A2(n_206),
.B(n_195),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_288),
.A2(n_289),
.B(n_278),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_256),
.A2(n_195),
.B(n_222),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_290),
.B(n_153),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_260),
.A2(n_220),
.B1(n_161),
.B2(n_216),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_252),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_217),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_295),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_240),
.Y(n_296)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_296),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_250),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_303),
.C(n_311),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_240),
.Y(n_298)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_298),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_299),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_229),
.Y(n_301)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_301),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_277),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_314),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_230),
.C(n_241),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_258),
.B1(n_257),
.B2(n_242),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_272),
.Y(n_308)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_308),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_284),
.A2(n_246),
.B1(n_247),
.B2(n_231),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_309),
.A2(n_269),
.B1(n_275),
.B2(n_274),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_310),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_220),
.C(n_200),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_239),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_268),
.A2(n_246),
.B1(n_162),
.B2(n_221),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_316),
.A2(n_263),
.B1(n_265),
.B2(n_270),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_267),
.A2(n_261),
.B(n_289),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_322),
.B(n_287),
.Y(n_324)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_319),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_320),
.B(n_32),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_291),
.A2(n_279),
.B1(n_273),
.B2(n_262),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

OAI32xp33_ASAP7_75t_L g322 ( 
.A1(n_278),
.A2(n_217),
.A3(n_200),
.B1(n_221),
.B2(n_162),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_324),
.A2(n_327),
.B(n_331),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_312),
.A2(n_267),
.B(n_288),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_319),
.Y(n_329)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_329),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_290),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_330),
.B(n_339),
.Y(n_365)
);

A2O1A1O1Ixp25_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_280),
.B(n_261),
.C(n_276),
.D(n_294),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_332),
.A2(n_335),
.B1(n_340),
.B2(n_349),
.Y(n_354)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_333),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_305),
.A2(n_263),
.B1(n_276),
.B2(n_281),
.Y(n_334)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_334),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_304),
.A2(n_276),
.B1(n_293),
.B2(n_179),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_293),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_310),
.A2(n_301),
.B1(n_298),
.B2(n_296),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_173),
.B(n_30),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_341),
.A2(n_316),
.B(n_322),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_345),
.B(n_303),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_297),
.B(n_62),
.C(n_60),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_325),
.C(n_311),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_309),
.A2(n_32),
.B1(n_30),
.B2(n_20),
.Y(n_349)
);

MAJx2_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_363),
.C(n_369),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_347),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_356),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_324),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_367),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_345),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_347),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_320),
.C(n_307),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_358),
.C(n_337),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_346),
.B(n_300),
.C(n_313),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_361),
.A2(n_333),
.B1(n_342),
.B2(n_331),
.Y(n_387)
);

FAx1_ASAP7_75t_SL g362 ( 
.A(n_327),
.B(n_323),
.CI(n_317),
.CON(n_362),
.SN(n_362)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_364),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_323),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_326),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_337),
.A2(n_317),
.B(n_315),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_343),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_315),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_336),
.B(n_313),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_370),
.B(n_338),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_368),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_376),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_375),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_334),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_358),
.C(n_366),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_364),
.A2(n_342),
.B1(n_348),
.B2(n_328),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_377),
.A2(n_354),
.B1(n_369),
.B2(n_360),
.Y(n_389)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_352),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_378),
.B(n_384),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_379),
.B(n_383),
.Y(n_398)
);

OAI21xp33_ASAP7_75t_L g381 ( 
.A1(n_366),
.A2(n_338),
.B(n_328),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_381),
.A2(n_361),
.B(n_360),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_382),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_367),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_365),
.B(n_348),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_386),
.B(n_300),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_359),
.Y(n_393)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_389),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_377),
.A2(n_363),
.B1(n_354),
.B2(n_353),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_390),
.B(n_391),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_374),
.C(n_376),
.Y(n_391)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_394),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_350),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_395),
.B(n_396),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_381),
.A2(n_359),
.B1(n_362),
.B2(n_341),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_397),
.A2(n_373),
.B1(n_382),
.B2(n_362),
.Y(n_405)
);

BUFx24_ASAP7_75t_SL g401 ( 
.A(n_372),
.Y(n_401)
);

OAI221xp5_ASAP7_75t_L g413 ( 
.A1(n_401),
.A2(n_32),
.B1(n_4),
.B2(n_6),
.C(n_7),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_385),
.C(n_380),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_404),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_399),
.A2(n_398),
.B(n_400),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_405),
.A2(n_408),
.B1(n_409),
.B2(n_32),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_397),
.A2(n_373),
.B1(n_384),
.B2(n_349),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_393),
.A2(n_335),
.B1(n_378),
.B2(n_319),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_410),
.B(n_395),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_391),
.A2(n_32),
.B(n_3),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_411),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_413),
.B(n_405),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_412),
.B(n_402),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_415),
.B(n_416),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_410),
.B(n_388),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_420),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_418),
.B(n_419),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_407),
.B(n_2),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_421),
.A2(n_423),
.B1(n_411),
.B2(n_409),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_6),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_422),
.B(n_7),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_408),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_423),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_426),
.B(n_428),
.Y(n_432)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_427),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_414),
.B(n_7),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_430),
.B(n_8),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_417),
.C(n_10),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_433),
.B(n_429),
.C(n_424),
.Y(n_435)
);

AO21x1_ASAP7_75t_L g436 ( 
.A1(n_434),
.A2(n_429),
.B(n_10),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_435),
.A2(n_436),
.B(n_431),
.Y(n_437)
);

AOI321xp33_ASAP7_75t_L g438 ( 
.A1(n_437),
.A2(n_8),
.A3(n_11),
.B1(n_12),
.B2(n_432),
.C(n_430),
.Y(n_438)
);

AOI21x1_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_12),
.B(n_8),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_11),
.C(n_12),
.Y(n_440)
);


endmodule