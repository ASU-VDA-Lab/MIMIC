module fake_netlist_1_12617_n_729 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_96, n_39, n_729);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_96;
input n_39;
output n_729;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_490;
wire n_247;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_699;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g98 ( .A(n_35), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_83), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_64), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_48), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_45), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_0), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_70), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_1), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_23), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_63), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_8), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_9), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_96), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_89), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_47), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_5), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_62), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_74), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_28), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_6), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_55), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_42), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_8), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_95), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_19), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_71), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_51), .Y(n_127) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_24), .Y(n_128) );
CKINVDCx16_ASAP7_75t_R g129 ( .A(n_17), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_2), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_56), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_33), .Y(n_132) );
INVxp33_ASAP7_75t_SL g133 ( .A(n_39), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_52), .Y(n_134) );
INVx4_ASAP7_75t_R g135 ( .A(n_91), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_49), .Y(n_136) );
AND2x2_ASAP7_75t_SL g137 ( .A(n_128), .B(n_97), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_129), .B(n_120), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_98), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_98), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_104), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_104), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_107), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_105), .B(n_1), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_107), .Y(n_145) );
AND2x6_ASAP7_75t_L g146 ( .A(n_110), .B(n_25), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_110), .Y(n_147) );
INVx1_ASAP7_75t_SL g148 ( .A(n_105), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_112), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_124), .B(n_2), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_112), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_121), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_121), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_123), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_123), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_126), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_144), .B(n_126), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_140), .B(n_131), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_152), .Y(n_161) );
BUFx10_ASAP7_75t_L g162 ( .A(n_144), .Y(n_162) );
AND2x6_ASAP7_75t_L g163 ( .A(n_144), .B(n_131), .Y(n_163) );
BUFx4f_ASAP7_75t_L g164 ( .A(n_146), .Y(n_164) );
INVxp67_ASAP7_75t_SL g165 ( .A(n_148), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_152), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_152), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_152), .Y(n_168) );
OR2x2_ASAP7_75t_L g169 ( .A(n_138), .B(n_129), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_140), .B(n_128), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_143), .B(n_103), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_155), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
INVx8_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_146), .A2(n_125), .B1(n_103), .B2(n_113), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_143), .B(n_108), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_155), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_145), .B(n_113), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_145), .B(n_132), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_151), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_146), .A2(n_130), .B1(n_125), .B2(n_115), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_146), .A2(n_130), .B1(n_115), .B2(n_119), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_184), .B(n_151), .Y(n_187) );
NOR2x1p5_ASAP7_75t_L g188 ( .A(n_165), .B(n_150), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_184), .B(n_153), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_170), .B(n_153), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_157), .B(n_137), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_170), .B(n_154), .Y(n_192) );
OR2x6_ASAP7_75t_SL g193 ( .A(n_169), .B(n_109), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_159), .A2(n_137), .B1(n_146), .B2(n_154), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_181), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_169), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_181), .A2(n_156), .B(n_149), .C(n_147), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_159), .A2(n_137), .B1(n_156), .B2(n_147), .Y(n_198) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_159), .Y(n_199) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_173), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_178), .B(n_141), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_180), .B(n_141), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_157), .B(n_133), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_157), .B(n_99), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_164), .A2(n_149), .B(n_142), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_157), .B(n_100), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_159), .A2(n_142), .B1(n_106), .B2(n_119), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_180), .B(n_101), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_183), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_183), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_180), .B(n_102), .Y(n_212) );
NAND2x1p5_ASAP7_75t_L g213 ( .A(n_164), .B(n_132), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_180), .B(n_111), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_173), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_171), .B(n_122), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_162), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_173), .Y(n_218) );
NOR2x1_ASAP7_75t_L g219 ( .A(n_160), .B(n_116), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_164), .B(n_114), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_159), .A2(n_117), .B1(n_116), .B2(n_134), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_159), .A2(n_117), .B1(n_127), .B2(n_118), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_164), .B(n_136), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_160), .A2(n_135), .B(n_4), .C(n_5), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_192), .B(n_159), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_198), .A2(n_163), .B1(n_162), .B2(n_185), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_198), .A2(n_163), .B1(n_162), .B2(n_186), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_203), .Y(n_228) );
OR2x2_ASAP7_75t_L g229 ( .A(n_216), .B(n_171), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_192), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_192), .B(n_163), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_195), .Y(n_232) );
NAND3xp33_ASAP7_75t_L g233 ( .A(n_194), .B(n_177), .C(n_182), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_217), .B(n_174), .Y(n_234) );
NOR2x1_ASAP7_75t_L g235 ( .A(n_188), .B(n_182), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_217), .B(n_174), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_208), .A2(n_174), .B1(n_163), .B2(n_162), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_192), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_190), .A2(n_174), .B(n_167), .C(n_175), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_195), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_188), .B(n_163), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_224), .A2(n_174), .B(n_167), .C(n_175), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_191), .A2(n_163), .B1(n_166), .B2(n_176), .Y(n_243) );
O2A1O1Ixp5_ASAP7_75t_L g244 ( .A1(n_197), .A2(n_179), .B(n_158), .C(n_172), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_216), .B(n_163), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_210), .Y(n_246) );
AO32x1_ASAP7_75t_L g247 ( .A1(n_210), .A2(n_172), .A3(n_168), .B1(n_161), .B2(n_158), .Y(n_247) );
OAI22x1_ASAP7_75t_L g248 ( .A1(n_208), .A2(n_163), .B1(n_4), .B2(n_6), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_187), .A2(n_179), .B(n_168), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_202), .A2(n_176), .B(n_166), .C(n_161), .Y(n_250) );
OR2x2_ASAP7_75t_SL g251 ( .A(n_193), .B(n_135), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_211), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_193), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_211), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_217), .B(n_166), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_189), .A2(n_176), .B(n_166), .C(n_9), .Y(n_256) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_244), .A2(n_206), .B(n_213), .Y(n_257) );
O2A1O1Ixp5_ASAP7_75t_L g258 ( .A1(n_242), .A2(n_204), .B(n_207), .C(n_205), .Y(n_258) );
INVx8_ASAP7_75t_L g259 ( .A(n_241), .Y(n_259) );
NOR2xp33_ASAP7_75t_SL g260 ( .A(n_253), .B(n_196), .Y(n_260) );
BUFx10_ASAP7_75t_L g261 ( .A(n_241), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_229), .B(n_209), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_230), .B(n_212), .Y(n_263) );
AOI221xp5_ASAP7_75t_SL g264 ( .A1(n_242), .A2(n_222), .B1(n_214), .B2(n_223), .C(n_220), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_232), .B(n_219), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_232), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_238), .B(n_217), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_235), .B(n_221), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g269 ( .A1(n_245), .A2(n_219), .B(n_213), .C(n_199), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_251), .B(n_221), .Y(n_270) );
AO31x2_ASAP7_75t_L g271 ( .A1(n_239), .A2(n_218), .A3(n_215), .B(n_201), .Y(n_271) );
AOI21xp33_ASAP7_75t_L g272 ( .A1(n_237), .A2(n_200), .B(n_213), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_239), .A2(n_218), .B(n_215), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_256), .A2(n_176), .B(n_215), .C(n_201), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_246), .Y(n_275) );
OAI22xp33_ASAP7_75t_L g276 ( .A1(n_226), .A2(n_201), .B1(n_218), .B2(n_10), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_248), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_L g278 ( .A1(n_228), .A2(n_3), .B(n_7), .C(n_10), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_266), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_259), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_270), .A2(n_227), .B(n_233), .C(n_250), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_266), .Y(n_282) );
OAI211xp5_ASAP7_75t_SL g283 ( .A1(n_278), .A2(n_244), .B(n_231), .C(n_225), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_262), .A2(n_246), .B1(n_254), .B2(n_252), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_263), .B(n_240), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_265), .B(n_255), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_273), .A2(n_247), .B(n_249), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_274), .A2(n_247), .B(n_255), .Y(n_288) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_257), .A2(n_236), .B(n_234), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_258), .A2(n_247), .B(n_236), .Y(n_290) );
OA21x2_ASAP7_75t_L g291 ( .A1(n_264), .A2(n_257), .B(n_277), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_265), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_260), .A2(n_234), .B1(n_243), .B2(n_11), .Y(n_293) );
AO31x2_ASAP7_75t_L g294 ( .A1(n_268), .A2(n_3), .A3(n_7), .B(n_11), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_263), .B(n_12), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_275), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_276), .A2(n_12), .B1(n_13), .B2(n_14), .C(n_15), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_275), .Y(n_299) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_269), .A2(n_54), .B(n_93), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_296), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_282), .Y(n_302) );
OAI21xp5_ASAP7_75t_L g303 ( .A1(n_281), .A2(n_264), .B(n_272), .Y(n_303) );
OA21x2_ASAP7_75t_L g304 ( .A1(n_288), .A2(n_271), .B(n_267), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_282), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_297), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_297), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_291), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_297), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_279), .Y(n_310) );
AO21x2_ASAP7_75t_L g311 ( .A1(n_290), .A2(n_271), .B(n_267), .Y(n_311) );
OA21x2_ASAP7_75t_L g312 ( .A1(n_287), .A2(n_271), .B(n_267), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_291), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_284), .A2(n_271), .B(n_275), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_291), .Y(n_315) );
INVx5_ASAP7_75t_L g316 ( .A(n_280), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_284), .A2(n_283), .B(n_295), .Y(n_317) );
OAI21xp5_ASAP7_75t_L g318 ( .A1(n_289), .A2(n_271), .B(n_275), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_292), .B(n_261), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_285), .B(n_261), .Y(n_320) );
AOI21xp5_ASAP7_75t_SL g321 ( .A1(n_298), .A2(n_280), .B(n_299), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_292), .B(n_259), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_291), .B(n_261), .Y(n_323) );
NOR2x1_ASAP7_75t_L g324 ( .A(n_296), .B(n_259), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_286), .B(n_13), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_299), .Y(n_326) );
OAI221xp5_ASAP7_75t_L g327 ( .A1(n_293), .A2(n_259), .B1(n_15), .B2(n_16), .C(n_17), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_289), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_294), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_286), .B(n_14), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_294), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_300), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_312), .B(n_294), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_302), .B(n_294), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_309), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_302), .B(n_294), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_302), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_308), .Y(n_338) );
INVx2_ASAP7_75t_SL g339 ( .A(n_310), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_310), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_320), .B(n_16), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_329), .B(n_300), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_312), .B(n_18), .Y(n_343) );
AO21x2_ASAP7_75t_L g344 ( .A1(n_303), .A2(n_18), .B(n_19), .Y(n_344) );
NOR2xp67_ASAP7_75t_L g345 ( .A(n_331), .B(n_59), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_328), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_305), .B(n_20), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_328), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_305), .B(n_20), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_310), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_312), .B(n_21), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_312), .B(n_21), .Y(n_352) );
OAI31xp33_ASAP7_75t_SL g353 ( .A1(n_327), .A2(n_22), .A3(n_23), .B(n_26), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_327), .A2(n_22), .B1(n_27), .B2(n_29), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_312), .B(n_94), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_328), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_312), .B(n_30), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_328), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_305), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_312), .B(n_311), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_310), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_311), .B(n_92), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_326), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_301), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_326), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_301), .Y(n_366) );
INVxp67_ASAP7_75t_L g367 ( .A(n_329), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_318), .B(n_31), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_326), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_329), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_314), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_301), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_308), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_311), .B(n_90), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_311), .B(n_32), .Y(n_375) );
INVx4_ASAP7_75t_L g376 ( .A(n_316), .Y(n_376) );
AO21x2_ASAP7_75t_L g377 ( .A1(n_303), .A2(n_34), .B(n_36), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_331), .B(n_88), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_331), .B(n_37), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_311), .B(n_87), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_301), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_331), .Y(n_382) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_318), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_314), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_323), .B(n_311), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_308), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_385), .B(n_323), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_363), .B(n_330), .Y(n_388) );
INVx5_ASAP7_75t_L g389 ( .A(n_376), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_361), .B(n_304), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_361), .Y(n_391) );
INVx5_ASAP7_75t_L g392 ( .A(n_376), .Y(n_392) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_376), .B(n_324), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_378), .A2(n_321), .B(n_332), .Y(n_394) );
NAND2x1p5_ASAP7_75t_L g395 ( .A(n_376), .B(n_316), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_363), .B(n_330), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_337), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_337), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_338), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_385), .B(n_304), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_365), .B(n_330), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_338), .Y(n_402) );
INVx4_ASAP7_75t_L g403 ( .A(n_376), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_359), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_385), .B(n_323), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_385), .B(n_304), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_359), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_385), .B(n_304), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_353), .B(n_317), .C(n_325), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_360), .B(n_304), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_360), .B(n_304), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_339), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_340), .B(n_304), .Y(n_413) );
BUFx12f_ASAP7_75t_L g414 ( .A(n_339), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_360), .B(n_323), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_343), .B(n_313), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_339), .B(n_325), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_343), .B(n_313), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_341), .A2(n_317), .B1(n_325), .B2(n_320), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_365), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_343), .B(n_315), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_340), .B(n_315), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_369), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_351), .B(n_315), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_369), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_372), .Y(n_426) );
NOR4xp25_ASAP7_75t_SL g427 ( .A(n_340), .B(n_332), .C(n_313), .D(n_316), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_351), .B(n_332), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_351), .B(n_309), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_372), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_352), .B(n_309), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_370), .B(n_335), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_352), .B(n_309), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_352), .B(n_307), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_350), .Y(n_435) );
AND2x4_ASAP7_75t_SL g436 ( .A(n_335), .B(n_307), .Y(n_436) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_364), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_338), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_381), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_333), .B(n_307), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_381), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_364), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_347), .B(n_324), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_370), .B(n_307), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_350), .Y(n_445) );
INVxp67_ASAP7_75t_L g446 ( .A(n_350), .Y(n_446) );
AND2x4_ASAP7_75t_SL g447 ( .A(n_335), .B(n_307), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_333), .B(n_307), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_333), .B(n_306), .Y(n_449) );
NAND4xp25_ASAP7_75t_L g450 ( .A(n_353), .B(n_324), .C(n_322), .D(n_319), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_366), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_366), .B(n_306), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_347), .Y(n_453) );
NOR2x1p5_ASAP7_75t_L g454 ( .A(n_362), .B(n_322), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_349), .B(n_319), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_349), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_341), .B(n_319), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_338), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_334), .B(n_316), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_386), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_373), .Y(n_461) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_378), .B(n_316), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_362), .B(n_306), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_362), .B(n_306), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_334), .B(n_316), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_336), .B(n_316), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_415), .B(n_335), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_415), .B(n_386), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_440), .B(n_335), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_389), .B(n_374), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_410), .B(n_411), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_417), .B(n_386), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_397), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_451), .B(n_386), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_399), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_440), .B(n_374), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_399), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_391), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_410), .B(n_336), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_411), .B(n_367), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_457), .B(n_316), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_402), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_403), .B(n_367), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_448), .B(n_374), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_453), .B(n_373), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_416), .B(n_373), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_398), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_456), .B(n_382), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_404), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_407), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_448), .B(n_380), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_402), .Y(n_492) );
NAND3xp33_ASAP7_75t_SL g493 ( .A(n_427), .B(n_354), .C(n_380), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_394), .A2(n_345), .B(n_379), .Y(n_494) );
NAND3x1_ASAP7_75t_L g495 ( .A(n_400), .B(n_380), .C(n_375), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_420), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_449), .B(n_375), .Y(n_497) );
OR2x6_ASAP7_75t_L g498 ( .A(n_403), .B(n_375), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_389), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_442), .B(n_382), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_403), .B(n_383), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_423), .B(n_383), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_425), .B(n_384), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_426), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_449), .B(n_387), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_416), .B(n_384), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_430), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_439), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_441), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_461), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_422), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_389), .B(n_384), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_387), .B(n_371), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_422), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_418), .B(n_371), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_387), .B(n_371), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_438), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_418), .B(n_357), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_405), .B(n_355), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_421), .B(n_357), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_421), .B(n_378), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_438), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_424), .B(n_357), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_405), .B(n_355), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_458), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_424), .B(n_355), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_458), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_460), .B(n_344), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_405), .B(n_368), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_460), .B(n_344), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_450), .B(n_316), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_389), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_388), .B(n_344), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_396), .B(n_344), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_437), .B(n_379), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_429), .B(n_368), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_459), .B(n_379), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_452), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_429), .B(n_368), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_412), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_431), .B(n_368), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_389), .B(n_368), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_401), .B(n_344), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_435), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_431), .B(n_306), .Y(n_545) );
NOR2xp33_ASAP7_75t_SL g546 ( .A(n_392), .B(n_345), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_465), .B(n_342), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_445), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_466), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_390), .B(n_342), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_400), .B(n_342), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_433), .B(n_306), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_406), .B(n_348), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_433), .B(n_348), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_446), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_392), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_390), .B(n_348), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_505), .B(n_406), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_478), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_467), .B(n_408), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_513), .B(n_408), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_485), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_471), .B(n_413), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_474), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_471), .B(n_409), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_485), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_479), .B(n_428), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_479), .B(n_428), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_516), .B(n_434), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_473), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_549), .B(n_414), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_511), .B(n_432), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_468), .B(n_413), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_557), .Y(n_574) );
NOR2xp33_ASAP7_75t_SL g575 ( .A(n_498), .B(n_392), .Y(n_575) );
NAND3xp33_ASAP7_75t_L g576 ( .A(n_544), .B(n_419), .C(n_392), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_487), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_514), .B(n_432), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_489), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_498), .A2(n_454), .B1(n_419), .B2(n_462), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_469), .B(n_434), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_553), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_490), .Y(n_583) );
CKINVDCx16_ASAP7_75t_R g584 ( .A(n_498), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_503), .B(n_432), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_496), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_504), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_499), .Y(n_588) );
INVxp67_ASAP7_75t_SL g589 ( .A(n_553), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_475), .Y(n_590) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_495), .A2(n_354), .B(n_395), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_503), .B(n_444), .Y(n_592) );
NAND2x1p5_ASAP7_75t_L g593 ( .A(n_499), .B(n_392), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_502), .B(n_444), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_551), .B(n_464), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_555), .B(n_414), .Y(n_596) );
NAND2x1p5_ASAP7_75t_L g597 ( .A(n_542), .B(n_393), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_519), .B(n_464), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_524), .B(n_463), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_538), .B(n_443), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_502), .B(n_444), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_551), .B(n_463), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_531), .A2(n_455), .B1(n_395), .B2(n_377), .Y(n_603) );
AND2x2_ASAP7_75t_SL g604 ( .A(n_542), .B(n_447), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_532), .B(n_556), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_507), .Y(n_606) );
NOR2xp33_ASAP7_75t_SL g607 ( .A(n_546), .B(n_462), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_508), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_509), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_529), .B(n_447), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_477), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_545), .B(n_436), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_540), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_548), .B(n_358), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_480), .B(n_358), .Y(n_615) );
NOR2x1p5_ASAP7_75t_L g616 ( .A(n_493), .B(n_322), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_481), .A2(n_377), .B1(n_436), .B2(n_316), .Y(n_617) );
NAND2x1_ASAP7_75t_L g618 ( .A(n_483), .B(n_358), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_488), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_480), .B(n_356), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_486), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_552), .B(n_356), .Y(n_622) );
NAND2xp33_ASAP7_75t_SL g623 ( .A(n_470), .B(n_483), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_488), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_501), .B(n_356), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_533), .B(n_346), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_554), .B(n_346), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_500), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_482), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_500), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_565), .B(n_515), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_562), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_628), .B(n_515), .Y(n_633) );
INVxp67_ASAP7_75t_L g634 ( .A(n_559), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_566), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_563), .B(n_550), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_613), .A2(n_533), .B1(n_543), .B2(n_534), .C(n_476), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_619), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_624), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_630), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_621), .Y(n_641) );
NOR2xp67_ASAP7_75t_L g642 ( .A(n_580), .B(n_494), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_582), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_589), .B(n_543), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_567), .B(n_534), .Y(n_645) );
A2O1A1Ixp33_ASAP7_75t_L g646 ( .A1(n_623), .A2(n_494), .B(n_501), .C(n_512), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_570), .B(n_506), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_577), .Y(n_648) );
INVx1_ASAP7_75t_SL g649 ( .A(n_605), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_579), .Y(n_650) );
INVx2_ASAP7_75t_SL g651 ( .A(n_604), .Y(n_651) );
AOI322xp5_ASAP7_75t_L g652 ( .A1(n_584), .A2(n_526), .A3(n_518), .B1(n_520), .B2(n_523), .C1(n_484), .C2(n_497), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_583), .B(n_547), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_567), .B(n_472), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_586), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_588), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_616), .A2(n_491), .B1(n_512), .B2(n_539), .Y(n_657) );
AOI211xp5_ASAP7_75t_SL g658 ( .A1(n_580), .A2(n_546), .B(n_523), .C(n_518), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_573), .B(n_521), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_568), .B(n_510), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_618), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_568), .B(n_526), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_587), .Y(n_663) );
OAI221xp5_ASAP7_75t_SL g664 ( .A1(n_603), .A2(n_520), .B1(n_536), .B2(n_541), .C(n_537), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_594), .B(n_522), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_594), .B(n_527), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_591), .A2(n_530), .B(n_528), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_561), .B(n_517), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_593), .A2(n_535), .B1(n_525), .B2(n_492), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_606), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_608), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_596), .B(n_530), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_564), .Y(n_673) );
OAI21xp33_ASAP7_75t_L g674 ( .A1(n_652), .A2(n_578), .B(n_572), .Y(n_674) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_646), .B(n_576), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_642), .A2(n_575), .B(n_591), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_632), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_664), .A2(n_609), .B1(n_600), .B2(n_585), .C(n_572), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_656), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_631), .B(n_601), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_635), .Y(n_681) );
OAI31xp33_ASAP7_75t_L g682 ( .A1(n_658), .A2(n_593), .A3(n_597), .B(n_571), .Y(n_682) );
AND2x2_ASAP7_75t_SL g683 ( .A(n_673), .B(n_607), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_637), .B(n_601), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_643), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_661), .B(n_597), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_636), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g688 ( .A1(n_651), .A2(n_617), .B1(n_585), .B2(n_592), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_667), .A2(n_592), .B(n_578), .C(n_625), .Y(n_689) );
OAI222xp33_ASAP7_75t_L g690 ( .A1(n_657), .A2(n_595), .B1(n_602), .B2(n_610), .C1(n_558), .C2(n_560), .Y(n_690) );
AOI322xp5_ASAP7_75t_L g691 ( .A1(n_641), .A2(n_599), .A3(n_598), .B1(n_569), .B2(n_581), .C1(n_574), .C2(n_620), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_649), .A2(n_625), .B(n_612), .C(n_615), .Y(n_692) );
AOI322xp5_ASAP7_75t_L g693 ( .A1(n_662), .A2(n_620), .A3(n_615), .B1(n_627), .B2(n_622), .C1(n_626), .C2(n_614), .Y(n_693) );
INVx1_ASAP7_75t_SL g694 ( .A(n_673), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_672), .A2(n_626), .B(n_614), .C(n_629), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g696 ( .A1(n_634), .A2(n_611), .B1(n_590), .B2(n_528), .C(n_346), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_686), .A2(n_670), .B(n_634), .Y(n_697) );
AOI222xp33_ASAP7_75t_L g698 ( .A1(n_678), .A2(n_670), .B1(n_644), .B2(n_647), .C1(n_669), .C2(n_639), .Y(n_698) );
AOI211xp5_ASAP7_75t_SL g699 ( .A1(n_676), .A2(n_647), .B(n_653), .C(n_633), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_679), .B(n_653), .Y(n_700) );
INVx1_ASAP7_75t_SL g701 ( .A(n_694), .Y(n_701) );
NOR2x1_ASAP7_75t_L g702 ( .A(n_686), .B(n_655), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_674), .A2(n_645), .B1(n_638), .B2(n_640), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_688), .A2(n_671), .B1(n_648), .B2(n_650), .C(n_663), .Y(n_704) );
AOI222xp33_ASAP7_75t_L g705 ( .A1(n_683), .A2(n_660), .B1(n_666), .B2(n_665), .C1(n_654), .C2(n_668), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_692), .A2(n_659), .B1(n_377), .B2(n_41), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_687), .Y(n_707) );
NAND2xp33_ASAP7_75t_SL g708 ( .A(n_682), .B(n_377), .Y(n_708) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_708), .A2(n_688), .B(n_690), .C(n_684), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_698), .A2(n_675), .B1(n_683), .B2(n_689), .Y(n_710) );
NAND4xp25_ASAP7_75t_L g711 ( .A(n_699), .B(n_691), .C(n_693), .D(n_695), .Y(n_711) );
NAND5xp2_ASAP7_75t_L g712 ( .A(n_705), .B(n_685), .C(n_696), .D(n_680), .E(n_681), .Y(n_712) );
AOI322xp5_ASAP7_75t_L g713 ( .A1(n_703), .A2(n_677), .A3(n_377), .B1(n_43), .B2(n_44), .C1(n_46), .C2(n_50), .Y(n_713) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_704), .A2(n_38), .B1(n_40), .B2(n_53), .C(n_57), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_709), .Y(n_715) );
NOR4xp75_ASAP7_75t_L g716 ( .A(n_714), .B(n_706), .C(n_701), .D(n_702), .Y(n_716) );
NOR5xp2_ASAP7_75t_L g717 ( .A(n_711), .B(n_707), .C(n_697), .D(n_700), .E(n_65), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_710), .B(n_58), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_715), .B(n_713), .Y(n_719) );
NOR4xp25_ASAP7_75t_L g720 ( .A(n_718), .B(n_712), .C(n_61), .D(n_66), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_717), .B(n_60), .Y(n_721) );
OAI21xp5_ASAP7_75t_L g722 ( .A1(n_719), .A2(n_716), .B(n_68), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_721), .A2(n_67), .B1(n_69), .B2(n_73), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_723), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_722), .Y(n_725) );
AOI222xp33_ASAP7_75t_SL g726 ( .A1(n_724), .A2(n_720), .B1(n_76), .B2(n_77), .C1(n_78), .C2(n_79), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g727 ( .A1(n_726), .A2(n_725), .B(n_81), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_727), .A2(n_75), .B(n_82), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_728), .A2(n_84), .B1(n_85), .B2(n_86), .Y(n_729) );
endmodule