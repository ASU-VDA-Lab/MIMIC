module fake_jpeg_1412_n_224 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_224);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_13),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_23),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_8),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_10),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_83),
.Y(n_88)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx5_ASAP7_75t_SL g97 ( 
.A(n_81),
.Y(n_97)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_63),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_93),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_74),
.B(n_60),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_74),
.B1(n_58),
.B2(n_72),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_92),
.B1(n_58),
.B2(n_52),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_94),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_55),
.B1(n_73),
.B2(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_76),
.B(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_65),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_55),
.B1(n_60),
.B2(n_52),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_56),
.B(n_97),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_87),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_54),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_51),
.B1(n_72),
.B2(n_75),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_81),
.B1(n_62),
.B2(n_75),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_61),
.B1(n_59),
.B2(n_56),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_53),
.B1(n_4),
.B2(n_5),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_61),
.B1(n_59),
.B2(n_57),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_3),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_0),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_116),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_0),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_97),
.B(n_62),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_104),
.B(n_110),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_131),
.Y(n_143)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_1),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_130),
.B(n_133),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_135),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_1),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_99),
.C(n_108),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_157),
.C(n_161),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_145),
.Y(n_178)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_110),
.A3(n_109),
.B1(n_98),
.B2(n_53),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_152),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_137),
.B(n_3),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_121),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_153),
.B(n_42),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_24),
.C(n_45),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_6),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_159),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_125),
.B1(n_12),
.B2(n_13),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_26),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_150),
.A2(n_134),
.B1(n_129),
.B2(n_122),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_167),
.B1(n_182),
.B2(n_15),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_138),
.B1(n_155),
.B2(n_143),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_141),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_170),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_122),
.B(n_125),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_171),
.A2(n_34),
.B(n_33),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_173),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_47),
.B(n_30),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_147),
.B(n_11),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_180),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_157),
.B(n_15),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_155),
.A2(n_41),
.B1(n_28),
.B2(n_31),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_139),
.C(n_161),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_190),
.C(n_191),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_174),
.B1(n_169),
.B2(n_168),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_25),
.C(n_38),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_39),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_16),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_194),
.B1(n_193),
.B2(n_188),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_182),
.B(n_175),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_183),
.B(n_17),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_168),
.C(n_181),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_178),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_199),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_183),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_204),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_171),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_192),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_205),
.B1(n_19),
.B2(n_20),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_206),
.Y(n_210)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_163),
.C(n_166),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_208),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_199),
.A2(n_164),
.B1(n_162),
.B2(n_32),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_201),
.B(n_198),
.Y(n_215)
);

AOI31xp67_ASAP7_75t_SL g218 ( 
.A1(n_215),
.A2(n_210),
.A3(n_207),
.B(n_208),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_218),
.B(n_216),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_217),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_220),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_214),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_19),
.B(n_20),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_223),
.Y(n_224)
);


endmodule