module fake_jpeg_5382_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_23),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_0),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_28),
.B1(n_18),
.B2(n_17),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_19),
.B1(n_22),
.B2(n_18),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_48),
.B(n_56),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_24),
.B1(n_23),
.B2(n_28),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_26),
.B1(n_36),
.B2(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_54),
.Y(n_75)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_55),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_27),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_17),
.B1(n_22),
.B2(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_60),
.Y(n_92)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_64),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_56),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_34),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_20),
.B1(n_50),
.B2(n_41),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_74),
.B(n_76),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_40),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_81),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_79),
.B(n_44),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_40),
.Y(n_94)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_43),
.A2(n_39),
.B(n_30),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_84),
.B(n_29),
.Y(n_109)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_41),
.B1(n_21),
.B2(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_93),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_98),
.B1(n_75),
.B2(n_74),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_40),
.B(n_55),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_89),
.A2(n_106),
.B(n_63),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_61),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_55),
.B1(n_53),
.B2(n_35),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_38),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_38),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_38),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_53),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_109),
.B1(n_82),
.B2(n_65),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_107),
.B(n_98),
.C(n_85),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_129),
.B(n_133),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_119),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_78),
.B1(n_76),
.B2(n_65),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_124),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_79),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_SL g135 ( 
.A1(n_121),
.A2(n_88),
.A3(n_105),
.B1(n_95),
.B2(n_87),
.C1(n_97),
.C2(n_104),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_73),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_108),
.B(n_29),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_81),
.B1(n_58),
.B2(n_57),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_29),
.B1(n_16),
.B2(n_31),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_90),
.Y(n_124)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_128),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_131),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_100),
.B1(n_87),
.B2(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_125),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_100),
.B(n_102),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_101),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_114),
.B(n_133),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_104),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_144),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_68),
.B1(n_83),
.B2(n_86),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_38),
.A3(n_92),
.B1(n_21),
.B2(n_31),
.C1(n_25),
.C2(n_16),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_92),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_130),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_116),
.B(n_124),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_60),
.B1(n_2),
.B2(n_3),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_38),
.C(n_60),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_123),
.C(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_112),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_96),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_161),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_117),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_141),
.C(n_153),
.Y(n_176)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_165),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_126),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_171),
.B(n_172),
.Y(n_184)
);

A2O1A1O1Ixp25_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_111),
.B(n_122),
.C(n_120),
.D(n_31),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_170),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_119),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_169),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_31),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_14),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_174),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_175),
.A2(n_140),
.B1(n_136),
.B2(n_156),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_178),
.C(n_187),
.Y(n_195)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_142),
.C(n_143),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_143),
.B1(n_150),
.B2(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_157),
.B1(n_172),
.B2(n_160),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_150),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_159),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_138),
.C(n_147),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_134),
.C(n_152),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_146),
.C(n_175),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_183),
.B(n_137),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_192),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_198),
.C(n_199),
.Y(n_203)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_200),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_R g196 ( 
.A(n_184),
.B(n_134),
.C(n_170),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_197),
.B(n_60),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_167),
.C(n_173),
.Y(n_199)
);

OA21x2_ASAP7_75t_SL g200 ( 
.A1(n_188),
.A2(n_173),
.B(n_13),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_196),
.B(n_189),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_208),
.C(n_209),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_178),
.B1(n_163),
.B2(n_179),
.Y(n_204)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_186),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_206),
.Y(n_211)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_195),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_216),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_207),
.A2(n_195),
.B(n_199),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_203),
.B(n_208),
.Y(n_218)
);

NOR2x1p5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_13),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_202),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_218),
.B(n_219),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_205),
.B(n_5),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_4),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_4),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_212),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_6),
.B(n_8),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_214),
.B(n_5),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_225),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_10),
.C2(n_11),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_227),
.B(n_223),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_10),
.Y(n_229)
);


endmodule