module fake_jpeg_23137_n_230 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_45),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

HAxp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_42),
.CON(n_47),
.SN(n_47)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_41),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_1),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_27),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_29),
.B1(n_19),
.B2(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_29),
.B1(n_19),
.B2(n_46),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_29),
.B1(n_19),
.B2(n_18),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_57),
.B1(n_58),
.B2(n_64),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_20),
.B1(n_32),
.B2(n_28),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_35),
.B1(n_20),
.B2(n_32),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_25),
.B1(n_22),
.B2(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_33),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_36),
.A2(n_35),
.B1(n_22),
.B2(n_28),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_75),
.B1(n_84),
.B2(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_17),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_77),
.Y(n_107)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_86),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_88),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_33),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_24),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_66),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_62),
.B1(n_53),
.B2(n_38),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_23),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_33),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_63),
.B1(n_42),
.B2(n_55),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_99),
.A2(n_87),
.B1(n_81),
.B2(n_85),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_47),
.B1(n_60),
.B2(n_43),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_103),
.B1(n_108),
.B2(n_116),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_60),
.B1(n_21),
.B2(n_23),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_78),
.A2(n_43),
.B(n_25),
.C(n_42),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_119),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_94),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_71),
.A2(n_38),
.B1(n_27),
.B2(n_62),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_38),
.C(n_53),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_1),
.C(n_3),
.Y(n_142)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_125),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_73),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_70),
.B(n_91),
.Y(n_126)
);

AOI221xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_144),
.B1(n_123),
.B2(n_145),
.C(n_125),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_128),
.B(n_136),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_82),
.B(n_70),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_131),
.B(n_143),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_112),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_137),
.Y(n_148)
);

AO22x1_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_88),
.B1(n_82),
.B2(n_76),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_90),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_140),
.B1(n_142),
.B2(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_81),
.B1(n_94),
.B2(n_4),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_121),
.B1(n_111),
.B2(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_117),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_4),
.B(n_5),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_145),
.B(n_7),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_6),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_7),
.B(n_8),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_149),
.B(n_156),
.Y(n_170)
);

NAND2x1_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_104),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_157),
.B(n_158),
.Y(n_182)
);

AOI22x1_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_113),
.B1(n_8),
.B2(n_7),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_159),
.B1(n_132),
.B2(n_124),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_110),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_162),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_165),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_129),
.C(n_127),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_152),
.C(n_147),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_174),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_175),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_127),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_150),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_167),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_181),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_159),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_154),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_182),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_177),
.C(n_180),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_147),
.B(n_154),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_194),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_162),
.C(n_158),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_196),
.C(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_153),
.B(n_165),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_143),
.C(n_153),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_184),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_197),
.B(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_204),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_176),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_207),
.B1(n_189),
.B2(n_190),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_187),
.B(n_163),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_201),
.B(n_205),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_202),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_192),
.A2(n_169),
.B1(n_181),
.B2(n_174),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_213),
.B1(n_204),
.B2(n_201),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_212),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_193),
.Y(n_212)
);

INVx13_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_169),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_188),
.B(n_196),
.Y(n_218)
);

OAI211xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_220),
.B(n_146),
.C(n_10),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_212),
.A2(n_214),
.B1(n_213),
.B2(n_211),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_218),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_SL g220 ( 
.A1(n_209),
.A2(n_151),
.B(n_170),
.C(n_163),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_215),
.C(n_210),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_106),
.C(n_220),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_224),
.B(n_9),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_220),
.A2(n_106),
.B(n_117),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_226),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_11),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_13),
.B(n_146),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_228),
.Y(n_230)
);


endmodule