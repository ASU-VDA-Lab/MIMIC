module fake_aes_7811_n_1159 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1159);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1159;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_627;
wire n_532;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_857;
wire n_786;
wire n_360;
wire n_345;
wire n_1090;
wire n_236;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1011;
wire n_1132;
wire n_1025;
wire n_880;
wire n_1101;
wire n_1155;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_230;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_1000;
wire n_893;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_1106;
wire n_982;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_1157;
wire n_876;
wire n_986;
wire n_886;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_622;
wire n_549;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_955;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_721;
wire n_438;
wire n_656;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_233;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_1042;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_924;
wire n_1043;
wire n_947;
wire n_378;
wire n_582;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_994;
wire n_930;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_919;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_1127;
wire n_269;
INVx1_ASAP7_75t_L g230 ( .A(n_98), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_194), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_190), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_170), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_120), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_111), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_166), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_89), .Y(n_237) );
BUFx10_ASAP7_75t_L g238 ( .A(n_95), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_167), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_113), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_182), .Y(n_241) );
INVxp33_ASAP7_75t_L g242 ( .A(n_156), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_32), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_9), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_109), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_102), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_84), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_22), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_75), .Y(n_249) );
INVxp67_ASAP7_75t_L g250 ( .A(n_64), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_78), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_96), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_164), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_142), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_150), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_198), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_146), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_68), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_97), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_225), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_140), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_126), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_79), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_160), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_229), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_155), .Y(n_266) );
NOR2xp67_ASAP7_75t_L g267 ( .A(n_60), .B(n_186), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_14), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_105), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_47), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_20), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_3), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_47), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_220), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_27), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_16), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_42), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_28), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_87), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_208), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_85), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_115), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_37), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_49), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_175), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_215), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_86), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_218), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_61), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_161), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_60), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_9), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_214), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_149), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_90), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_116), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_151), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_8), .Y(n_298) );
BUFx10_ASAP7_75t_L g299 ( .A(n_178), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_196), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_212), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_101), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_169), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_135), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_81), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_82), .Y(n_306) );
BUFx10_ASAP7_75t_L g307 ( .A(n_171), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_53), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_5), .Y(n_309) );
CKINVDCx16_ASAP7_75t_R g310 ( .A(n_127), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_204), .B(n_172), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_124), .Y(n_312) );
CKINVDCx16_ASAP7_75t_R g313 ( .A(n_88), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_21), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_104), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_211), .Y(n_316) );
INVxp33_ASAP7_75t_L g317 ( .A(n_0), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_40), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_217), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_173), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_157), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_144), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_195), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_80), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_193), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_153), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_54), .B(n_184), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_83), .Y(n_328) );
INVxp33_ASAP7_75t_L g329 ( .A(n_93), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_25), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_221), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_210), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_10), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_8), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_16), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_11), .Y(n_336) );
INVxp33_ASAP7_75t_L g337 ( .A(n_134), .Y(n_337) );
INVx1_ASAP7_75t_SL g338 ( .A(n_76), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_136), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_203), .Y(n_340) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_137), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_159), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_187), .Y(n_343) );
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_108), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_197), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_91), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_62), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_119), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_11), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_199), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_168), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_94), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_206), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_139), .Y(n_354) );
OAI21x1_ASAP7_75t_L g355 ( .A1(n_237), .A2(n_74), .B(n_73), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_341), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_268), .Y(n_357) );
INVx5_ASAP7_75t_L g358 ( .A(n_341), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_317), .B(n_0), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_268), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_270), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_244), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_317), .B(n_1), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_270), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_341), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_341), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_232), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_246), .B(n_1), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_237), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_294), .B(n_2), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_323), .B(n_2), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_284), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_247), .Y(n_373) );
OA21x2_ASAP7_75t_L g374 ( .A1(n_264), .A2(n_3), .B(n_4), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_264), .Y(n_375) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_327), .B(n_77), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_283), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_247), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_242), .B(n_6), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_298), .Y(n_380) );
INVx5_ASAP7_75t_L g381 ( .A(n_323), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_336), .B(n_7), .Y(n_382) );
OA21x2_ASAP7_75t_L g383 ( .A1(n_285), .A2(n_7), .B(n_10), .Y(n_383) );
BUFx3_ASAP7_75t_L g384 ( .A(n_234), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_243), .B(n_12), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_285), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_298), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_242), .B(n_12), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_284), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_372), .B(n_329), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_359), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_369), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_358), .Y(n_393) );
BUFx10_ASAP7_75t_L g394 ( .A(n_371), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_369), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_369), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_379), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_371), .B(n_330), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_372), .B(n_329), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_358), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_358), .Y(n_401) );
BUFx10_ASAP7_75t_L g402 ( .A(n_371), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_371), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_389), .B(n_337), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_358), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_389), .B(n_337), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_371), .B(n_310), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_379), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_367), .B(n_313), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_375), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_358), .Y(n_411) );
INVx2_ASAP7_75t_SL g412 ( .A(n_381), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_386), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_379), .B(n_344), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_359), .A2(n_273), .B1(n_275), .B2(n_271), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_384), .B(n_315), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_358), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_363), .A2(n_292), .B1(n_308), .B2(n_277), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_388), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_386), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_358), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_381), .B(n_230), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_374), .Y(n_425) );
BUFx10_ASAP7_75t_L g426 ( .A(n_376), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_358), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_384), .B(n_315), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_356), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_388), .B(n_238), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_356), .Y(n_431) );
INVx4_ASAP7_75t_SL g432 ( .A(n_384), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_384), .B(n_352), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_356), .Y(n_434) );
INVx5_ASAP7_75t_L g435 ( .A(n_381), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_381), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_388), .B(n_352), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_394), .B(n_376), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_425), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_430), .B(n_368), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_399), .B(n_363), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_425), .Y(n_442) );
OAI22xp5_ASAP7_75t_SL g443 ( .A1(n_408), .A2(n_373), .B1(n_362), .B2(n_378), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_397), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_390), .B(n_363), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_403), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_403), .Y(n_447) );
O2A1O1Ixp5_ASAP7_75t_L g448 ( .A1(n_407), .A2(n_368), .B(n_370), .C(n_382), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_399), .B(n_370), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_397), .A2(n_408), .B1(n_421), .B2(n_426), .Y(n_450) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_437), .A2(n_355), .B(n_376), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_394), .B(n_376), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_426), .A2(n_383), .B1(n_374), .B2(n_385), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_426), .A2(n_378), .B1(n_342), .B2(n_346), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_391), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_404), .B(n_381), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_406), .B(n_381), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_390), .B(n_231), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_416), .B(n_385), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_398), .Y(n_460) );
NOR2xp67_ASAP7_75t_L g461 ( .A(n_409), .B(n_357), .Y(n_461) );
INVx3_ASAP7_75t_L g462 ( .A(n_398), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_398), .B(n_231), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_394), .B(n_233), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_398), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_426), .A2(n_383), .B1(n_374), .B2(n_360), .Y(n_466) );
OR2x6_ASAP7_75t_L g467 ( .A(n_413), .B(n_355), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_402), .B(n_241), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_392), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_417), .B(n_304), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_420), .B(n_373), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_413), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_395), .Y(n_473) );
BUFx12f_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_429), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_418), .A2(n_342), .B1(n_346), .B2(n_304), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_418), .A2(n_272), .B1(n_276), .B2(n_248), .Y(n_477) );
NAND2xp33_ASAP7_75t_L g478 ( .A(n_412), .B(n_251), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_413), .B(n_272), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_424), .B(n_235), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_395), .A2(n_383), .B1(n_374), .B2(n_360), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_432), .B(n_387), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_396), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_429), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_429), .Y(n_485) );
BUFx4f_ASAP7_75t_SL g486 ( .A(n_410), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_410), .B(n_269), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_428), .B(n_357), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_414), .B(n_269), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_414), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_428), .B(n_361), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_431), .Y(n_492) );
AND3x1_ASAP7_75t_L g493 ( .A(n_415), .B(n_362), .C(n_333), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_415), .B(n_291), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_431), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_433), .B(n_361), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_422), .B(n_328), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_412), .A2(n_318), .B1(n_250), .B2(n_289), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_431), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_432), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_432), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_412), .A2(n_355), .B(n_239), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_432), .B(n_328), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_432), .B(n_340), .Y(n_504) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_434), .B(n_364), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_436), .B(n_236), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_434), .A2(n_374), .B1(n_383), .B2(n_377), .Y(n_507) );
INVx2_ASAP7_75t_SL g508 ( .A(n_393), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_393), .B(n_278), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_436), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_400), .A2(n_245), .B(n_240), .Y(n_511) );
BUFx3_ASAP7_75t_L g512 ( .A(n_435), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_435), .B(n_340), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_435), .B(n_249), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_400), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_435), .B(n_345), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_401), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_401), .A2(n_253), .B(n_252), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_435), .B(n_345), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_401), .B(n_380), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_405), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_474), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_444), .B(n_335), .Y(n_523) );
OR2x6_ASAP7_75t_L g524 ( .A(n_470), .B(n_330), .Y(n_524) );
INVx4_ASAP7_75t_L g525 ( .A(n_486), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_449), .B(n_445), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_439), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_441), .A2(n_334), .B(n_347), .C(n_309), .Y(n_528) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_482), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_464), .A2(n_419), .B(n_411), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_438), .A2(n_350), .B1(n_351), .B2(n_348), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_490), .B(n_350), .Y(n_532) );
INVx3_ASAP7_75t_L g533 ( .A(n_482), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_438), .A2(n_354), .B1(n_383), .B2(n_349), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_451), .A2(n_267), .B(n_387), .C(n_254), .Y(n_535) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_439), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_452), .A2(n_354), .B1(n_383), .B2(n_314), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_442), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_470), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_459), .B(n_238), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_464), .A2(n_423), .B(n_419), .Y(n_541) );
AND2x2_ASAP7_75t_SL g542 ( .A(n_476), .B(n_258), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_461), .B(n_255), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_479), .B(n_256), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_452), .A2(n_259), .B1(n_260), .B2(n_257), .Y(n_545) );
BUFx2_ASAP7_75t_L g546 ( .A(n_493), .Y(n_546) );
AOI33xp33_ASAP7_75t_L g547 ( .A1(n_455), .A2(n_305), .A3(n_262), .B1(n_263), .B2(n_265), .B3(n_353), .Y(n_547) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_512), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_458), .B(n_299), .Y(n_549) );
AOI21x1_ASAP7_75t_L g550 ( .A1(n_467), .A2(n_427), .B(n_311), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_454), .B(n_299), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_494), .B(n_299), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_460), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_456), .A2(n_311), .B(n_274), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_457), .A2(n_280), .B(n_266), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_450), .A2(n_258), .B1(n_286), .B2(n_281), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_465), .A2(n_288), .B(n_290), .C(n_287), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_460), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_448), .A2(n_293), .B(n_297), .C(n_295), .Y(n_559) );
O2A1O1Ixp5_ASAP7_75t_L g560 ( .A1(n_502), .A2(n_300), .B(n_302), .C(n_301), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_462), .B(n_303), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_462), .A2(n_440), .B1(n_443), .B2(n_446), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_477), .B(n_307), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_471), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_510), .A2(n_320), .B(n_319), .Y(n_565) );
OR2x6_ASAP7_75t_L g566 ( .A(n_483), .B(n_258), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_509), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_440), .B(n_307), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_453), .A2(n_322), .B(n_321), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_453), .A2(n_325), .B(n_324), .Y(n_570) );
INVx3_ASAP7_75t_L g571 ( .A(n_446), .Y(n_571) );
A2O1A1Ixp33_ASAP7_75t_L g572 ( .A1(n_488), .A2(n_326), .B(n_332), .C(n_331), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_469), .Y(n_573) );
NOR2xp33_ASAP7_75t_SL g574 ( .A(n_498), .B(n_261), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_463), .B(n_279), .Y(n_575) );
AO21x1_ASAP7_75t_L g576 ( .A1(n_480), .A2(n_343), .B(n_339), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_468), .A2(n_312), .B1(n_296), .B2(n_282), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_447), .A2(n_258), .B1(n_234), .B2(n_338), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_447), .B(n_13), .Y(n_579) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_507), .A2(n_365), .B(n_356), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_488), .B(n_306), .Y(n_581) );
BUFx4f_ASAP7_75t_L g582 ( .A(n_473), .Y(n_582) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_512), .Y(n_583) );
O2A1O1Ixp5_ASAP7_75t_L g584 ( .A1(n_480), .A2(n_366), .B(n_365), .C(n_316), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_506), .A2(n_365), .B(n_366), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_506), .A2(n_365), .B(n_366), .Y(n_586) );
O2A1O1Ixp33_ASAP7_75t_SL g587 ( .A1(n_514), .A2(n_123), .B(n_228), .C(n_227), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_487), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_491), .B(n_13), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_491), .B(n_14), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_489), .B(n_15), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_SL g592 ( .A1(n_514), .A2(n_121), .B(n_224), .C(n_223), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_496), .B(n_15), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_497), .B(n_17), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_496), .B(n_17), .Y(n_595) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_508), .Y(n_596) );
NAND2x1p5_ASAP7_75t_L g597 ( .A(n_472), .B(n_18), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_478), .A2(n_19), .B1(n_20), .B2(n_21), .Y(n_598) );
NOR2xp67_ASAP7_75t_SL g599 ( .A(n_503), .B(n_19), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_520), .Y(n_600) );
INVx3_ASAP7_75t_L g601 ( .A(n_500), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_520), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_513), .B(n_22), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_511), .B(n_23), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_504), .B(n_24), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_518), .B(n_24), .Y(n_606) );
OR2x6_ASAP7_75t_L g607 ( .A(n_501), .B(n_26), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_505), .B(n_28), .Y(n_608) );
BUFx2_ASAP7_75t_L g609 ( .A(n_516), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_481), .A2(n_29), .B1(n_30), .B2(n_31), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_519), .B(n_30), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_515), .B(n_31), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_481), .A2(n_32), .B1(n_33), .B2(n_34), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_517), .B(n_33), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_515), .B(n_34), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_521), .B(n_35), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_SL g617 ( .A1(n_475), .A2(n_141), .B(n_222), .C(n_219), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_499), .B(n_35), .Y(n_618) );
CKINVDCx10_ASAP7_75t_R g619 ( .A(n_484), .Y(n_619) );
INVx3_ASAP7_75t_L g620 ( .A(n_485), .Y(n_620) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_485), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_492), .B(n_36), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_495), .B(n_36), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_449), .B(n_37), .Y(n_624) );
BUFx12f_ASAP7_75t_L g625 ( .A(n_470), .Y(n_625) );
INVx11_ASAP7_75t_L g626 ( .A(n_474), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_449), .B(n_38), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_449), .B(n_38), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_502), .A2(n_143), .B(n_216), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_449), .A2(n_39), .B(n_40), .C(n_41), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_470), .B(n_39), .Y(n_631) );
O2A1O1Ixp33_ASAP7_75t_SL g632 ( .A1(n_451), .A2(n_145), .B(n_213), .C(n_209), .Y(n_632) );
NOR2xp67_ASAP7_75t_L g633 ( .A(n_454), .B(n_43), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_449), .B(n_44), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_439), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_438), .A2(n_44), .B1(n_45), .B2(n_46), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_438), .A2(n_45), .B1(n_46), .B2(n_48), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_438), .A2(n_48), .B1(n_49), .B2(n_50), .Y(n_638) );
INVx3_ASAP7_75t_L g639 ( .A(n_474), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_449), .B(n_51), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_486), .B(n_51), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_438), .A2(n_52), .B1(n_53), .B2(n_54), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_444), .B(n_55), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_526), .B(n_55), .Y(n_644) );
XNOR2xp5_ASAP7_75t_L g645 ( .A(n_524), .B(n_56), .Y(n_645) );
OAI22x1_ASAP7_75t_L g646 ( .A1(n_539), .A2(n_56), .B1(n_57), .B2(n_58), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_524), .B(n_57), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_624), .Y(n_648) );
O2A1O1Ixp33_ASAP7_75t_SL g649 ( .A1(n_535), .A2(n_148), .B(n_207), .C(n_205), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_627), .Y(n_650) );
INVxp67_ASAP7_75t_SL g651 ( .A(n_536), .Y(n_651) );
AO31x2_ASAP7_75t_L g652 ( .A1(n_569), .A2(n_59), .A3(n_61), .B(n_62), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_527), .A2(n_152), .B(n_202), .Y(n_653) );
NOR2xp67_ASAP7_75t_L g654 ( .A(n_525), .B(n_92), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_538), .A2(n_147), .B(n_201), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_567), .B(n_59), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_523), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_573), .B(n_63), .Y(n_658) );
BUFx10_ASAP7_75t_L g659 ( .A(n_524), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_625), .B(n_65), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_566), .A2(n_542), .B1(n_582), .B2(n_579), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_561), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_566), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_561), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_635), .A2(n_154), .B(n_200), .Y(n_665) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_548), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_564), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_643), .Y(n_668) );
AO31x2_ASAP7_75t_L g669 ( .A1(n_570), .A2(n_69), .A3(n_70), .B(n_71), .Y(n_669) );
INVx3_ASAP7_75t_SL g670 ( .A(n_525), .Y(n_670) );
INVx2_ASAP7_75t_SL g671 ( .A(n_619), .Y(n_671) );
AO31x2_ASAP7_75t_L g672 ( .A1(n_534), .A2(n_69), .A3(n_70), .B(n_71), .Y(n_672) );
A2O1A1Ixp33_ASAP7_75t_L g673 ( .A1(n_628), .A2(n_72), .B(n_99), .C(n_100), .Y(n_673) );
INVx1_ASAP7_75t_SL g674 ( .A(n_566), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_612), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_588), .B(n_72), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_633), .A2(n_103), .B1(n_106), .B2(n_107), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_551), .B(n_110), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g679 ( .A1(n_634), .A2(n_112), .B(n_114), .C(n_117), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_640), .A2(n_118), .B(n_122), .C(n_125), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_620), .Y(n_681) );
NOR2xp67_ASAP7_75t_L g682 ( .A(n_637), .B(n_128), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_582), .A2(n_129), .B1(n_130), .B2(n_131), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_546), .B(n_132), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_547), .B(n_133), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_528), .B(n_138), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_SL g687 ( .A1(n_559), .A2(n_158), .B(n_162), .C(n_163), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_563), .B(n_165), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_616), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_631), .Y(n_690) );
BUFx2_ASAP7_75t_L g691 ( .A(n_607), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_579), .A2(n_174), .B1(n_176), .B2(n_177), .Y(n_692) );
OA21x2_ASAP7_75t_L g693 ( .A1(n_560), .A2(n_179), .B(n_180), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_620), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_530), .A2(n_181), .B(n_183), .Y(n_695) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_548), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_604), .A2(n_185), .B1(n_188), .B2(n_189), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_571), .Y(n_698) );
OR2x2_ASAP7_75t_L g699 ( .A(n_552), .B(n_226), .Y(n_699) );
AND2x6_ASAP7_75t_L g700 ( .A(n_529), .B(n_191), .Y(n_700) );
NOR4xp25_ASAP7_75t_L g701 ( .A(n_630), .B(n_192), .C(n_613), .D(n_610), .Y(n_701) );
BUFx3_ASAP7_75t_L g702 ( .A(n_522), .Y(n_702) );
O2A1O1Ixp33_ASAP7_75t_L g703 ( .A1(n_572), .A2(n_557), .B(n_589), .C(n_593), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_574), .B(n_596), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_600), .B(n_602), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_541), .A2(n_537), .B(n_555), .Y(n_706) );
OA21x2_ASAP7_75t_L g707 ( .A1(n_554), .A2(n_622), .B(n_615), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_568), .A2(n_540), .B(n_581), .Y(n_708) );
OAI21x1_ASAP7_75t_L g709 ( .A1(n_601), .A2(n_584), .B(n_571), .Y(n_709) );
BUFx8_ASAP7_75t_L g710 ( .A(n_619), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_544), .A2(n_575), .B(n_549), .Y(n_711) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_548), .Y(n_712) );
INVx3_ASAP7_75t_L g713 ( .A(n_529), .Y(n_713) );
OAI22x1_ASAP7_75t_L g714 ( .A1(n_637), .A2(n_642), .B1(n_597), .B2(n_641), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_522), .B(n_639), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_590), .Y(n_716) );
NAND3x1_ASAP7_75t_L g717 ( .A(n_642), .B(n_598), .C(n_639), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_607), .B(n_532), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_591), .B(n_594), .C(n_605), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_558), .Y(n_720) );
OAI21xp5_ASAP7_75t_L g721 ( .A1(n_545), .A2(n_565), .B(n_595), .Y(n_721) );
OAI21xp5_ASAP7_75t_L g722 ( .A1(n_606), .A2(n_618), .B(n_603), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_607), .A2(n_638), .B1(n_636), .B2(n_556), .Y(n_723) );
OAI21x1_ASAP7_75t_L g724 ( .A1(n_585), .A2(n_586), .B(n_623), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g725 ( .A1(n_611), .A2(n_553), .B(n_608), .Y(n_725) );
AO21x2_ASAP7_75t_L g726 ( .A1(n_632), .A2(n_576), .B(n_617), .Y(n_726) );
NOR2xp67_ASAP7_75t_L g727 ( .A(n_533), .B(n_583), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_543), .A2(n_621), .B(n_609), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_614), .A2(n_599), .B(n_578), .C(n_531), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_577), .A2(n_533), .B(n_592), .Y(n_730) );
NAND3xp33_ASAP7_75t_SL g731 ( .A(n_626), .B(n_587), .C(n_529), .Y(n_731) );
OAI21xp5_ASAP7_75t_L g732 ( .A1(n_621), .A2(n_583), .B(n_596), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_596), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_526), .B(n_397), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_524), .A2(n_486), .B1(n_490), .B2(n_438), .Y(n_735) );
NOR2x1_ASAP7_75t_SL g736 ( .A(n_566), .B(n_607), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_536), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_526), .B(n_397), .Y(n_738) );
AO31x2_ASAP7_75t_L g739 ( .A1(n_535), .A2(n_570), .A3(n_569), .B(n_534), .Y(n_739) );
INVx4_ASAP7_75t_SL g740 ( .A(n_524), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_526), .B(n_397), .Y(n_741) );
BUFx3_ASAP7_75t_L g742 ( .A(n_522), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g743 ( .A1(n_628), .A2(n_640), .B(n_634), .C(n_594), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_526), .B(n_397), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_524), .A2(n_486), .B1(n_490), .B2(n_438), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_526), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_524), .A2(n_486), .B1(n_490), .B2(n_438), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_536), .Y(n_748) );
BUFx2_ASAP7_75t_L g749 ( .A(n_625), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_524), .A2(n_486), .B1(n_490), .B2(n_438), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_526), .B(n_397), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_539), .B(n_470), .Y(n_752) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_619), .Y(n_753) );
AO31x2_ASAP7_75t_L g754 ( .A1(n_535), .A2(n_570), .A3(n_569), .B(n_534), .Y(n_754) );
AO21x2_ASAP7_75t_L g755 ( .A1(n_535), .A2(n_629), .B(n_502), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_526), .B(n_524), .Y(n_756) );
AO31x2_ASAP7_75t_L g757 ( .A1(n_535), .A2(n_570), .A3(n_569), .B(n_534), .Y(n_757) );
OAI21xp5_ASAP7_75t_L g758 ( .A1(n_560), .A2(n_451), .B(n_534), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_526), .B(n_397), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_526), .B(n_397), .Y(n_760) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_536), .Y(n_761) );
OAI21x1_ASAP7_75t_L g762 ( .A1(n_580), .A2(n_502), .B(n_550), .Y(n_762) );
OAI21x1_ASAP7_75t_L g763 ( .A1(n_580), .A2(n_502), .B(n_550), .Y(n_763) );
OAI21xp5_ASAP7_75t_L g764 ( .A1(n_560), .A2(n_451), .B(n_466), .Y(n_764) );
BUFx3_ASAP7_75t_L g765 ( .A(n_670), .Y(n_765) );
OAI21xp5_ASAP7_75t_L g766 ( .A1(n_708), .A2(n_743), .B(n_703), .Y(n_766) );
BUFx2_ASAP7_75t_L g767 ( .A(n_740), .Y(n_767) );
OAI21xp5_ASAP7_75t_L g768 ( .A1(n_764), .A2(n_719), .B(n_721), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_661), .A2(n_723), .B1(n_691), .B2(n_747), .Y(n_769) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_746), .Y(n_770) );
OAI21x1_ASAP7_75t_SL g771 ( .A1(n_736), .A2(n_732), .B(n_692), .Y(n_771) );
OAI21xp5_ASAP7_75t_L g772 ( .A1(n_764), .A2(n_719), .B(n_758), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_710), .Y(n_773) );
INVx3_ASAP7_75t_L g774 ( .A(n_666), .Y(n_774) );
AO21x1_ASAP7_75t_L g775 ( .A1(n_685), .A2(n_663), .B(n_686), .Y(n_775) );
AOI21xp33_ASAP7_75t_L g776 ( .A1(n_714), .A2(n_745), .B(n_735), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_705), .Y(n_777) );
OAI21xp5_ASAP7_75t_L g778 ( .A1(n_706), .A2(n_650), .B(n_648), .Y(n_778) );
AO21x2_ASAP7_75t_L g779 ( .A1(n_762), .A2(n_763), .B(n_755), .Y(n_779) );
BUFx8_ASAP7_75t_L g780 ( .A(n_671), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_644), .Y(n_781) );
OAI21x1_ASAP7_75t_SL g782 ( .A1(n_750), .A2(n_683), .B(n_677), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_658), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_720), .Y(n_784) );
INVx1_ASAP7_75t_SL g785 ( .A(n_702), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_734), .B(n_738), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_756), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_656), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_675), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_752), .A2(n_647), .B1(n_657), .B2(n_690), .Y(n_790) );
NOR2x1_ASAP7_75t_SL g791 ( .A(n_704), .B(n_666), .Y(n_791) );
CKINVDCx6p67_ASAP7_75t_R g792 ( .A(n_753), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_741), .B(n_744), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g794 ( .A(n_674), .B(n_740), .Y(n_794) );
INVx4_ASAP7_75t_SL g795 ( .A(n_700), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_674), .A2(n_751), .B1(n_760), .B2(n_759), .Y(n_796) );
OAI211xp5_ASAP7_75t_L g797 ( .A1(n_667), .A2(n_677), .B(n_711), .C(n_660), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_645), .A2(n_717), .B1(n_718), .B2(n_678), .Y(n_798) );
INVx2_ASAP7_75t_SL g799 ( .A(n_710), .Y(n_799) );
OAI21xp5_ASAP7_75t_L g800 ( .A1(n_701), .A2(n_722), .B(n_729), .Y(n_800) );
INVx3_ASAP7_75t_L g801 ( .A(n_666), .Y(n_801) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_761), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_689), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_716), .B(n_668), .Y(n_804) );
NAND2x1_ASAP7_75t_L g805 ( .A(n_700), .B(n_696), .Y(n_805) );
OA21x2_ASAP7_75t_L g806 ( .A1(n_724), .A2(n_709), .B(n_725), .Y(n_806) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_761), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_681), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_694), .Y(n_809) );
OR2x6_ASAP7_75t_L g810 ( .A(n_749), .B(n_742), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_652), .Y(n_811) );
AO31x2_ASAP7_75t_L g812 ( .A1(n_679), .A2(n_680), .A3(n_673), .B(n_695), .Y(n_812) );
OA21x2_ASAP7_75t_L g813 ( .A1(n_725), .A2(n_682), .B(n_730), .Y(n_813) );
AND2x4_ASAP7_75t_L g814 ( .A(n_727), .B(n_664), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_662), .B(n_676), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_659), .Y(n_816) );
AO21x2_ASAP7_75t_L g817 ( .A1(n_726), .A2(n_701), .B(n_731), .Y(n_817) );
AND2x4_ASAP7_75t_L g818 ( .A(n_727), .B(n_713), .Y(n_818) );
NAND2x1p5_ASAP7_75t_L g819 ( .A(n_712), .B(n_715), .Y(n_819) );
NOR2xp33_ASAP7_75t_SL g820 ( .A(n_659), .B(n_700), .Y(n_820) );
INVx2_ASAP7_75t_SL g821 ( .A(n_713), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_688), .B(n_699), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_652), .Y(n_823) );
OR2x2_ASAP7_75t_L g824 ( .A(n_733), .B(n_646), .Y(n_824) );
NAND2x1p5_ASAP7_75t_L g825 ( .A(n_654), .B(n_684), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_669), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_728), .B(n_698), .Y(n_827) );
NAND2x1p5_ASAP7_75t_L g828 ( .A(n_654), .B(n_737), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_669), .Y(n_829) );
BUFx4f_ASAP7_75t_L g830 ( .A(n_700), .Y(n_830) );
OA21x2_ASAP7_75t_L g831 ( .A1(n_653), .A2(n_665), .B(n_655), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_669), .Y(n_832) );
OR2x2_ASAP7_75t_L g833 ( .A(n_672), .B(n_651), .Y(n_833) );
OR2x6_ASAP7_75t_L g834 ( .A(n_748), .B(n_693), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_672), .B(n_757), .Y(n_835) );
AND2x4_ASAP7_75t_L g836 ( .A(n_739), .B(n_757), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_672), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_687), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_707), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_739), .Y(n_840) );
NAND2x1p5_ASAP7_75t_L g841 ( .A(n_697), .B(n_649), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_757), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_754), .B(n_526), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_754), .B(n_625), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_705), .Y(n_845) );
AND2x4_ASAP7_75t_L g846 ( .A(n_740), .B(n_746), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_710), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_734), .B(n_526), .Y(n_848) );
INVx3_ASAP7_75t_L g849 ( .A(n_666), .Y(n_849) );
OR2x2_ASAP7_75t_L g850 ( .A(n_746), .B(n_524), .Y(n_850) );
OR2x2_ASAP7_75t_L g851 ( .A(n_746), .B(n_524), .Y(n_851) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_746), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_705), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_734), .B(n_526), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_734), .B(n_526), .Y(n_855) );
OR2x2_ASAP7_75t_L g856 ( .A(n_746), .B(n_524), .Y(n_856) );
AO21x1_ASAP7_75t_L g857 ( .A1(n_661), .A2(n_692), .B(n_613), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_708), .A2(n_743), .B(n_706), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_705), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_705), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_734), .B(n_526), .Y(n_861) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_708), .A2(n_743), .B(n_706), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_734), .B(n_526), .Y(n_863) );
A2O1A1Ixp33_ASAP7_75t_L g864 ( .A1(n_703), .A2(n_708), .B(n_743), .C(n_719), .Y(n_864) );
INVx4_ASAP7_75t_L g865 ( .A(n_670), .Y(n_865) );
OAI211xp5_ASAP7_75t_L g866 ( .A1(n_667), .A2(n_562), .B(n_454), .C(n_633), .Y(n_866) );
NAND2x1p5_ASAP7_75t_L g867 ( .A(n_671), .B(n_525), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_756), .B(n_524), .Y(n_868) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_746), .Y(n_869) );
A2O1A1Ixp33_ASAP7_75t_L g870 ( .A1(n_703), .A2(n_708), .B(n_743), .C(n_719), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_705), .Y(n_871) );
AOI21xp5_ASAP7_75t_L g872 ( .A1(n_708), .A2(n_743), .B(n_706), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_734), .B(n_526), .Y(n_873) );
BUFx2_ASAP7_75t_L g874 ( .A(n_740), .Y(n_874) );
CKINVDCx12_ASAP7_75t_R g875 ( .A(n_710), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_769), .A2(n_798), .B1(n_844), .B2(n_857), .Y(n_876) );
OR2x2_ASAP7_75t_L g877 ( .A(n_843), .B(n_777), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_777), .B(n_845), .Y(n_878) );
INVxp67_ASAP7_75t_L g879 ( .A(n_770), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_780), .Y(n_880) );
NAND2x1_ASAP7_75t_L g881 ( .A(n_839), .B(n_771), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_811), .Y(n_882) );
OAI211xp5_ASAP7_75t_L g883 ( .A1(n_866), .A2(n_790), .B(n_797), .C(n_776), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_823), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_845), .B(n_853), .Y(n_885) );
AO21x1_ASAP7_75t_SL g886 ( .A1(n_795), .A2(n_830), .B(n_820), .Y(n_886) );
AO21x2_ASAP7_75t_L g887 ( .A1(n_800), .A2(n_862), .B(n_858), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_826), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_826), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_829), .Y(n_890) );
AO21x2_ASAP7_75t_L g891 ( .A1(n_872), .A2(n_768), .B(n_772), .Y(n_891) );
OR2x2_ASAP7_75t_SL g892 ( .A(n_824), .B(n_813), .Y(n_892) );
INVx2_ASAP7_75t_SL g893 ( .A(n_830), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_840), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_829), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_842), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_796), .A2(n_782), .B1(n_860), .B2(n_853), .Y(n_897) );
OAI221xp5_ASAP7_75t_L g898 ( .A1(n_848), .A2(n_863), .B1(n_854), .B2(n_861), .C(n_855), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_859), .B(n_860), .Y(n_899) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_873), .A2(n_786), .B1(n_793), .B2(n_871), .C(n_859), .Y(n_900) );
OR2x2_ASAP7_75t_L g901 ( .A(n_871), .B(n_852), .Y(n_901) );
CKINVDCx5p33_ASAP7_75t_R g902 ( .A(n_780), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_832), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_778), .B(n_766), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_837), .Y(n_905) );
BUFx2_ASAP7_75t_L g906 ( .A(n_795), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_784), .B(n_835), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_869), .B(n_804), .Y(n_908) );
INVx5_ASAP7_75t_L g909 ( .A(n_802), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_803), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_803), .B(n_787), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_781), .B(n_850), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_827), .Y(n_913) );
AND2x2_ASAP7_75t_L g914 ( .A(n_864), .B(n_870), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_808), .Y(n_915) );
BUFx3_ASAP7_75t_L g916 ( .A(n_765), .Y(n_916) );
INVx2_ASAP7_75t_L g917 ( .A(n_806), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_808), .Y(n_918) );
AND2x4_ASAP7_75t_L g919 ( .A(n_774), .B(n_801), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_809), .Y(n_920) );
OR2x2_ASAP7_75t_L g921 ( .A(n_851), .B(n_856), .Y(n_921) );
INVx2_ASAP7_75t_L g922 ( .A(n_836), .Y(n_922) );
INVx2_ASAP7_75t_L g923 ( .A(n_836), .Y(n_923) );
INVx2_ASAP7_75t_SL g924 ( .A(n_810), .Y(n_924) );
HB1xp67_ASAP7_75t_L g925 ( .A(n_810), .Y(n_925) );
INVx2_ASAP7_75t_L g926 ( .A(n_779), .Y(n_926) );
AO21x2_ASAP7_75t_L g927 ( .A1(n_817), .A2(n_838), .B(n_775), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_833), .Y(n_928) );
BUFx2_ASAP7_75t_L g929 ( .A(n_807), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_789), .B(n_783), .Y(n_930) );
INVx3_ASAP7_75t_L g931 ( .A(n_805), .Y(n_931) );
BUFx3_ASAP7_75t_L g932 ( .A(n_865), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_834), .Y(n_933) );
AO21x2_ASAP7_75t_L g934 ( .A1(n_822), .A2(n_788), .B(n_791), .Y(n_934) );
OR2x2_ASAP7_75t_L g935 ( .A(n_815), .B(n_868), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_819), .B(n_794), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_813), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_846), .B(n_785), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_846), .B(n_767), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_849), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_792), .A2(n_814), .B1(n_874), .B2(n_816), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_814), .B(n_867), .Y(n_942) );
INVx2_ASAP7_75t_SL g943 ( .A(n_865), .Y(n_943) );
AO21x2_ASAP7_75t_L g944 ( .A1(n_818), .A2(n_841), .B(n_812), .Y(n_944) );
NOR2xp33_ASAP7_75t_L g945 ( .A(n_898), .B(n_799), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_907), .B(n_812), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_877), .B(n_818), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_905), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_905), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_907), .B(n_812), .Y(n_950) );
BUFx2_ASAP7_75t_L g951 ( .A(n_929), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_877), .B(n_825), .Y(n_952) );
AND2x4_ASAP7_75t_SL g953 ( .A(n_878), .B(n_821), .Y(n_953) );
INVx2_ASAP7_75t_SL g954 ( .A(n_909), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_904), .B(n_828), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_914), .B(n_831), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_914), .B(n_831), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_878), .B(n_773), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_897), .B(n_847), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_885), .B(n_875), .Y(n_960) );
BUFx3_ASAP7_75t_L g961 ( .A(n_909), .Y(n_961) );
OR2x2_ASAP7_75t_L g962 ( .A(n_928), .B(n_901), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_885), .B(n_899), .Y(n_963) );
BUFx2_ASAP7_75t_L g964 ( .A(n_929), .Y(n_964) );
INVx5_ASAP7_75t_L g965 ( .A(n_906), .Y(n_965) );
INVxp67_ASAP7_75t_L g966 ( .A(n_901), .Y(n_966) );
AND2x4_ASAP7_75t_L g967 ( .A(n_922), .B(n_923), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_899), .B(n_882), .Y(n_968) );
INVx3_ASAP7_75t_L g969 ( .A(n_881), .Y(n_969) );
OR2x2_ASAP7_75t_L g970 ( .A(n_928), .B(n_921), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_922), .B(n_923), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_891), .B(n_884), .Y(n_972) );
OR2x2_ASAP7_75t_L g973 ( .A(n_921), .B(n_908), .Y(n_973) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_894), .Y(n_974) );
INVx1_ASAP7_75t_SL g975 ( .A(n_936), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_884), .B(n_888), .Y(n_976) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_896), .Y(n_977) );
INVx2_ASAP7_75t_SL g978 ( .A(n_909), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_917), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_889), .B(n_890), .Y(n_980) );
INVxp67_ASAP7_75t_SL g981 ( .A(n_913), .Y(n_981) );
INVx2_ASAP7_75t_SL g982 ( .A(n_909), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_890), .B(n_895), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_910), .B(n_911), .Y(n_984) );
OR2x6_ASAP7_75t_SL g985 ( .A(n_880), .B(n_902), .Y(n_985) );
AND2x4_ASAP7_75t_L g986 ( .A(n_944), .B(n_933), .Y(n_986) );
INVxp67_ASAP7_75t_L g987 ( .A(n_913), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_876), .A2(n_900), .B1(n_935), .B2(n_879), .Y(n_988) );
NOR2xp33_ASAP7_75t_R g989 ( .A(n_880), .B(n_902), .Y(n_989) );
INVx3_ASAP7_75t_L g990 ( .A(n_931), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_910), .B(n_915), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_911), .B(n_903), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_963), .B(n_918), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_946), .B(n_891), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_963), .B(n_920), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_948), .Y(n_996) );
HB1xp67_ASAP7_75t_L g997 ( .A(n_966), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_992), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_946), .B(n_887), .Y(n_999) );
INVx2_ASAP7_75t_L g1000 ( .A(n_979), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_948), .Y(n_1001) );
HB1xp67_ASAP7_75t_L g1002 ( .A(n_966), .Y(n_1002) );
INVx1_ASAP7_75t_SL g1003 ( .A(n_989), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_949), .Y(n_1004) );
AND2x4_ASAP7_75t_SL g1005 ( .A(n_954), .B(n_978), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_946), .B(n_887), .Y(n_1006) );
AND2x4_ASAP7_75t_L g1007 ( .A(n_972), .B(n_944), .Y(n_1007) );
OR2x2_ASAP7_75t_L g1008 ( .A(n_962), .B(n_892), .Y(n_1008) );
INVx3_ASAP7_75t_L g1009 ( .A(n_969), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_950), .B(n_887), .Y(n_1010) );
HB1xp67_ASAP7_75t_L g1011 ( .A(n_951), .Y(n_1011) );
BUFx2_ASAP7_75t_L g1012 ( .A(n_981), .Y(n_1012) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_962), .B(n_892), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_950), .B(n_937), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_984), .B(n_918), .Y(n_1015) );
INVx4_ASAP7_75t_L g1016 ( .A(n_965), .Y(n_1016) );
CKINVDCx14_ASAP7_75t_R g1017 ( .A(n_985), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_945), .A2(n_934), .B1(n_935), .B2(n_944), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_950), .B(n_937), .Y(n_1019) );
NAND2x1p5_ASAP7_75t_L g1020 ( .A(n_965), .B(n_906), .Y(n_1020) );
OR2x2_ASAP7_75t_L g1021 ( .A(n_970), .B(n_912), .Y(n_1021) );
OR2x2_ASAP7_75t_L g1022 ( .A(n_970), .B(n_926), .Y(n_1022) );
INVx2_ASAP7_75t_SL g1023 ( .A(n_965), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_984), .B(n_920), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g1025 ( .A(n_964), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_971), .B(n_927), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_988), .A2(n_934), .B1(n_924), .B2(n_925), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_971), .B(n_927), .Y(n_1028) );
OR2x2_ASAP7_75t_L g1029 ( .A(n_973), .B(n_926), .Y(n_1029) );
INVx1_ASAP7_75t_SL g1030 ( .A(n_985), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_992), .B(n_915), .Y(n_1031) );
AND2x4_ASAP7_75t_L g1032 ( .A(n_1007), .B(n_956), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_996), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_998), .B(n_968), .Y(n_1034) );
NAND2xp5_ASAP7_75t_SL g1035 ( .A(n_1030), .B(n_965), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_999), .B(n_957), .Y(n_1036) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_1007), .B(n_957), .Y(n_1037) );
NOR2x1p5_ASAP7_75t_L g1038 ( .A(n_1016), .B(n_981), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_997), .B(n_968), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_999), .B(n_972), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_996), .Y(n_1041) );
AND2x4_ASAP7_75t_L g1042 ( .A(n_1007), .B(n_986), .Y(n_1042) );
INVx2_ASAP7_75t_L g1043 ( .A(n_1000), .Y(n_1043) );
NAND2xp5_ASAP7_75t_SL g1044 ( .A(n_1016), .B(n_965), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1006), .B(n_971), .Y(n_1045) );
NAND2xp5_ASAP7_75t_SL g1046 ( .A(n_1016), .B(n_965), .Y(n_1046) );
INVx3_ASAP7_75t_SL g1047 ( .A(n_1005), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_1006), .B(n_976), .Y(n_1048) );
OR2x2_ASAP7_75t_L g1049 ( .A(n_1029), .B(n_973), .Y(n_1049) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_1029), .B(n_974), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1001), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_1010), .B(n_976), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1001), .Y(n_1053) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_1008), .B(n_974), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_1002), .B(n_987), .Y(n_1055) );
OAI22xp33_ASAP7_75t_L g1056 ( .A1(n_1020), .A2(n_965), .B1(n_959), .B2(n_954), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1004), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_1010), .B(n_980), .Y(n_1058) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_1008), .B(n_977), .Y(n_1059) );
OR2x2_ASAP7_75t_L g1060 ( .A(n_1013), .B(n_977), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_993), .B(n_987), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_994), .B(n_980), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_994), .B(n_983), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1014), .B(n_983), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1014), .B(n_986), .Y(n_1065) );
OR2x2_ASAP7_75t_L g1066 ( .A(n_1013), .B(n_975), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_995), .B(n_988), .Y(n_1067) );
NOR2x1p5_ASAP7_75t_L g1068 ( .A(n_1009), .B(n_961), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1019), .B(n_986), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1019), .B(n_986), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1026), .B(n_967), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1040), .B(n_1026), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_1036), .B(n_1031), .Y(n_1073) );
OAI22xp33_ASAP7_75t_SL g1074 ( .A1(n_1047), .A2(n_985), .B1(n_1020), .B2(n_1023), .Y(n_1074) );
BUFx3_ASAP7_75t_L g1075 ( .A(n_1047), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_1036), .B(n_1015), .Y(n_1076) );
OR2x2_ASAP7_75t_L g1077 ( .A(n_1049), .B(n_1022), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1040), .B(n_1028), .Y(n_1078) );
NAND2xp5_ASAP7_75t_SL g1079 ( .A(n_1047), .B(n_1023), .Y(n_1079) );
OAI21xp33_ASAP7_75t_SL g1080 ( .A1(n_1038), .A2(n_1003), .B(n_1017), .Y(n_1080) );
INVx1_ASAP7_75t_SL g1081 ( .A(n_1049), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1048), .B(n_1052), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_1064), .B(n_1024), .Y(n_1083) );
NAND2xp33_ASAP7_75t_SL g1084 ( .A(n_1038), .B(n_1012), .Y(n_1084) );
OR2x2_ASAP7_75t_L g1085 ( .A(n_1039), .B(n_1022), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1033), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1041), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1041), .Y(n_1088) );
NOR2xp33_ASAP7_75t_L g1089 ( .A(n_1067), .B(n_958), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1064), .B(n_1028), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1051), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1051), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1053), .Y(n_1093) );
AOI21xp5_ASAP7_75t_L g1094 ( .A1(n_1044), .A2(n_1005), .B(n_1020), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1053), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_1054), .B(n_1012), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1057), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1062), .B(n_1021), .Y(n_1098) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1043), .Y(n_1099) );
INVx1_ASAP7_75t_SL g1100 ( .A(n_1075), .Y(n_1100) );
OAI21xp5_ASAP7_75t_L g1101 ( .A1(n_1080), .A2(n_1046), .B(n_1027), .Y(n_1101) );
AND2x4_ASAP7_75t_L g1102 ( .A(n_1075), .B(n_1068), .Y(n_1102) );
AOI221xp5_ASAP7_75t_L g1103 ( .A1(n_1089), .A2(n_1055), .B1(n_1061), .B2(n_1034), .C(n_1048), .Y(n_1103) );
AOI21xp33_ASAP7_75t_L g1104 ( .A1(n_1074), .A2(n_959), .B(n_943), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g1105 ( .A1(n_1081), .A2(n_1058), .B1(n_1052), .B2(n_1062), .C(n_1063), .Y(n_1105) );
NOR2xp33_ASAP7_75t_L g1106 ( .A(n_1098), .B(n_916), .Y(n_1106) );
INVxp67_ASAP7_75t_L g1107 ( .A(n_1079), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1077), .Y(n_1108) );
OAI22xp5_ASAP7_75t_L g1109 ( .A1(n_1079), .A2(n_1068), .B1(n_1018), .B2(n_1056), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1110 ( .A(n_1082), .B(n_1063), .Y(n_1110) );
INVx1_ASAP7_75t_SL g1111 ( .A(n_1096), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1082), .B(n_1058), .Y(n_1112) );
OAI22xp33_ASAP7_75t_L g1113 ( .A1(n_1094), .A2(n_1035), .B1(n_1054), .B2(n_1059), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1072), .B(n_1045), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1078), .B(n_1032), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1078), .B(n_1045), .Y(n_1116) );
OAI21x1_ASAP7_75t_SL g1117 ( .A1(n_1101), .A2(n_1084), .B(n_1083), .Y(n_1117) );
OAI221xp5_ASAP7_75t_L g1118 ( .A1(n_1101), .A2(n_883), .B1(n_1066), .B2(n_1085), .C(n_941), .Y(n_1118) );
OAI21xp33_ASAP7_75t_SL g1119 ( .A1(n_1105), .A2(n_1090), .B(n_1076), .Y(n_1119) );
AOI21xp5_ASAP7_75t_SL g1120 ( .A1(n_1109), .A2(n_932), .B(n_916), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1108), .Y(n_1121) );
OAI211xp5_ASAP7_75t_L g1122 ( .A1(n_1104), .A2(n_960), .B(n_943), .C(n_1066), .Y(n_1122) );
NOR2xp33_ASAP7_75t_L g1123 ( .A(n_1100), .B(n_1073), .Y(n_1123) );
AOI221xp5_ASAP7_75t_L g1124 ( .A1(n_1103), .A2(n_1088), .B1(n_1087), .B2(n_1097), .C(n_1095), .Y(n_1124) );
AOI221xp5_ASAP7_75t_L g1125 ( .A1(n_1109), .A2(n_1086), .B1(n_1093), .B2(n_1092), .C(n_1091), .Y(n_1125) );
AOI211xp5_ASAP7_75t_L g1126 ( .A1(n_1113), .A2(n_1060), .B(n_1059), .C(n_1032), .Y(n_1126) );
OAI22xp33_ASAP7_75t_L g1127 ( .A1(n_1107), .A2(n_1060), .B1(n_1050), .B2(n_1011), .Y(n_1127) );
OAI221xp5_ASAP7_75t_SL g1128 ( .A1(n_1111), .A2(n_1021), .B1(n_1069), .B2(n_1070), .C(n_1065), .Y(n_1128) );
NOR2xp33_ASAP7_75t_L g1129 ( .A(n_1106), .B(n_1037), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1110), .B(n_1037), .Y(n_1130) );
NOR3xp33_ASAP7_75t_SL g1131 ( .A(n_1112), .B(n_938), .C(n_942), .Y(n_1131) );
NOR2xp33_ASAP7_75t_L g1132 ( .A(n_1114), .B(n_924), .Y(n_1132) );
NOR2xp33_ASAP7_75t_L g1133 ( .A(n_1116), .B(n_1042), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1115), .B(n_1071), .Y(n_1134) );
NOR3xp33_ASAP7_75t_L g1135 ( .A(n_1102), .B(n_939), .C(n_990), .Y(n_1135) );
OAI211xp5_ASAP7_75t_SL g1136 ( .A1(n_1102), .A2(n_952), .B(n_975), .C(n_947), .Y(n_1136) );
AOI221xp5_ASAP7_75t_L g1137 ( .A1(n_1125), .A2(n_1119), .B1(n_1117), .B2(n_1118), .C(n_1124), .Y(n_1137) );
NAND3xp33_ASAP7_75t_L g1138 ( .A(n_1126), .B(n_1120), .C(n_1122), .Y(n_1138) );
OAI211xp5_ASAP7_75t_L g1139 ( .A1(n_1135), .A2(n_1131), .B(n_1128), .C(n_1123), .Y(n_1139) );
NAND3xp33_ASAP7_75t_SL g1140 ( .A(n_1129), .B(n_1121), .C(n_1130), .Y(n_1140) );
OAI211xp5_ASAP7_75t_L g1141 ( .A1(n_1132), .A2(n_1136), .B(n_1133), .C(n_1134), .Y(n_1141) );
AOI21xp5_ASAP7_75t_L g1142 ( .A1(n_1127), .A2(n_953), .B(n_954), .Y(n_1142) );
AND3x1_ASAP7_75t_L g1143 ( .A(n_1137), .B(n_893), .C(n_955), .Y(n_1143) );
OR2x2_ASAP7_75t_L g1144 ( .A(n_1138), .B(n_1050), .Y(n_1144) );
NAND4xp25_ASAP7_75t_SL g1145 ( .A(n_1139), .B(n_955), .C(n_952), .D(n_947), .Y(n_1145) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_1140), .B(n_1099), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1144), .B(n_1141), .Y(n_1147) );
NAND2xp5_ASAP7_75t_SL g1148 ( .A(n_1143), .B(n_1142), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1146), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1149), .Y(n_1150) );
XNOR2xp5_ASAP7_75t_L g1151 ( .A(n_1147), .B(n_1145), .Y(n_1151) );
NAND2xp5_ASAP7_75t_SL g1152 ( .A(n_1150), .B(n_1148), .Y(n_1152) );
AOI22xp5_ASAP7_75t_L g1153 ( .A1(n_1151), .A2(n_934), .B1(n_893), .B2(n_953), .Y(n_1153) );
AOI22xp5_ASAP7_75t_L g1154 ( .A1(n_1152), .A2(n_930), .B1(n_978), .B2(n_982), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1153), .B(n_1099), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_1155), .A2(n_1025), .B1(n_982), .B2(n_961), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_1156), .A2(n_1154), .B1(n_886), .B2(n_961), .Y(n_1157) );
OAI21x1_ASAP7_75t_SL g1158 ( .A1(n_1157), .A2(n_886), .B(n_991), .Y(n_1158) );
AOI21xp5_ASAP7_75t_L g1159 ( .A1(n_1158), .A2(n_919), .B(n_940), .Y(n_1159) );
endmodule