module fake_jpeg_2772_n_192 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_192);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_13),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_SL g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_67),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_71),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_62),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_56),
.B1(n_62),
.B2(n_45),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_83),
.B1(n_73),
.B2(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_61),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_56),
.B1(n_62),
.B2(n_51),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_99),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_54),
.B1(n_46),
.B2(n_59),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_90),
.B1(n_50),
.B2(n_63),
.Y(n_103)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_98),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_54),
.B1(n_59),
.B2(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_96),
.Y(n_108)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_95),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_100),
.B1(n_60),
.B2(n_3),
.Y(n_113)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_73),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_57),
.B1(n_43),
.B2(n_63),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_47),
.B(n_53),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_118),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_112),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_78),
.B1(n_63),
.B2(n_60),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_111),
.B1(n_6),
.B2(n_8),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_86),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_60),
.B1(n_1),
.B2(n_2),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_0),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_116),
.B(n_6),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_19),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_10),
.C(n_11),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_87),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_108),
.B(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_129),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_107),
.B(n_22),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_12),
.C(n_13),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_14),
.Y(n_146)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_8),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_130),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_9),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_103),
.B1(n_105),
.B2(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_136),
.Y(n_152)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_9),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_34),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_111),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_12),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_145),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_10),
.B(n_11),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_144),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_15),
.B(n_16),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_149),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_20),
.C(n_23),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_137),
.C(n_131),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_139),
.A2(n_24),
.B(n_26),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_151),
.B(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_132),
.CI(n_125),
.CON(n_161),
.SN(n_161)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_168),
.Y(n_177)
);

NOR2xp67_ASAP7_75t_R g162 ( 
.A(n_154),
.B(n_145),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_162),
.B(n_164),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_143),
.B1(n_138),
.B2(n_147),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_171),
.A2(n_173),
.B1(n_161),
.B2(n_169),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_163),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_148),
.C(n_165),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_164),
.A2(n_151),
.B(n_142),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_150),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_175),
.B(n_152),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_181),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_184),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_170),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_179),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_185),
.B(n_182),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_37),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_39),
.B(n_40),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g191 ( 
.A(n_190),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_172),
.B1(n_144),
.B2(n_166),
.Y(n_192)
);


endmodule