module real_aes_9028_n_254 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_254);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_254;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_519;
wire n_815;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_725;
wire n_455;
wire n_504;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_449;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_809;
wire n_482;
wire n_679;
wire n_633;
wire n_520;
wire n_472;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_741;
wire n_314;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_668;
wire n_797;
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_0), .A2(n_196), .B1(n_298), .B2(n_361), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_1), .Y(n_523) );
AOI222xp33_ASAP7_75t_L g337 ( .A1(n_2), .A2(n_82), .B1(n_238), .B2(n_338), .C1(n_341), .C2(n_345), .Y(n_337) );
INVx1_ASAP7_75t_L g350 ( .A(n_3), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_4), .A2(n_57), .B1(n_330), .B2(n_406), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_5), .B(n_324), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_6), .A2(n_13), .B1(n_429), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_7), .A2(n_119), .B1(n_424), .B2(n_426), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_8), .A2(n_161), .B1(n_381), .B2(n_505), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_9), .A2(n_139), .B1(n_460), .B2(n_461), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_10), .A2(n_47), .B1(n_428), .B2(n_429), .Y(n_427) );
AOI222xp33_ASAP7_75t_L g677 ( .A1(n_11), .A2(n_116), .B1(n_204), .B2(n_475), .C1(n_678), .C2(n_679), .Y(n_677) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_12), .A2(n_52), .B1(n_507), .B2(n_509), .Y(n_506) );
AOI222xp33_ASAP7_75t_L g593 ( .A1(n_14), .A2(n_84), .B1(n_129), .B2(n_403), .C1(n_594), .C2(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_15), .B(n_468), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g694 ( .A1(n_16), .A2(n_157), .B1(n_312), .B2(n_652), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_17), .A2(n_114), .B1(n_556), .B2(n_720), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_18), .Y(n_385) );
AO22x2_ASAP7_75t_L g278 ( .A1(n_19), .A2(n_86), .B1(n_279), .B2(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g752 ( .A(n_19), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_20), .B(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_21), .A2(n_190), .B1(n_481), .B2(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_22), .A2(n_252), .B1(n_293), .B2(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_23), .A2(n_136), .B1(n_651), .B2(n_775), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_24), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_25), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_26), .A2(n_253), .B1(n_363), .B2(n_460), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_27), .A2(n_150), .B1(n_354), .B2(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g398 ( .A(n_28), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_29), .A2(n_237), .B1(n_355), .B2(n_454), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_30), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_31), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_32), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_33), .A2(n_230), .B1(n_293), .B2(n_298), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_34), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_35), .B(n_442), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_36), .Y(n_808) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_37), .A2(n_178), .B1(n_476), .B2(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_38), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_39), .Y(n_546) );
INVx1_ASAP7_75t_L g448 ( .A(n_40), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_41), .A2(n_163), .B1(n_330), .B2(n_476), .Y(n_691) );
AO22x2_ASAP7_75t_L g282 ( .A1(n_42), .A2(n_87), .B1(n_279), .B2(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g753 ( .A(n_42), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_43), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_44), .A2(n_135), .B1(n_710), .B2(n_711), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_45), .Y(n_730) );
INVx1_ASAP7_75t_L g760 ( .A(n_46), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_48), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_49), .A2(n_81), .B1(n_428), .B2(n_587), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_50), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_51), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_53), .A2(n_58), .B1(n_485), .B2(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_54), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_55), .B(n_811), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_56), .A2(n_118), .B1(n_525), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_59), .A2(n_69), .B1(n_293), .B2(n_426), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_60), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_61), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_62), .A2(n_210), .B1(n_272), .B2(n_289), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_63), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_64), .A2(n_245), .B1(n_357), .B2(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_65), .A2(n_140), .B1(n_381), .B2(n_471), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_66), .A2(n_183), .B1(n_312), .B2(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_67), .A2(n_191), .B1(n_460), .B2(n_654), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_68), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_70), .A2(n_182), .B1(n_328), .B2(n_541), .Y(n_727) );
XNOR2x2_ASAP7_75t_L g268 ( .A(n_71), .B(n_269), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_72), .Y(n_640) );
AO22x2_ASAP7_75t_L g632 ( .A1(n_73), .A2(n_633), .B1(n_656), .B2(n_657), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_73), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_74), .A2(n_153), .B1(n_623), .B2(n_625), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_75), .A2(n_219), .B1(n_651), .B2(n_652), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_76), .A2(n_101), .B1(n_515), .B2(n_517), .Y(n_514) );
AOI211xp5_ASAP7_75t_L g534 ( .A1(n_77), .A2(n_403), .B(n_535), .C(n_543), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_78), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_79), .A2(n_212), .B1(n_507), .B2(n_591), .Y(n_590) );
AOI22xp5_ASAP7_75t_SL g353 ( .A1(n_80), .A2(n_138), .B1(n_354), .B2(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g462 ( .A(n_83), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_85), .A2(n_225), .B1(n_604), .B2(n_605), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_88), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_89), .Y(n_708) );
INVx1_ASAP7_75t_L g261 ( .A(n_90), .Y(n_261) );
AOI211xp5_ASAP7_75t_L g254 ( .A1(n_91), .A2(n_255), .B(n_263), .C(n_754), .Y(n_254) );
AOI22xp5_ASAP7_75t_SL g391 ( .A1(n_92), .A2(n_392), .B1(n_434), .B2(n_435), .Y(n_391) );
INVx1_ASAP7_75t_L g435 ( .A(n_92), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_93), .A2(n_122), .B1(n_304), .B2(n_306), .Y(n_303) );
INVx1_ASAP7_75t_L g488 ( .A(n_94), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_95), .A2(n_127), .B1(n_461), .B2(n_553), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_96), .Y(n_706) );
AOI22xp5_ASAP7_75t_SL g360 ( .A1(n_97), .A2(n_224), .B1(n_361), .B2(n_363), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_98), .A2(n_173), .B1(n_345), .B2(n_381), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_99), .A2(n_192), .B1(n_461), .B2(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g258 ( .A(n_100), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_102), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_103), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_104), .A2(n_137), .B1(n_341), .B2(n_346), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_105), .A2(n_175), .B1(n_312), .B2(n_315), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_106), .B(n_444), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_107), .A2(n_228), .B1(n_456), .B2(n_517), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_108), .A2(n_205), .B1(n_341), .B2(n_471), .Y(n_470) );
AOI211xp5_ASAP7_75t_L g518 ( .A1(n_109), .A2(n_519), .B(n_520), .C(n_528), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_110), .A2(n_158), .B1(n_290), .B2(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_111), .B(n_442), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_112), .A2(n_167), .B1(n_480), .B2(n_481), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_113), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_115), .B(n_629), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_117), .Y(n_621) );
INVx1_ASAP7_75t_L g473 ( .A(n_120), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_121), .B(n_444), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_123), .A2(n_198), .B1(n_426), .B2(n_802), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_124), .A2(n_220), .B1(n_486), .B2(n_526), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g771 ( .A1(n_125), .A2(n_246), .B1(n_306), .B2(n_458), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_126), .A2(n_200), .B1(n_505), .B2(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_128), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_130), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_131), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_132), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_133), .B(n_324), .Y(n_539) );
INVx2_ASAP7_75t_L g262 ( .A(n_134), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_141), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_142), .Y(n_806) );
INVx1_ASAP7_75t_L g767 ( .A(n_143), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_144), .A2(n_217), .B1(n_334), .B2(n_505), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_145), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_146), .A2(n_195), .B1(n_328), .B2(n_333), .Y(n_327) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_147), .Y(n_532) );
AND2x6_ASAP7_75t_L g257 ( .A(n_148), .B(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_148), .Y(n_746) );
AO22x2_ASAP7_75t_L g286 ( .A1(n_149), .A2(n_216), .B1(n_279), .B2(n_283), .Y(n_286) );
INVx1_ASAP7_75t_L g768 ( .A(n_151), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_152), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_154), .A2(n_236), .B1(n_357), .B2(n_458), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_155), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_156), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_159), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g457 ( .A1(n_160), .A2(n_240), .B1(n_354), .B2(n_458), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_162), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_164), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_165), .A2(n_250), .B1(n_315), .B2(n_654), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_166), .A2(n_174), .B1(n_405), .B2(n_407), .Y(n_404) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_168), .A2(n_187), .B1(n_485), .B2(n_486), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_169), .A2(n_702), .B1(n_735), .B2(n_736), .Y(n_701) );
INVx1_ASAP7_75t_L g735 ( .A(n_169), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_170), .A2(n_203), .B1(n_420), .B2(n_422), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_171), .A2(n_239), .B1(n_480), .B2(n_517), .Y(n_655) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_172), .A2(n_233), .B1(n_363), .B2(n_481), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_176), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_177), .A2(n_206), .B1(n_345), .B2(n_381), .Y(n_765) );
AO22x2_ASAP7_75t_L g288 ( .A1(n_179), .A2(n_232), .B1(n_279), .B2(n_280), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_180), .A2(n_243), .B1(n_475), .B2(n_476), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_181), .A2(n_208), .B1(n_519), .B2(n_607), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_184), .A2(n_207), .B1(n_306), .B2(n_432), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_185), .A2(n_234), .B1(n_548), .B2(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g566 ( .A(n_186), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_188), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_189), .A2(n_201), .B1(n_525), .B2(n_583), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_193), .A2(n_247), .B1(n_408), .B2(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g395 ( .A(n_194), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_197), .B(n_442), .Y(n_441) );
AOI22xp33_ASAP7_75t_SL g697 ( .A1(n_199), .A2(n_235), .B1(n_560), .B2(n_649), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_202), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_209), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_211), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_213), .Y(n_561) );
AOI22xp33_ASAP7_75t_SL g455 ( .A1(n_214), .A2(n_222), .B1(n_426), .B2(n_456), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_215), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_216), .B(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_218), .B(n_444), .Y(n_688) );
INVx1_ASAP7_75t_L g763 ( .A(n_221), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_223), .Y(n_813) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_226), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_227), .A2(n_599), .B1(n_600), .B2(n_631), .Y(n_598) );
INVx1_ASAP7_75t_L g631 ( .A(n_227), .Y(n_631) );
INVx1_ASAP7_75t_L g761 ( .A(n_229), .Y(n_761) );
XNOR2xp5_ASAP7_75t_L g493 ( .A(n_231), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g749 ( .A(n_232), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_241), .Y(n_374) );
INVx1_ASAP7_75t_L g279 ( .A(n_242), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_242), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_244), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_244), .A2(n_787), .B1(n_791), .B2(n_815), .Y(n_790) );
OA22x2_ASAP7_75t_L g575 ( .A1(n_248), .A2(n_576), .B1(n_577), .B2(n_596), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_248), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_249), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_251), .A2(n_756), .B1(n_778), .B2(n_779), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_251), .Y(n_778) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_257), .B(n_259), .Y(n_256) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_258), .Y(n_745) );
OA21x2_ASAP7_75t_L g785 ( .A1(n_259), .A2(n_744), .B(n_786), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_662), .B1(n_739), .B2(n_740), .C(n_741), .Y(n_263) );
INVx1_ASAP7_75t_L g739 ( .A(n_264), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_491), .B1(n_660), .B2(n_661), .Y(n_264) );
INVx1_ASAP7_75t_L g660 ( .A(n_265), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B1(n_388), .B2(n_389), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OAI22xp5_ASAP7_75t_SL g267 ( .A1(n_268), .A2(n_348), .B1(n_386), .B2(n_387), .Y(n_267) );
INVx1_ASAP7_75t_L g386 ( .A(n_268), .Y(n_386) );
NAND4xp75_ASAP7_75t_L g269 ( .A(n_270), .B(n_302), .C(n_318), .D(n_337), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_292), .Y(n_270) );
INVx2_ASAP7_75t_L g705 ( .A(n_272), .Y(n_705) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx5_ASAP7_75t_SL g458 ( .A(n_273), .Y(n_458) );
INVx2_ASAP7_75t_SL g480 ( .A(n_273), .Y(n_480) );
INVx11_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx11_ASAP7_75t_L g362 ( .A(n_274), .Y(n_362) );
AND2x6_ASAP7_75t_L g274 ( .A(n_275), .B(n_284), .Y(n_274) );
AND2x4_ASAP7_75t_L g326 ( .A(n_275), .B(n_297), .Y(n_326) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g377 ( .A(n_276), .B(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_282), .Y(n_276) );
AND2x2_ASAP7_75t_L g291 ( .A(n_277), .B(n_282), .Y(n_291) );
AND2x2_ASAP7_75t_L g295 ( .A(n_277), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g332 ( .A(n_278), .B(n_286), .Y(n_332) );
AND2x2_ASAP7_75t_L g336 ( .A(n_278), .B(n_282), .Y(n_336) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g283 ( .A(n_281), .Y(n_283) );
INVx2_ASAP7_75t_L g296 ( .A(n_282), .Y(n_296) );
INVx1_ASAP7_75t_L g317 ( .A(n_282), .Y(n_317) );
AND2x4_ASAP7_75t_L g290 ( .A(n_284), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g305 ( .A(n_284), .B(n_295), .Y(n_305) );
AND2x6_ASAP7_75t_L g340 ( .A(n_284), .B(n_336), .Y(n_340) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
AND2x2_ASAP7_75t_L g297 ( .A(n_285), .B(n_288), .Y(n_297) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_286), .B(n_288), .Y(n_301) );
AND2x2_ASAP7_75t_L g309 ( .A(n_286), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g310 ( .A(n_288), .Y(n_310) );
INVx1_ASAP7_75t_L g344 ( .A(n_288), .Y(n_344) );
INVx3_ASAP7_75t_L g776 ( .A(n_289), .Y(n_776) );
BUFx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx6_ASAP7_75t_L g430 ( .A(n_290), .Y(n_430) );
BUFx3_ASAP7_75t_L g485 ( .A(n_290), .Y(n_485) );
BUFx3_ASAP7_75t_L g649 ( .A(n_290), .Y(n_649) );
AND2x2_ASAP7_75t_L g314 ( .A(n_291), .B(n_309), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_291), .B(n_297), .Y(n_322) );
AND2x6_ASAP7_75t_L g445 ( .A(n_291), .B(n_297), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_291), .B(n_309), .Y(n_522) );
INVx4_ASAP7_75t_L g554 ( .A(n_293), .Y(n_554) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g421 ( .A(n_294), .Y(n_421) );
BUFx3_ASAP7_75t_L g456 ( .A(n_294), .Y(n_456) );
BUFx3_ASAP7_75t_L g516 ( .A(n_294), .Y(n_516) );
BUFx3_ASAP7_75t_L g654 ( .A(n_294), .Y(n_654) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
AND2x4_ASAP7_75t_L g299 ( .A(n_295), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g308 ( .A(n_295), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_295), .B(n_309), .Y(n_569) );
AND2x2_ASAP7_75t_L g343 ( .A(n_296), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g366 ( .A(n_296), .Y(n_366) );
INVx1_ASAP7_75t_L g378 ( .A(n_297), .Y(n_378) );
INVx1_ASAP7_75t_L g717 ( .A(n_298), .Y(n_717) );
BUFx2_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g363 ( .A(n_299), .Y(n_363) );
BUFx2_ASAP7_75t_SL g422 ( .A(n_299), .Y(n_422) );
BUFx2_ASAP7_75t_L g461 ( .A(n_299), .Y(n_461) );
BUFx3_ASAP7_75t_L g517 ( .A(n_299), .Y(n_517) );
BUFx3_ASAP7_75t_L g607 ( .A(n_299), .Y(n_607) );
AND2x2_ASAP7_75t_L g365 ( .A(n_300), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x6_ASAP7_75t_L g316 ( .A(n_301), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_311), .Y(n_302) );
INVx3_ASAP7_75t_L g433 ( .A(n_304), .Y(n_433) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_304), .Y(n_565) );
BUFx3_ASAP7_75t_L g587 ( .A(n_304), .Y(n_587) );
BUFx3_ASAP7_75t_L g710 ( .A(n_304), .Y(n_710) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g358 ( .A(n_305), .Y(n_358) );
BUFx2_ASAP7_75t_SL g519 ( .A(n_305), .Y(n_519) );
BUFx4f_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g712 ( .A(n_307), .Y(n_712) );
BUFx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx3_ASAP7_75t_L g354 ( .A(n_308), .Y(n_354) );
BUFx3_ASAP7_75t_L g481 ( .A(n_308), .Y(n_481) );
INVx1_ASAP7_75t_L g335 ( .A(n_310), .Y(n_335) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_312), .Y(n_802) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx3_ASAP7_75t_L g355 ( .A(n_313), .Y(n_355) );
BUFx3_ASAP7_75t_L g425 ( .A(n_313), .Y(n_425) );
INVx5_ASAP7_75t_L g486 ( .A(n_313), .Y(n_486) );
INVx4_ASAP7_75t_L g584 ( .A(n_313), .Y(n_584) );
INVx2_ASAP7_75t_L g651 ( .A(n_313), .Y(n_651) );
INVx8_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g426 ( .A(n_316), .Y(n_426) );
INVx6_ASAP7_75t_SL g526 ( .A(n_316), .Y(n_526) );
INVx1_ASAP7_75t_SL g556 ( .A(n_316), .Y(n_556) );
INVx1_ASAP7_75t_L g331 ( .A(n_317), .Y(n_331) );
OA211x2_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B(n_323), .C(n_327), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_320), .A2(n_396), .B1(n_805), .B2(n_806), .Y(n_804) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g369 ( .A(n_321), .Y(n_369) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g399 ( .A(n_322), .Y(n_399) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g442 ( .A(n_325), .Y(n_442) );
INVx5_ASAP7_75t_L g508 ( .A(n_325), .Y(n_508) );
INVx2_ASAP7_75t_L g690 ( .A(n_325), .Y(n_690) );
INVx4_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx3_ASAP7_75t_L g471 ( .A(n_330), .Y(n_471) );
BUFx2_ASAP7_75t_L g505 ( .A(n_330), .Y(n_505) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
AND2x4_ASAP7_75t_L g342 ( .A(n_332), .B(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g346 ( .A(n_332), .B(n_347), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g373 ( .A(n_332), .B(n_366), .Y(n_373) );
BUFx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_334), .Y(n_381) );
BUFx2_ASAP7_75t_SL g451 ( .A(n_334), .Y(n_451) );
BUFx3_ASAP7_75t_L g476 ( .A(n_334), .Y(n_476) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g417 ( .A(n_335), .Y(n_417) );
INVx1_ASAP7_75t_L g416 ( .A(n_336), .Y(n_416) );
INVx4_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI22xp5_ASAP7_75t_SL g382 ( .A1(n_339), .A2(n_383), .B1(n_384), .B2(n_385), .Y(n_382) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_339), .A2(n_621), .B(n_622), .Y(n_620) );
INVx4_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx3_ASAP7_75t_L g403 ( .A(n_340), .Y(n_403) );
INVx2_ASAP7_75t_L g449 ( .A(n_340), .Y(n_449) );
INVx2_ASAP7_75t_L g497 ( .A(n_340), .Y(n_497) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_340), .Y(n_678) );
INVx2_ASAP7_75t_SL g731 ( .A(n_340), .Y(n_731) );
INVx2_ASAP7_75t_L g384 ( .A(n_341), .Y(n_384) );
INVx4_ASAP7_75t_L g624 ( .A(n_341), .Y(n_624) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_342), .Y(n_406) );
BUFx4f_ASAP7_75t_SL g594 ( .A(n_342), .Y(n_594) );
BUFx2_ASAP7_75t_L g642 ( .A(n_342), .Y(n_642) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_342), .Y(n_679) );
INVx1_ASAP7_75t_L g347 ( .A(n_344), .Y(n_347) );
INVx1_ASAP7_75t_L g501 ( .A(n_345), .Y(n_501) );
BUFx4f_ASAP7_75t_L g625 ( .A(n_345), .Y(n_625) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_346), .Y(n_408) );
BUFx12f_ASAP7_75t_L g475 ( .A(n_346), .Y(n_475) );
INVx1_ASAP7_75t_SL g387 ( .A(n_348), .Y(n_387) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
XNOR2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
NAND3x1_ASAP7_75t_SL g351 ( .A(n_352), .B(n_359), .C(n_367), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_356), .Y(n_352) );
BUFx2_ASAP7_75t_L g513 ( .A(n_354), .Y(n_513) );
INVx1_ASAP7_75t_L g581 ( .A(n_354), .Y(n_581) );
INVx3_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx3_ASAP7_75t_L g460 ( .A(n_358), .Y(n_460) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
INVx1_ASAP7_75t_L g530 ( .A(n_361), .Y(n_530) );
INVx4_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_SL g428 ( .A(n_362), .Y(n_428) );
INVx3_ASAP7_75t_L g560 ( .A(n_362), .Y(n_560) );
NOR3xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_375), .C(n_382), .Y(n_367) );
OAI22xp5_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_370), .B1(n_371), .B2(n_374), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_369), .A2(n_636), .B1(n_637), .B2(n_638), .Y(n_635) );
INVx3_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g645 ( .A(n_372), .Y(n_645) );
INVx4_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx3_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_373), .A2(n_545), .B1(n_767), .B2(n_768), .Y(n_766) );
OAI21xp5_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_379), .B(n_380), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_376), .A2(n_725), .B1(n_760), .B2(n_761), .Y(n_759) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g397 ( .A(n_377), .Y(n_397) );
INVx1_ASAP7_75t_SL g542 ( .A(n_381), .Y(n_542) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OA22x2_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_436), .B1(n_489), .B2(n_490), .Y(n_390) );
INVx1_ASAP7_75t_L g489 ( .A(n_391), .Y(n_489) );
INVx2_ASAP7_75t_SL g434 ( .A(n_392), .Y(n_434) );
AND2x2_ASAP7_75t_SL g392 ( .A(n_393), .B(n_418), .Y(n_392) );
NOR3xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_400), .C(n_409), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_398), .B2(n_399), .Y(n_394) );
OAI221xp5_ASAP7_75t_SL g723 ( .A1(n_396), .A2(n_724), .B1(n_725), .B2(n_726), .C(n_727), .Y(n_723) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g637 ( .A(n_397), .Y(n_637) );
INVx2_ASAP7_75t_L g538 ( .A(n_399), .Y(n_538) );
OA211x2_ASAP7_75t_L g673 ( .A1(n_399), .A2(n_674), .B(n_675), .C(n_676), .Y(n_673) );
BUFx3_ASAP7_75t_L g725 ( .A(n_399), .Y(n_725) );
OAI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B(n_404), .Y(n_400) );
OAI21xp33_ASAP7_75t_L g639 ( .A1(n_402), .A2(n_640), .B(n_641), .Y(n_639) );
INVx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_SL g499 ( .A(n_405), .Y(n_499) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g545 ( .A(n_406), .Y(n_545) );
BUFx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g733 ( .A(n_408), .Y(n_733) );
BUFx2_ASAP7_75t_L g811 ( .A(n_408), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_412), .B2(n_413), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_413), .A2(n_645), .B1(n_813), .B2(n_814), .Y(n_812) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
CKINVDCx16_ASAP7_75t_R g414 ( .A(n_415), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_415), .A2(n_644), .B1(n_645), .B2(n_646), .Y(n_643) );
OR2x6_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
AND4x1_ASAP7_75t_L g418 ( .A(n_419), .B(n_423), .C(n_427), .D(n_431), .Y(n_418) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g454 ( .A(n_430), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_430), .A2(n_558), .B1(n_559), .B2(n_561), .Y(n_557) );
INVx3_ASAP7_75t_L g671 ( .A(n_430), .Y(n_671) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI221xp5_ASAP7_75t_SL g793 ( .A1(n_433), .A2(n_714), .B1(n_794), .B2(n_795), .C(n_796), .Y(n_793) );
INVx1_ASAP7_75t_L g490 ( .A(n_436), .Y(n_490) );
XOR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_463), .Y(n_436) );
XOR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_462), .Y(n_437) );
NAND4xp75_ASAP7_75t_SL g438 ( .A(n_439), .B(n_452), .C(n_457), .D(n_459), .Y(n_438) );
NOR2xp67_ASAP7_75t_SL g439 ( .A(n_440), .B(n_447), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_443), .C(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g510 ( .A(n_444), .Y(n_510) );
BUFx4f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g468 ( .A(n_445), .Y(n_468) );
BUFx2_ASAP7_75t_L g591 ( .A(n_445), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B(n_450), .Y(n_447) );
OAI21xp5_ASAP7_75t_SL g472 ( .A1(n_449), .A2(n_473), .B(n_474), .Y(n_472) );
OAI21xp5_ASAP7_75t_SL g684 ( .A1(n_449), .A2(n_685), .B(n_686), .Y(n_684) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
INVx1_ASAP7_75t_L g612 ( .A(n_458), .Y(n_612) );
XOR2x2_ASAP7_75t_SL g463 ( .A(n_464), .B(n_488), .Y(n_463) );
NAND2x1p5_ASAP7_75t_L g464 ( .A(n_465), .B(n_477), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_472), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .C(n_470), .Y(n_466) );
INVx2_ASAP7_75t_L g549 ( .A(n_475), .Y(n_549) );
BUFx4f_ASAP7_75t_SL g595 ( .A(n_475), .Y(n_595) );
NOR2x1_ASAP7_75t_L g477 ( .A(n_478), .B(n_483), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_482), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .Y(n_483) );
INVx1_ASAP7_75t_L g614 ( .A(n_485), .Y(n_614) );
INVx1_ASAP7_75t_SL g661 ( .A(n_491), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_572), .B1(n_573), .B2(n_659), .Y(n_491) );
INVx1_ASAP7_75t_L g659 ( .A(n_492), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_531), .B1(n_570), .B2(n_571), .Y(n_492) );
INVx1_ASAP7_75t_L g571 ( .A(n_493), .Y(n_571) );
NAND3x1_ASAP7_75t_L g494 ( .A(n_495), .B(n_511), .C(n_518), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_503), .Y(n_495) );
OAI222xp33_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_499), .B2(n_500), .C1(n_501), .C2(n_502), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_508), .Y(n_629) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_514), .Y(n_511) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g617 ( .A(n_519), .Y(n_617) );
OAI22xp5_ASAP7_75t_SL g520 ( .A1(n_521), .A2(n_523), .B1(n_524), .B2(n_527), .Y(n_520) );
BUFx2_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g652 ( .A(n_526), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g570 ( .A(n_531), .Y(n_570) );
XNOR2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_550), .Y(n_533) );
OAI211xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_537), .B(n_539), .C(n_540), .Y(n_535) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_545), .B1(n_546), .B2(n_547), .Y(n_543) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NOR3xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_557), .C(n_562), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx4_ASAP7_75t_L g604 ( .A(n_554), .Y(n_604) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B1(n_566), .B2(n_567), .Y(n_562) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_567), .A2(n_616), .B1(n_617), .B2(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g799 ( .A(n_568), .Y(n_799) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AO22x1_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B1(n_597), .B2(n_658), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_SL g596 ( .A(n_577), .Y(n_596) );
NAND4xp75_ASAP7_75t_L g577 ( .A(n_578), .B(n_585), .C(n_589), .D(n_593), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_584), .Y(n_609) );
INVx2_ASAP7_75t_L g721 ( .A(n_584), .Y(n_721) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
AND2x2_ASAP7_75t_SL g589 ( .A(n_590), .B(n_592), .Y(n_589) );
INVx1_ASAP7_75t_L g729 ( .A(n_594), .Y(n_729) );
INVx1_ASAP7_75t_L g658 ( .A(n_597), .Y(n_658) );
XNOR2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_632), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_SL g600 ( .A(n_601), .B(n_619), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_610), .C(n_615), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_608), .Y(n_602) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_626), .Y(n_619) );
INVx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .C(n_630), .Y(n_626) );
INVx1_ASAP7_75t_SL g656 ( .A(n_633), .Y(n_656) );
AND2x2_ASAP7_75t_SL g633 ( .A(n_634), .B(n_647), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_639), .C(n_643), .Y(n_634) );
AND4x1_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .C(n_653), .D(n_655), .Y(n_647) );
INVx1_ASAP7_75t_L g707 ( .A(n_649), .Y(n_707) );
BUFx2_ASAP7_75t_L g715 ( .A(n_654), .Y(n_715) );
CKINVDCx16_ASAP7_75t_R g740 ( .A(n_662), .Y(n_740) );
AOI22xp5_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_701), .B1(n_737), .B2(n_738), .Y(n_662) );
INVx1_ASAP7_75t_L g737 ( .A(n_663), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_681), .B1(n_699), .B2(n_700), .Y(n_663) );
INVx2_ASAP7_75t_SL g699 ( .A(n_664), .Y(n_699) );
XOR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_680), .Y(n_664) );
NAND4xp75_ASAP7_75t_L g665 ( .A(n_666), .B(n_669), .C(n_673), .D(n_677), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx2_ASAP7_75t_SL g764 ( .A(n_678), .Y(n_764) );
INVx4_ASAP7_75t_SL g700 ( .A(n_681), .Y(n_700) );
XOR2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_698), .Y(n_681) );
NAND3x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_692), .C(n_695), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_687), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .C(n_691), .Y(n_687) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g738 ( .A(n_701), .Y(n_738) );
INVx1_ASAP7_75t_L g736 ( .A(n_702), .Y(n_736) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_722), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_713), .Y(n_703) );
OAI221xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_706), .B1(n_707), .B2(n_708), .C(n_709), .Y(n_704) );
OAI221xp5_ASAP7_75t_SL g797 ( .A1(n_707), .A2(n_798), .B1(n_799), .B2(n_800), .C(n_801), .Y(n_797) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OAI221xp5_ASAP7_75t_SL g713 ( .A1(n_714), .A2(n_716), .B1(n_717), .B2(n_718), .C(n_719), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx3_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_SL g722 ( .A(n_723), .B(n_728), .Y(n_722) );
OAI222xp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_730), .B1(n_731), .B2(n_732), .C1(n_733), .C2(n_734), .Y(n_728) );
OAI221xp5_ASAP7_75t_L g807 ( .A1(n_729), .A2(n_731), .B1(n_808), .B2(n_809), .C(n_810), .Y(n_807) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
NOR2x1_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .Y(n_742) );
OR2x2_ASAP7_75t_SL g818 ( .A(n_743), .B(n_748), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_745), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_745), .B(n_782), .Y(n_786) );
CKINVDCx16_ASAP7_75t_R g782 ( .A(n_746), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
OAI322xp33_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_780), .A3(n_781), .B1(n_783), .B2(n_787), .C1(n_788), .C2(n_816), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_756), .Y(n_779) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_769), .Y(n_757) );
NOR3xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_762), .C(n_766), .Y(n_758) );
OAI21xp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B(n_765), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_773), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_777), .Y(n_773) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g815 ( .A(n_791), .Y(n_815) );
AND2x2_ASAP7_75t_SL g791 ( .A(n_792), .B(n_803), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_797), .Y(n_792) );
NOR3xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_807), .C(n_812), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
endmodule