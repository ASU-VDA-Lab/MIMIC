module fake_jpeg_8382_n_69 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_69);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_23),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_6),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_27),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_8),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_9),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_14),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_60),
.Y(n_62)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_61),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_54),
.C(n_52),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_55),
.Y(n_65)
);

AOI31xp33_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_53),
.A3(n_58),
.B(n_59),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_46),
.A3(n_19),
.B1(n_20),
.B2(n_22),
.C1(n_24),
.C2(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_18),
.Y(n_69)
);


endmodule