module real_aes_6373_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_150;
wire n_147;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g546 ( .A1(n_0), .A2(n_151), .B(n_547), .C(n_550), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_1), .B(n_491), .Y(n_551) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_2), .B(n_89), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g436 ( .A(n_2), .Y(n_436) );
INVx1_ASAP7_75t_L g185 ( .A(n_3), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_4), .B(n_143), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_5), .A2(n_460), .B(n_485), .Y(n_484) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_6), .A2(n_128), .B(n_476), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_7), .A2(n_35), .B1(n_137), .B2(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_8), .B(n_128), .Y(n_154) );
AND2x6_ASAP7_75t_L g152 ( .A(n_9), .B(n_153), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_10), .A2(n_152), .B(n_450), .C(n_452), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_11), .B(n_36), .Y(n_105) );
INVx1_ASAP7_75t_L g133 ( .A(n_12), .Y(n_133) );
INVx1_ASAP7_75t_L g178 ( .A(n_13), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_14), .B(n_141), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_15), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_16), .B(n_143), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_17), .B(n_129), .Y(n_190) );
AO32x2_ASAP7_75t_L g212 ( .A1(n_18), .A2(n_128), .A3(n_158), .B1(n_169), .B2(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_19), .B(n_137), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_20), .B(n_129), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_21), .A2(n_54), .B1(n_137), .B2(n_215), .Y(n_216) );
AOI22xp33_ASAP7_75t_SL g237 ( .A1(n_22), .A2(n_81), .B1(n_137), .B2(n_141), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_23), .B(n_137), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_24), .A2(n_169), .B(n_450), .C(n_511), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_25), .A2(n_169), .B(n_450), .C(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_26), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_27), .B(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_28), .A2(n_460), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_29), .B(n_171), .Y(n_209) );
INVx2_ASAP7_75t_L g139 ( .A(n_30), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_31), .A2(n_462), .B(n_470), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_32), .B(n_137), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_33), .B(n_171), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_34), .B(n_223), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_37), .B(n_509), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_38), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g113 ( .A1(n_39), .A2(n_78), .B1(n_114), .B2(n_115), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_39), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_40), .B(n_143), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_41), .B(n_460), .Y(n_477) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_42), .A2(n_79), .B1(n_431), .B2(n_743), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_42), .Y(n_743) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_43), .A2(n_462), .B(n_464), .C(n_470), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_44), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g548 ( .A(n_45), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_46), .A2(n_103), .B1(n_111), .B2(n_755), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_47), .A2(n_90), .B1(n_215), .B2(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g465 ( .A(n_48), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_49), .B(n_137), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_50), .B(n_137), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_51), .B(n_740), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_51), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_52), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_53), .B(n_149), .Y(n_148) );
AOI22xp33_ASAP7_75t_SL g194 ( .A1(n_55), .A2(n_59), .B1(n_137), .B2(n_141), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_56), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_57), .B(n_137), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_58), .B(n_137), .Y(n_220) );
INVx1_ASAP7_75t_L g153 ( .A(n_60), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_61), .B(n_460), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_62), .B(n_491), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_63), .A2(n_149), .B(n_181), .C(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_64), .B(n_137), .Y(n_186) );
INVx1_ASAP7_75t_L g132 ( .A(n_65), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_66), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_67), .B(n_143), .Y(n_501) );
AO32x2_ASAP7_75t_L g233 ( .A1(n_68), .A2(n_128), .A3(n_169), .B1(n_234), .B2(n_238), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_69), .B(n_144), .Y(n_453) );
INVx1_ASAP7_75t_L g164 ( .A(n_70), .Y(n_164) );
INVx1_ASAP7_75t_L g204 ( .A(n_71), .Y(n_204) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_72), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_73), .B(n_467), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_74), .A2(n_450), .B(n_470), .C(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_75), .B(n_141), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_76), .Y(n_486) );
INVx1_ASAP7_75t_L g110 ( .A(n_77), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_78), .Y(n_114) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_79), .A2(n_120), .B1(n_430), .B2(n_431), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_79), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_80), .B(n_466), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_82), .B(n_215), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_83), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_84), .B(n_141), .Y(n_208) );
INVx2_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_86), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_87), .B(n_168), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_88), .B(n_141), .Y(n_140) );
OR2x2_ASAP7_75t_L g434 ( .A(n_89), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g724 ( .A(n_89), .Y(n_724) );
OR2x2_ASAP7_75t_L g748 ( .A(n_89), .B(n_734), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_91), .A2(n_101), .B1(n_141), .B2(n_142), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_92), .B(n_460), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_93), .Y(n_731) );
INVx1_ASAP7_75t_L g500 ( .A(n_94), .Y(n_500) );
INVxp67_ASAP7_75t_L g489 ( .A(n_95), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_96), .B(n_141), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_97), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g446 ( .A(n_98), .Y(n_446) );
INVx1_ASAP7_75t_L g524 ( .A(n_99), .Y(n_524) );
AND2x2_ASAP7_75t_L g472 ( .A(n_100), .B(n_171), .Y(n_472) );
BUFx4f_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx12_ASAP7_75t_R g757 ( .A(n_104), .Y(n_757) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g435 ( .A(n_105), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO221x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_735), .B1(n_738), .B2(n_749), .C(n_751), .Y(n_111) );
OAI222xp33_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_116), .B1(n_725), .B2(n_726), .C1(n_731), .C2(n_732), .Y(n_112) );
INVx1_ASAP7_75t_L g725 ( .A(n_113), .Y(n_725) );
INVxp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI22xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_432), .B1(n_437), .B2(n_721), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_119), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_727) );
INVx2_ASAP7_75t_L g430 ( .A(n_120), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_120), .A2(n_430), .B1(n_741), .B2(n_742), .Y(n_740) );
NAND2x1p5_ASAP7_75t_L g120 ( .A(n_121), .B(n_354), .Y(n_120) );
AND2x2_ASAP7_75t_SL g121 ( .A(n_122), .B(n_312), .Y(n_121) );
NOR4xp25_ASAP7_75t_L g122 ( .A(n_123), .B(n_252), .C(n_288), .D(n_302), .Y(n_122) );
OAI221xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_196), .B1(n_228), .B2(n_239), .C(n_243), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_124), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_172), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_155), .Y(n_126) );
AND2x2_ASAP7_75t_L g249 ( .A(n_127), .B(n_156), .Y(n_249) );
INVx3_ASAP7_75t_L g257 ( .A(n_127), .Y(n_257) );
AND2x2_ASAP7_75t_L g311 ( .A(n_127), .B(n_175), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_127), .B(n_174), .Y(n_347) );
AND2x2_ASAP7_75t_L g405 ( .A(n_127), .B(n_267), .Y(n_405) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_134), .B(n_154), .Y(n_127) );
INVx4_ASAP7_75t_L g195 ( .A(n_128), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_128), .A2(n_477), .B(n_478), .Y(n_476) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_128), .Y(n_483) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g158 ( .A(n_129), .Y(n_158) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_130), .B(n_131), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
OAI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_146), .B(n_152), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_140), .B(n_143), .Y(n_135) );
INVx3_ASAP7_75t_L g203 ( .A(n_137), .Y(n_203) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_137), .Y(n_526) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g215 ( .A(n_138), .Y(n_215) );
BUFx3_ASAP7_75t_L g236 ( .A(n_138), .Y(n_236) );
AND2x6_ASAP7_75t_L g450 ( .A(n_138), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g142 ( .A(n_139), .Y(n_142) );
INVx1_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
INVx2_ASAP7_75t_L g179 ( .A(n_141), .Y(n_179) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_143), .A2(n_161), .B(n_162), .Y(n_160) );
O2A1O1Ixp5_ASAP7_75t_SL g202 ( .A1(n_143), .A2(n_203), .B(n_204), .C(n_205), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_143), .B(n_489), .Y(n_488) );
INVx5_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OAI22xp5_ASAP7_75t_SL g234 ( .A1(n_144), .A2(n_168), .B1(n_235), .B2(n_237), .Y(n_234) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_145), .Y(n_168) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_145), .Y(n_183) );
INVx1_ASAP7_75t_L g223 ( .A(n_145), .Y(n_223) );
AND2x2_ASAP7_75t_L g448 ( .A(n_145), .B(n_150), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_145), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_151), .Y(n_146) );
INVx2_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_151), .A2(n_165), .B(n_185), .C(n_186), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_151), .A2(n_168), .B1(n_193), .B2(n_194), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_151), .A2(n_168), .B1(n_214), .B2(n_216), .Y(n_213) );
BUFx3_ASAP7_75t_L g169 ( .A(n_152), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g176 ( .A1(n_152), .A2(n_177), .B(n_184), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_152), .A2(n_202), .B(n_206), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_152), .A2(n_219), .B(n_224), .Y(n_218) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_152), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g460 ( .A(n_152), .B(n_448), .Y(n_460) );
INVx4_ASAP7_75t_SL g471 ( .A(n_152), .Y(n_471) );
AND2x2_ASAP7_75t_L g240 ( .A(n_155), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g254 ( .A(n_155), .B(n_175), .Y(n_254) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_156), .B(n_175), .Y(n_269) );
AND2x2_ASAP7_75t_L g281 ( .A(n_156), .B(n_257), .Y(n_281) );
OR2x2_ASAP7_75t_L g283 ( .A(n_156), .B(n_241), .Y(n_283) );
AND2x2_ASAP7_75t_L g318 ( .A(n_156), .B(n_241), .Y(n_318) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_156), .Y(n_363) );
INVx1_ASAP7_75t_L g371 ( .A(n_156), .Y(n_371) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_170), .Y(n_156) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_157), .A2(n_176), .B(n_187), .Y(n_175) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_158), .B(n_456), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_163), .B(n_169), .Y(n_159) );
O2A1O1Ixp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_166), .C(n_167), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_165), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_167), .A2(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx4_ASAP7_75t_L g549 ( .A(n_168), .Y(n_549) );
NAND3xp33_ASAP7_75t_L g191 ( .A(n_169), .B(n_192), .C(n_195), .Y(n_191) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_171), .A2(n_201), .B(n_209), .Y(n_200) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_171), .A2(n_218), .B(n_227), .Y(n_217) );
INVx2_ASAP7_75t_L g238 ( .A(n_171), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_171), .A2(n_459), .B(n_461), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_171), .A2(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g517 ( .A(n_171), .Y(n_517) );
OAI221xp5_ASAP7_75t_L g288 ( .A1(n_172), .A2(n_289), .B1(n_293), .B2(n_297), .C(n_298), .Y(n_288) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g248 ( .A(n_173), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_188), .Y(n_173) );
INVx2_ASAP7_75t_L g247 ( .A(n_174), .Y(n_247) );
AND2x2_ASAP7_75t_L g300 ( .A(n_174), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g319 ( .A(n_174), .B(n_257), .Y(n_319) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g382 ( .A(n_175), .B(n_257), .Y(n_382) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_180), .C(n_181), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_179), .A2(n_453), .B(n_454), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_179), .A2(n_480), .B(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_181), .A2(n_524), .B(n_525), .C(n_526), .Y(n_523) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_182), .A2(n_207), .B(n_208), .Y(n_206) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g467 ( .A(n_183), .Y(n_467) );
AND2x2_ASAP7_75t_L g304 ( .A(n_188), .B(n_249), .Y(n_304) );
OAI322xp33_ASAP7_75t_L g372 ( .A1(n_188), .A2(n_328), .A3(n_373), .B1(n_375), .B2(n_378), .C1(n_380), .C2(n_384), .Y(n_372) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2x1_ASAP7_75t_L g255 ( .A(n_189), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g268 ( .A(n_189), .Y(n_268) );
AND2x2_ASAP7_75t_L g377 ( .A(n_189), .B(n_257), .Y(n_377) );
AND2x2_ASAP7_75t_L g409 ( .A(n_189), .B(n_281), .Y(n_409) );
OR2x2_ASAP7_75t_L g412 ( .A(n_189), .B(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
INVx1_ASAP7_75t_L g242 ( .A(n_190), .Y(n_242) );
AO21x1_ASAP7_75t_L g241 ( .A1(n_192), .A2(n_195), .B(n_242), .Y(n_241) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_195), .A2(n_445), .B(n_455), .Y(n_444) );
INVx3_ASAP7_75t_L g491 ( .A(n_195), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_195), .B(n_503), .Y(n_502) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_195), .A2(n_521), .B(n_528), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_195), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_210), .Y(n_197) );
INVx1_ASAP7_75t_L g425 ( .A(n_198), .Y(n_425) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
OR2x2_ASAP7_75t_L g230 ( .A(n_199), .B(n_217), .Y(n_230) );
INVx2_ASAP7_75t_L g265 ( .A(n_199), .Y(n_265) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g287 ( .A(n_200), .Y(n_287) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_200), .Y(n_295) );
OR2x2_ASAP7_75t_L g419 ( .A(n_200), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g244 ( .A(n_210), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g284 ( .A(n_210), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g336 ( .A(n_210), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_217), .Y(n_210) );
AND2x2_ASAP7_75t_L g231 ( .A(n_211), .B(n_232), .Y(n_231) );
NOR2xp67_ASAP7_75t_L g291 ( .A(n_211), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g345 ( .A(n_211), .B(n_233), .Y(n_345) );
OR2x2_ASAP7_75t_L g353 ( .A(n_211), .B(n_287), .Y(n_353) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
BUFx2_ASAP7_75t_L g262 ( .A(n_212), .Y(n_262) );
AND2x2_ASAP7_75t_L g272 ( .A(n_212), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g296 ( .A(n_212), .B(n_217), .Y(n_296) );
AND2x2_ASAP7_75t_L g360 ( .A(n_212), .B(n_233), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_217), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_217), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g273 ( .A(n_217), .Y(n_273) );
INVx1_ASAP7_75t_L g278 ( .A(n_217), .Y(n_278) );
AND2x2_ASAP7_75t_L g290 ( .A(n_217), .B(n_291), .Y(n_290) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_217), .Y(n_368) );
INVx1_ASAP7_75t_L g420 ( .A(n_217), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_222), .Y(n_219) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
AND2x2_ASAP7_75t_L g397 ( .A(n_229), .B(n_306), .Y(n_397) );
INVx2_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g324 ( .A(n_231), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g423 ( .A(n_231), .B(n_358), .Y(n_423) );
INVx1_ASAP7_75t_L g245 ( .A(n_232), .Y(n_245) );
AND2x2_ASAP7_75t_L g271 ( .A(n_232), .B(n_265), .Y(n_271) );
BUFx2_ASAP7_75t_L g330 ( .A(n_232), .Y(n_330) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_233), .Y(n_251) );
INVx1_ASAP7_75t_L g261 ( .A(n_233), .Y(n_261) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_236), .Y(n_469) );
INVx2_ASAP7_75t_L g550 ( .A(n_236), .Y(n_550) );
INVx1_ASAP7_75t_L g514 ( .A(n_238), .Y(n_514) );
NOR2xp67_ASAP7_75t_L g399 ( .A(n_239), .B(n_246), .Y(n_399) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AOI32xp33_ASAP7_75t_L g243 ( .A1(n_240), .A2(n_244), .A3(n_246), .B1(n_248), .B2(n_250), .Y(n_243) );
AND2x2_ASAP7_75t_L g383 ( .A(n_240), .B(n_256), .Y(n_383) );
AND2x2_ASAP7_75t_L g421 ( .A(n_240), .B(n_319), .Y(n_421) );
INVx1_ASAP7_75t_L g301 ( .A(n_241), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_245), .B(n_307), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_246), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_246), .B(n_249), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_246), .B(n_318), .Y(n_400) );
OR2x2_ASAP7_75t_L g414 ( .A(n_246), .B(n_283), .Y(n_414) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g341 ( .A(n_247), .B(n_249), .Y(n_341) );
OR2x2_ASAP7_75t_L g350 ( .A(n_247), .B(n_337), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_249), .B(n_300), .Y(n_322) );
INVx2_ASAP7_75t_L g337 ( .A(n_251), .Y(n_337) );
OR2x2_ASAP7_75t_L g352 ( .A(n_251), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g367 ( .A(n_251), .B(n_368), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g424 ( .A1(n_251), .A2(n_344), .B(n_425), .C(n_426), .Y(n_424) );
OAI321xp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_258), .A3(n_263), .B1(n_266), .B2(n_270), .C(n_274), .Y(n_252) );
INVx1_ASAP7_75t_L g365 ( .A(n_253), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g376 ( .A(n_254), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g328 ( .A(n_256), .Y(n_328) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_257), .B(n_371), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g395 ( .A1(n_258), .A2(n_396), .B1(n_398), .B2(n_400), .C(n_401), .Y(n_395) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
AND2x2_ASAP7_75t_L g333 ( .A(n_260), .B(n_307), .Y(n_333) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_261), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_262), .Y(n_306) );
A2O1A1Ixp33_ASAP7_75t_L g348 ( .A1(n_263), .A2(n_304), .B(n_349), .C(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g315 ( .A(n_265), .B(n_272), .Y(n_315) );
BUFx2_ASAP7_75t_L g325 ( .A(n_265), .Y(n_325) );
INVx1_ASAP7_75t_L g340 ( .A(n_265), .Y(n_340) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
OR2x2_ASAP7_75t_L g346 ( .A(n_268), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g429 ( .A(n_268), .Y(n_429) );
INVx1_ASAP7_75t_L g422 ( .A(n_269), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
AND2x2_ASAP7_75t_L g275 ( .A(n_271), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g379 ( .A(n_271), .B(n_296), .Y(n_379) );
INVx1_ASAP7_75t_L g308 ( .A(n_272), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_279), .B1(n_282), .B2(n_284), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_276), .B(n_392), .Y(n_391) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g344 ( .A(n_277), .B(n_345), .Y(n_344) );
BUFx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_SL g307 ( .A(n_278), .B(n_287), .Y(n_307) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g299 ( .A(n_281), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g309 ( .A(n_283), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
OAI221xp5_ASAP7_75t_L g403 ( .A1(n_286), .A2(n_404), .B1(n_406), .B2(n_407), .C(n_408), .Y(n_403) );
INVx1_ASAP7_75t_L g292 ( .A(n_287), .Y(n_292) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_287), .Y(n_358) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_290), .B(n_409), .Y(n_408) );
OAI21xp5_ASAP7_75t_L g298 ( .A1(n_291), .A2(n_296), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_294), .B(n_304), .Y(n_401) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g370 ( .A(n_295), .Y(n_370) );
AND2x2_ASAP7_75t_L g329 ( .A(n_296), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g418 ( .A(n_296), .Y(n_418) );
INVx1_ASAP7_75t_L g334 ( .A(n_299), .Y(n_334) );
INVx1_ASAP7_75t_L g389 ( .A(n_300), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_305), .B1(n_308), .B2(n_309), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_306), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g374 ( .A(n_307), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_307), .B(n_345), .Y(n_411) );
OR2x2_ASAP7_75t_L g384 ( .A(n_308), .B(n_337), .Y(n_384) );
INVx1_ASAP7_75t_L g323 ( .A(n_309), .Y(n_323) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_311), .B(n_362), .Y(n_361) );
NOR3xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_331), .C(n_342), .Y(n_312) );
OAI211xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B(n_320), .C(n_326), .Y(n_313) );
INVxp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_315), .A2(n_386), .B1(n_390), .B2(n_393), .C(n_395), .Y(n_385) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x2_ASAP7_75t_L g327 ( .A(n_318), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g381 ( .A(n_318), .B(n_382), .Y(n_381) );
OAI211xp5_ASAP7_75t_L g366 ( .A1(n_319), .A2(n_367), .B(n_369), .C(n_371), .Y(n_366) );
INVx2_ASAP7_75t_L g413 ( .A(n_319), .Y(n_413) );
OAI21xp5_ASAP7_75t_SL g320 ( .A1(n_321), .A2(n_323), .B(n_324), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g392 ( .A(n_325), .B(n_345), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
OAI21xp5_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_334), .B(n_335), .Y(n_331) );
INVxp67_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI21xp5_ASAP7_75t_SL g335 ( .A1(n_336), .A2(n_338), .B(n_341), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_336), .B(n_365), .Y(n_364) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_341), .B(n_428), .Y(n_427) );
OAI21xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_346), .B(n_348), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g369 ( .A(n_345), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND4x1_ASAP7_75t_L g354 ( .A(n_355), .B(n_385), .C(n_402), .D(n_424), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_372), .Y(n_355) );
OAI211xp5_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_361), .B(n_364), .C(n_366), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_360), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_371), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g406 ( .A(n_381), .Y(n_406) );
INVx2_ASAP7_75t_SL g394 ( .A(n_382), .Y(n_394) );
OR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g407 ( .A(n_392), .Y(n_407) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NOR2xp33_ASAP7_75t_SL g402 ( .A(n_403), .B(n_410), .Y(n_402) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
OAI221xp5_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_412), .B1(n_414), .B2(n_415), .C(n_416), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g728 ( .A(n_433), .Y(n_728) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g723 ( .A(n_435), .B(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g734 ( .A(n_435), .Y(n_734) );
INVx2_ASAP7_75t_L g729 ( .A(n_437), .Y(n_729) );
OR3x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_619), .C(n_684), .Y(n_437) );
NAND4xp25_ASAP7_75t_SL g438 ( .A(n_439), .B(n_560), .C(n_586), .D(n_609), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_492), .B1(n_530), .B2(n_537), .C(n_552), .Y(n_439) );
CKINVDCx14_ASAP7_75t_R g440 ( .A(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_441), .A2(n_553), .B1(n_577), .B2(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_473), .Y(n_441) );
INVx1_ASAP7_75t_SL g613 ( .A(n_442), .Y(n_613) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_457), .Y(n_442) );
OR2x2_ASAP7_75t_L g535 ( .A(n_443), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g555 ( .A(n_443), .B(n_474), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_443), .B(n_482), .Y(n_568) );
AND2x2_ASAP7_75t_L g585 ( .A(n_443), .B(n_457), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_443), .B(n_533), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_443), .B(n_584), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_443), .B(n_473), .Y(n_706) );
AOI211xp5_ASAP7_75t_SL g717 ( .A1(n_443), .A2(n_623), .B(n_718), .C(n_719), .Y(n_717) );
INVx5_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_444), .B(n_474), .Y(n_589) );
AND2x2_ASAP7_75t_L g592 ( .A(n_444), .B(n_475), .Y(n_592) );
OR2x2_ASAP7_75t_L g637 ( .A(n_444), .B(n_474), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_444), .B(n_482), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B(n_449), .Y(n_445) );
INVx5_ASAP7_75t_L g463 ( .A(n_450), .Y(n_463) );
INVx5_ASAP7_75t_SL g536 ( .A(n_457), .Y(n_536) );
AND2x2_ASAP7_75t_L g554 ( .A(n_457), .B(n_555), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_457), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g640 ( .A(n_457), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g672 ( .A(n_457), .B(n_482), .Y(n_672) );
OR2x2_ASAP7_75t_L g678 ( .A(n_457), .B(n_568), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_457), .B(n_628), .Y(n_687) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_472), .Y(n_457) );
BUFx2_ASAP7_75t_L g509 ( .A(n_460), .Y(n_509) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_463), .A2(n_471), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_SL g544 ( .A1(n_463), .A2(n_471), .B(n_545), .C(n_546), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B(n_468), .C(n_469), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_466), .A2(n_469), .B(n_500), .C(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_482), .Y(n_473) );
AND2x2_ASAP7_75t_L g569 ( .A(n_474), .B(n_536), .Y(n_569) );
INVx1_ASAP7_75t_SL g582 ( .A(n_474), .Y(n_582) );
OR2x2_ASAP7_75t_L g617 ( .A(n_474), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g623 ( .A(n_474), .B(n_482), .Y(n_623) );
AND2x2_ASAP7_75t_L g681 ( .A(n_474), .B(n_533), .Y(n_681) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_475), .B(n_536), .Y(n_608) );
INVx3_ASAP7_75t_L g533 ( .A(n_482), .Y(n_533) );
OR2x2_ASAP7_75t_L g574 ( .A(n_482), .B(n_536), .Y(n_574) );
AND2x2_ASAP7_75t_L g584 ( .A(n_482), .B(n_582), .Y(n_584) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_482), .Y(n_632) );
AND2x2_ASAP7_75t_L g641 ( .A(n_482), .B(n_555), .Y(n_641) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_490), .Y(n_482) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_491), .A2(n_543), .B(n_551), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_492), .A2(n_658), .B1(n_660), .B2(n_662), .C(n_665), .Y(n_657) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_504), .Y(n_493) );
AND2x2_ASAP7_75t_L g631 ( .A(n_494), .B(n_612), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_494), .B(n_690), .Y(n_694) );
OR2x2_ASAP7_75t_L g715 ( .A(n_494), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_494), .B(n_720), .Y(n_719) );
BUFx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx5_ASAP7_75t_L g562 ( .A(n_495), .Y(n_562) );
AND2x2_ASAP7_75t_L g639 ( .A(n_495), .B(n_506), .Y(n_639) );
AND2x2_ASAP7_75t_L g700 ( .A(n_495), .B(n_579), .Y(n_700) );
AND2x2_ASAP7_75t_L g713 ( .A(n_495), .B(n_533), .Y(n_713) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_518), .Y(n_504) );
AND2x4_ASAP7_75t_L g540 ( .A(n_505), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g558 ( .A(n_505), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g565 ( .A(n_505), .Y(n_565) );
AND2x2_ASAP7_75t_L g634 ( .A(n_505), .B(n_612), .Y(n_634) );
AND2x2_ASAP7_75t_L g644 ( .A(n_505), .B(n_562), .Y(n_644) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_505), .Y(n_652) );
AND2x2_ASAP7_75t_L g664 ( .A(n_505), .B(n_542), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_505), .B(n_596), .Y(n_668) );
AND2x2_ASAP7_75t_L g705 ( .A(n_505), .B(n_700), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_505), .B(n_579), .Y(n_716) );
OR2x2_ASAP7_75t_L g718 ( .A(n_505), .B(n_654), .Y(n_718) );
INVx5_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g604 ( .A(n_506), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g614 ( .A(n_506), .B(n_559), .Y(n_614) );
AND2x2_ASAP7_75t_L g626 ( .A(n_506), .B(n_542), .Y(n_626) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_506), .Y(n_656) );
AND2x4_ASAP7_75t_L g690 ( .A(n_506), .B(n_541), .Y(n_690) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_515), .Y(n_506) );
AOI21xp5_ASAP7_75t_SL g507 ( .A1(n_508), .A2(n_510), .B(n_514), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
BUFx2_ASAP7_75t_L g539 ( .A(n_518), .Y(n_539) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g579 ( .A(n_519), .Y(n_579) );
AND2x2_ASAP7_75t_L g612 ( .A(n_519), .B(n_542), .Y(n_612) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g559 ( .A(n_520), .B(n_542), .Y(n_559) );
BUFx2_ASAP7_75t_L g605 ( .A(n_520), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_532), .B(n_613), .Y(n_692) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_533), .B(n_555), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_533), .B(n_536), .Y(n_594) );
AND2x2_ASAP7_75t_L g649 ( .A(n_533), .B(n_585), .Y(n_649) );
AOI221xp5_ASAP7_75t_SL g586 ( .A1(n_534), .A2(n_587), .B1(n_595), .B2(n_597), .C(n_601), .Y(n_586) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g581 ( .A(n_535), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g622 ( .A(n_535), .B(n_623), .Y(n_622) );
OAI321xp33_ASAP7_75t_L g629 ( .A1(n_535), .A2(n_588), .A3(n_630), .B1(n_632), .B2(n_633), .C(n_635), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_536), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_539), .B(n_690), .Y(n_708) );
AND2x2_ASAP7_75t_L g595 ( .A(n_540), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_540), .B(n_599), .Y(n_598) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_541), .Y(n_571) );
AND2x2_ASAP7_75t_L g578 ( .A(n_541), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_541), .B(n_653), .Y(n_683) );
INVx1_ASAP7_75t_L g720 ( .A(n_541), .Y(n_720) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_556), .B(n_557), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_554), .A2(n_664), .B(n_713), .C(n_714), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_555), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_555), .B(n_593), .Y(n_659) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g602 ( .A(n_559), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_559), .B(n_562), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_559), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_559), .B(n_644), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_563), .B1(n_575), .B2(n_580), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g576 ( .A(n_562), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g599 ( .A(n_562), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g611 ( .A(n_562), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_562), .B(n_605), .Y(n_647) );
OR2x2_ASAP7_75t_L g654 ( .A(n_562), .B(n_579), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_562), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g704 ( .A(n_562), .B(n_690), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .B1(n_570), .B2(n_572), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g610 ( .A(n_565), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_568), .A2(n_583), .B1(n_651), .B2(n_655), .Y(n_650) );
INVx1_ASAP7_75t_L g698 ( .A(n_569), .Y(n_698) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_573), .A2(n_610), .B1(n_613), .B2(n_614), .C(n_615), .Y(n_609) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g588 ( .A(n_574), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_578), .B(n_644), .Y(n_676) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_579), .Y(n_596) );
INVx1_ASAP7_75t_L g600 ( .A(n_579), .Y(n_600) );
NAND2xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g618 ( .A(n_585), .Y(n_618) );
AND2x2_ASAP7_75t_L g627 ( .A(n_585), .B(n_628), .Y(n_627) );
NAND2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx2_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g671 ( .A(n_592), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_595), .A2(n_621), .B1(n_624), .B2(n_627), .C(n_629), .Y(n_620) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_599), .B(n_656), .Y(n_655) );
AOI21xp33_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_603), .B(n_606), .Y(n_601) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
CKINVDCx16_ASAP7_75t_R g703 ( .A(n_606), .Y(n_703) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
OR2x2_ASAP7_75t_L g645 ( .A(n_608), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g666 ( .A(n_611), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_611), .B(n_671), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_614), .B(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
NAND4xp25_ASAP7_75t_L g619 ( .A(n_620), .B(n_638), .C(n_657), .D(n_670), .Y(n_619) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g628 ( .A(n_623), .Y(n_628) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g661 ( .A(n_632), .B(n_637), .Y(n_661) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI211xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B(n_642), .C(n_650), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_640), .A2(n_682), .B(n_710), .C(n_717), .Y(n_709) );
INVx1_ASAP7_75t_SL g669 ( .A(n_641), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B1(n_647), .B2(n_648), .Y(n_642) );
INVx1_ASAP7_75t_L g673 ( .A(n_647), .Y(n_673) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_653), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_653), .B(n_664), .Y(n_697) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g674 ( .A(n_664), .Y(n_674) );
AOI21xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B(n_669), .Y(n_665) );
INVxp33_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI322xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_673), .A3(n_674), .B1(n_675), .B2(n_677), .C1(n_679), .C2(n_682), .Y(n_670) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND3xp33_ASAP7_75t_SL g684 ( .A(n_685), .B(n_702), .C(n_709), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B1(n_691), .B2(n_693), .C(n_695), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g701 ( .A(n_690), .Y(n_701) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_705), .B2(n_706), .C(n_707), .Y(n_702) );
NAND2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVxp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g730 ( .A(n_722), .Y(n_730) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_724), .B(n_734), .Y(n_733) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_SL g750 ( .A(n_736), .Y(n_750) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NOR3xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_744), .C(n_747), .Y(n_738) );
INVx1_ASAP7_75t_L g746 ( .A(n_740), .Y(n_746) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g754 ( .A(n_748), .Y(n_754) );
BUFx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
endmodule