module fake_jpeg_26452_n_273 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_49),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_16),
.B1(n_31),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_17),
.B1(n_24),
.B2(n_32),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_56),
.Y(n_65)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_16),
.Y(n_56)
);

INVx5_ASAP7_75t_SL g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_40),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_68),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_21),
.B1(n_31),
.B2(n_38),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_39),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_37),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_33),
.B1(n_39),
.B2(n_35),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_63),
.A2(n_73),
.B1(n_82),
.B2(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_70),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_40),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_37),
.B(n_32),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_47),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_17),
.B(n_19),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_36),
.B1(n_35),
.B2(n_40),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_43),
.A2(n_36),
.B1(n_35),
.B2(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_51),
.B1(n_53),
.B2(n_44),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_87),
.A2(n_90),
.B1(n_83),
.B2(n_20),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_40),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_93),
.B(n_101),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_53),
.B1(n_44),
.B2(n_45),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_88),
.C(n_97),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_37),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_59),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_95),
.B(n_104),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_103),
.B1(n_67),
.B2(n_80),
.Y(n_118)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_37),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_37),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_30),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_30),
.Y(n_119)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_110),
.B(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_122),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_106),
.A2(n_82),
.B1(n_68),
.B2(n_73),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_113),
.A2(n_116),
.B1(n_131),
.B2(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_69),
.B1(n_79),
.B2(n_81),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_135),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_135),
.B1(n_115),
.B2(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_120),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_67),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_92),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_27),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_69),
.B1(n_74),
.B2(n_66),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_123),
.A2(n_89),
.B1(n_105),
.B2(n_96),
.Y(n_144)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_126),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_66),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_24),
.B(n_20),
.Y(n_129)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_132),
.B(n_122),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_86),
.B(n_19),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_132),
.B(n_133),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_98),
.B(n_29),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_85),
.A2(n_83),
.B1(n_23),
.B2(n_22),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

HAxp5_ASAP7_75t_SL g148 ( 
.A(n_136),
.B(n_116),
.CON(n_148),
.SN(n_148)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_137),
.B(n_11),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_98),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_151),
.Y(n_180)
);

AOI22x1_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_93),
.B1(n_89),
.B2(n_96),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_142),
.A2(n_10),
.B1(n_14),
.B2(n_4),
.Y(n_177)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_143),
.B(n_146),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_144),
.A2(n_149),
.B1(n_2),
.B2(n_5),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_93),
.C(n_105),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_120),
.C(n_114),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g183 ( 
.A(n_148),
.B(n_1),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_104),
.B(n_94),
.C(n_91),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_0),
.B(n_1),
.Y(n_175)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_129),
.B1(n_110),
.B2(n_133),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_158),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g158 ( 
.A(n_126),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_111),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_160),
.B(n_162),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_111),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_142),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_173),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_131),
.B1(n_124),
.B2(n_91),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_111),
.B1(n_23),
.B2(n_22),
.Y(n_172)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_22),
.C(n_29),
.Y(n_173)
);

A2O1A1O1Ixp25_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_140),
.B(n_153),
.C(n_159),
.D(n_164),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_175),
.B(n_176),
.Y(n_195)
);

XNOR2x2_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_9),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_177),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_7),
.C(n_14),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_178),
.B(n_184),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_156),
.B(n_148),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_163),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_145),
.B1(n_161),
.B2(n_141),
.Y(n_199)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_186),
.B(n_167),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_197),
.A2(n_205),
.B(n_210),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_198),
.B(n_150),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_185),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_201),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_179),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_202),
.B(n_207),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_147),
.B1(n_159),
.B2(n_150),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_206),
.B1(n_208),
.B2(n_11),
.Y(n_225)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_180),
.B1(n_182),
.B2(n_174),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_175),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_183),
.B1(n_181),
.B2(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_169),
.C(n_165),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_211),
.B(n_215),
.Y(n_231)
);

NOR3xp33_ASAP7_75t_SL g215 ( 
.A(n_199),
.B(n_157),
.C(n_176),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_188),
.C(n_178),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_217),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_150),
.C(n_170),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_218),
.B(n_225),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_155),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_222),
.Y(n_237)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_208),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_155),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_226),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_11),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_203),
.B1(n_205),
.B2(n_196),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_236),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_216),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_238),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_203),
.B1(n_196),
.B2(n_200),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_226),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_239),
.A2(n_219),
.B1(n_225),
.B2(n_215),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_194),
.B1(n_210),
.B2(n_209),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_244),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_246),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_218),
.C(n_195),
.Y(n_246)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_212),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_233),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_192),
.C(n_5),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_249),
.C(n_233),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_192),
.C(n_5),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_257),
.B(n_13),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_247),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_253),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_248),
.B(n_231),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_249),
.B(n_227),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_255),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_240),
.B(n_250),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_6),
.Y(n_257)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_258),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_262),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_250),
.B(n_241),
.Y(n_262)
);

OAI21x1_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_246),
.B(n_6),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_267),
.B(n_265),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_260),
.B(n_7),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_268),
.A2(n_269),
.B(n_13),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_12),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_15),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_271),
.A2(n_15),
.B(n_2),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_15),
.Y(n_273)
);


endmodule