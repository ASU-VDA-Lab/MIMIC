module fake_jpeg_26870_n_76 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_76);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_76;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_28;
wire n_38;
wire n_44;
wire n_36;
wire n_74;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_75;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;
wire n_70;
wire n_66;

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_14),
.B(n_24),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_13),
.A2(n_11),
.B(n_27),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_0),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_32),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_30),
.B(n_32),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_26),
.C(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_50),
.C(n_52),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_15),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_48),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_12),
.B(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_3),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_18),
.B1(n_23),
.B2(n_22),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_4),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_55),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_21),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_62),
.C(n_46),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_20),
.B1(n_19),
.B2(n_10),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_63),
.B1(n_53),
.B2(n_7),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_4),
.C(n_5),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_68),
.Y(n_70)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_67),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_47),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_57),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.B(n_70),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_71),
.B1(n_58),
.B2(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_61),
.Y(n_76)
);


endmodule