module real_jpeg_32386_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_323;
wire n_176;
wire n_166;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_0),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g377 ( 
.A(n_0),
.Y(n_377)
);

NAND2x1p5_ASAP7_75t_L g62 ( 
.A(n_1),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_1),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_R g285 ( 
.A(n_1),
.B(n_286),
.Y(n_285)
);

NAND2x1_ASAP7_75t_L g291 ( 
.A(n_1),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_1),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_1),
.B(n_386),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_1),
.B(n_155),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_1),
.B(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_1),
.B(n_283),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_41),
.Y(n_40)
);

AND2x4_ASAP7_75t_L g65 ( 
.A(n_2),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_2),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_2),
.B(n_124),
.Y(n_123)
);

NAND2x1p5_ASAP7_75t_L g188 ( 
.A(n_2),
.B(n_107),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_2),
.B(n_247),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_2),
.B(n_469),
.Y(n_468)
);

NAND2x1_ASAP7_75t_L g91 ( 
.A(n_3),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_3),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_3),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_3),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_3),
.B(n_326),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_3),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_3),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_3),
.B(n_419),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_5),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_5),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_5),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_5),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_5),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_5),
.B(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_5),
.B(n_433),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_6),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_6),
.Y(n_177)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_8),
.A2(n_19),
.B(n_22),
.Y(n_18)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_9),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_9),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_9),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_10),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_10),
.B(n_46),
.Y(n_53)
);

NAND2x1_ASAP7_75t_L g69 ( 
.A(n_10),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_10),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_10),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_10),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_10),
.B(n_283),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_10),
.B(n_477),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_10),
.B(n_500),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_11),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_11),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_12),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_38),
.Y(n_37)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_13),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_13),
.B(n_60),
.Y(n_59)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_13),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_13),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_13),
.B(n_35),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_13),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_SL g235 ( 
.A(n_13),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_14),
.B(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_14),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_14),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_14),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_14),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_14),
.B(n_472),
.Y(n_471)
);

NAND2x1_ASAP7_75t_SL g481 ( 
.A(n_14),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_14),
.B(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_15),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_16),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_16),
.Y(n_260)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_16),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_17),
.B(n_76),
.Y(n_75)
);

NAND2x1_ASAP7_75t_L g106 ( 
.A(n_17),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_17),
.B(n_121),
.Y(n_120)
);

AND2x4_ASAP7_75t_SL g175 ( 
.A(n_17),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_17),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_17),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_17),
.B(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_17),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1O1Ixp25_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_235),
.B(n_459),
.C(n_552),
.D(n_569),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_338),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_273),
.B(n_334),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g338 ( 
.A(n_27),
.B(n_339),
.C(n_341),
.Y(n_338)
);

AOI22x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_191),
.B1(n_227),
.B2(n_269),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_29),
.B(n_192),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_115),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_30),
.B(n_271),
.C(n_272),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_78),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_55),
.Y(n_31)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_32),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_44),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_33),
.A2(n_50),
.B(n_262),
.C(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.C(n_40),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_34),
.A2(n_37),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_34),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_34),
.A2(n_111),
.B1(n_204),
.B2(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_37),
.A2(n_112),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_37),
.B(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_37),
.B(n_359),
.Y(n_383)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_39),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_40),
.A2(n_110),
.B1(n_113),
.B2(n_114),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_40),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_40),
.Y(n_498)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_42),
.Y(n_210)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_42),
.Y(n_243)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_42),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_45),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_45),
.B(n_54),
.Y(n_263)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_49),
.Y(n_332)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_50),
.A2(n_54),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_50),
.A2(n_54),
.B1(n_81),
.B2(n_489),
.Y(n_565)
);

NOR3xp33_ASAP7_75t_L g569 ( 
.A(n_50),
.B(n_81),
.C(n_467),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_52),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_52),
.Y(n_247)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_52),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_54),
.B(n_253),
.C(n_519),
.Y(n_518)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_55),
.B(n_78),
.C(n_268),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_68),
.C(n_73),
.Y(n_55)
);

INVxp67_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

XNOR2x1_ASAP7_75t_L g146 ( 
.A(n_57),
.B(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.C(n_65),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_59),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_62),
.B(n_65),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_63),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_65),
.B(n_184),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g363 ( 
.A1(n_65),
.A2(n_183),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_65),
.B(n_365),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_69),
.A2(n_75),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_71),
.Y(n_388)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_77),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_94),
.C(n_109),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_79),
.A2(n_80),
.B1(n_94),
.B2(n_95),
.Y(n_223)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

OAI22x1_ASAP7_75t_L g179 ( 
.A1(n_81),
.A2(n_91),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_81),
.A2(n_197),
.B1(n_199),
.B2(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_81),
.Y(n_489)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2x1_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_87),
.B(n_91),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_87),
.Y(n_181)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_89),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.C(n_106),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2x2_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_98),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_99),
.Y(n_435)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_102),
.B(n_242),
.C(n_491),
.Y(n_528)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_103),
.A2(n_245),
.B1(n_246),
.B2(n_248),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_103),
.Y(n_248)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_109),
.Y(n_222)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_111),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_112),
.B(n_174),
.C(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_113),
.A2(n_494),
.B1(n_495),
.B2(n_498),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_170),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_145),
.C(n_150),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_117),
.B(n_145),
.C(n_150),
.Y(n_271)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_118),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_132),
.C(n_142),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_119),
.B(n_142),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.C(n_127),
.Y(n_119)
);

XNOR2x1_ASAP7_75t_L g280 ( 
.A(n_120),
.B(n_172),
.Y(n_280)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_123),
.Y(n_254)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_126),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_127),
.B(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_130),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_132),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.C(n_138),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_133),
.B(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_136),
.B(n_138),
.Y(n_202)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_138),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_138),
.A2(n_197),
.B1(n_199),
.B2(n_466),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_138),
.A2(n_466),
.B1(n_525),
.B2(n_526),
.Y(n_524)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_140),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_141),
.Y(n_327)
);

BUFx2_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_146),
.B(n_151),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.C(n_164),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_152),
.A2(n_153),
.B1(n_157),
.B2(n_158),
.Y(n_219)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_164),
.B(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_164),
.A2(n_282),
.B(n_285),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_168),
.Y(n_286)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_169),
.Y(n_474)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_170),
.Y(n_272)
);

XOR2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_171),
.B(n_179),
.C(n_182),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_176),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_177),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_183),
.A2(n_184),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_189),
.C(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_184),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_184),
.B(n_214),
.C(n_235),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_186),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_188),
.B(n_506),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_190),
.B(n_197),
.C(n_466),
.Y(n_484)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_220),
.C(n_224),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_193),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.C(n_217),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_194),
.B(n_218),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g562 ( 
.A(n_197),
.B(n_489),
.C(n_490),
.Y(n_562)
);

XOR2x2_ASAP7_75t_SL g276 ( 
.A(n_200),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.C(n_206),
.Y(n_200)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_201),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_203),
.B(n_207),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_204),
.Y(n_319)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.C(n_214),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_208),
.A2(n_214),
.B1(n_215),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_208),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_211),
.B(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_215),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_214),
.A2(n_215),
.B1(n_467),
.B2(n_527),
.Y(n_526)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_215),
.B(n_466),
.C(n_467),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_216),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_221),
.B(n_225),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NOR2xp67_ASAP7_75t_L g335 ( 
.A(n_228),
.B(n_270),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_228),
.B(n_270),
.Y(n_337)
);

XNOR2x1_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_267),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_250),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_230),
.Y(n_549)
);

XOR2x2_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_238),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_231),
.B(n_239),
.C(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_249),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g513 ( 
.A(n_241),
.Y(n_513)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_246),
.Y(n_491)
);

INVxp33_ASAP7_75t_SL g550 ( 
.A(n_250),
.Y(n_550)
);

OAI22x1_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_250)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_261),
.Y(n_251)
);

INVxp33_ASAP7_75t_SL g539 ( 
.A(n_252),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_257),
.Y(n_519)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g540 ( 
.A(n_261),
.Y(n_540)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_265),
.B(n_539),
.C(n_540),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_267),
.A2(n_548),
.B(n_551),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_301),
.B(n_333),
.Y(n_273)
);

NOR2x1_ASAP7_75t_L g339 ( 
.A(n_274),
.B(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_299),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_275),
.B(n_299),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.C(n_296),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_296),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.C(n_287),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_287),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.C(n_291),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_289),
.B(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_290),
.B(n_291),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx5_ASAP7_75t_L g324 ( 
.A(n_295),
.Y(n_324)
);

XNOR2x2_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_304),
.Y(n_340)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_308),
.C(n_312),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_306),
.B(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_313),
.Y(n_344)
);

XNOR2x1_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.C(n_320),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_314),
.B(n_348),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_317),
.A2(n_318),
.B1(n_320),
.B2(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_325),
.C(n_328),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_321),
.A2(n_322),
.B1(n_328),
.B2(n_329),
.Y(n_449)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_324),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_325),
.B(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B(n_337),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_366),
.B(n_457),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_345),
.Y(n_342)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_343),
.Y(n_458)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_346),
.B(n_458),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_350),
.C(n_353),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_347),
.B(n_453),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_350),
.A2(n_351),
.B1(n_353),
.B2(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_353),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.C(n_363),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_354),
.A2(n_355),
.B1(n_363),
.B2(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_357),
.B(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_363),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_451),
.B(n_456),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_440),
.B(n_450),
.Y(n_367)
);

AOI21x1_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_410),
.B(n_439),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_402),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_384),
.B1(n_400),
.B2(n_401),
.Y(n_370)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_371),
.Y(n_400)
);

AOI221xp5_ASAP7_75t_L g439 ( 
.A1(n_371),
.A2(n_384),
.B1(n_400),
.B2(n_401),
.C(n_402),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_373),
.B1(n_382),
.B2(n_383),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_372),
.B(n_383),
.C(n_401),
.Y(n_441)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_378),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_378),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

INVx8_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx8_ASAP7_75t_L g420 ( 
.A(n_377),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx6_ASAP7_75t_L g417 ( 
.A(n_381),
.Y(n_417)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_384),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_389),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_385),
.B(n_390),
.C(n_394),
.Y(n_447)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_394),
.B1(n_398),
.B2(n_399),
.Y(n_389)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_390),
.Y(n_398)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_394),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_405),
.C(n_406),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_403),
.A2(n_404),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_405),
.A2(n_406),
.B1(n_407),
.B2(n_424),
.Y(n_423)
);

CKINVDCx12_ASAP7_75t_R g424 ( 
.A(n_405),
.Y(n_424)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_425),
.B(n_438),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_421),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_421),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_418),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_418),
.Y(n_427)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx5_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_431),
.B(n_437),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_427),
.B(n_428),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_436),
.Y(n_431)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_441),
.B(n_442),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_446),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_443),
.B(n_447),
.C(n_448),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_455),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_SL g456 ( 
.A(n_452),
.B(n_455),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_530),
.Y(n_459)
);

OAI211xp5_ASAP7_75t_L g552 ( 
.A1(n_460),
.A2(n_553),
.B(n_556),
.C(n_557),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_510),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_461),
.B(n_510),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_492),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_479),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_463),
.B(n_479),
.C(n_492),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_470),
.C(n_475),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_465),
.B(n_508),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_467),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_467),
.A2(n_527),
.B1(n_564),
.B2(n_565),
.Y(n_563)
);

BUFx4f_ASAP7_75t_SL g467 ( 
.A(n_468),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_471),
.A2(n_475),
.B1(n_476),
.B2(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_471),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_487),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_484),
.B1(n_485),
.B2(n_486),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_481),
.Y(n_485)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_484),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_484),
.B(n_485),
.C(n_487),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_488),
.B(n_490),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_R g492 ( 
.A(n_493),
.B(n_504),
.C(n_507),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_493),
.B(n_505),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_498),
.C(n_499),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_499),
.Y(n_515)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_507),
.B(n_522),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_520),
.C(n_523),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_542),
.Y(n_541)
);

MAJx2_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_514),
.C(n_517),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_512),
.B(n_535),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_518),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_521),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_523),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_528),
.C(n_529),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_529),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_544),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_531),
.A2(n_554),
.B(n_555),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_541),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_532),
.B(n_541),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_536),
.C(n_538),
.Y(n_532)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_534),
.B(n_546),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_538),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_545),
.B(n_547),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_545),
.B(n_547),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_550),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_549),
.B(n_550),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g557 ( 
.A(n_558),
.B(n_561),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_568),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_567),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_561),
.A2(n_562),
.B1(n_563),
.B2(n_566),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_563),
.Y(n_566)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);


endmodule