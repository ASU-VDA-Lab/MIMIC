module fake_jpeg_31616_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_1),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_59),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_1),
.Y(n_79)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_69),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_68),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_79),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_43),
.B1(n_52),
.B2(n_50),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_58),
.B1(n_56),
.B2(n_55),
.Y(n_91)
);

HAxp5_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_47),
.CON(n_72),
.SN(n_72)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_2),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_47),
.C(n_49),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_89),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_96),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_54),
.B1(n_46),
.B2(n_4),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_98),
.B1(n_6),
.B2(n_7),
.Y(n_111)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_53),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_104),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_73),
.B(n_82),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_22),
.B(n_24),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_98),
.A3(n_85),
.B1(n_97),
.B2(n_53),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_28),
.B(n_30),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_3),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_109),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

NOR3xp33_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_5),
.C(n_6),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_8),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_114),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_15),
.A3(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_35),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_122),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_127),
.B1(n_112),
.B2(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_103),
.C(n_113),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_134),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_117),
.B1(n_124),
.B2(n_129),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_137),
.A2(n_130),
.B(n_128),
.C(n_121),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_137),
.C(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_136),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_141),
.B(n_121),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_134),
.B(n_138),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_127),
.Y(n_146)
);


endmodule