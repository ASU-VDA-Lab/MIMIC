module real_jpeg_15359_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_0),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_581),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_1),
.B(n_582),
.Y(n_581)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_2),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_2),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_2),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g498 ( 
.A(n_3),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_4),
.A2(n_101),
.B1(n_104),
.B2(n_105),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_4),
.A2(n_104),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_4),
.A2(n_104),
.B1(n_213),
.B2(n_218),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_4),
.A2(n_104),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_5),
.A2(n_273),
.B1(n_275),
.B2(n_276),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_5),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_5),
.A2(n_275),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g462 ( 
.A1(n_5),
.A2(n_275),
.B1(n_463),
.B2(n_464),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_5),
.A2(n_275),
.B1(n_519),
.B2(n_522),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_6),
.A2(n_37),
.B1(n_42),
.B2(n_44),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_6),
.A2(n_44),
.B1(n_146),
.B2(n_149),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_6),
.A2(n_44),
.B1(n_267),
.B2(n_270),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_6),
.A2(n_44),
.B1(n_343),
.B2(n_346),
.Y(n_342)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_7),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_7),
.Y(n_180)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_7),
.Y(n_252)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_8),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_8),
.Y(n_158)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_8),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_8),
.Y(n_461)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_8),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_9),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_9),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_9),
.A2(n_93),
.B1(n_182),
.B2(n_185),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_9),
.A2(n_93),
.B1(n_201),
.B2(n_204),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_9),
.A2(n_93),
.B1(n_226),
.B2(n_229),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_10),
.Y(n_582)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_11),
.Y(n_339)
);

OAI32xp33_ASAP7_75t_L g322 ( 
.A1(n_12),
.A2(n_323),
.A3(n_326),
.B1(n_329),
.B2(n_336),
.Y(n_322)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_12),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_12),
.A2(n_335),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_12),
.B(n_26),
.Y(n_400)
);

OAI32xp33_ASAP7_75t_L g437 ( 
.A1(n_12),
.A2(n_438),
.A3(n_442),
.B1(n_443),
.B2(n_446),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g467 ( 
.A1(n_12),
.A2(n_335),
.B1(n_468),
.B2(n_469),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_12),
.B(n_110),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_12),
.B(n_172),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_12),
.B(n_66),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_13),
.A2(n_298),
.B1(n_301),
.B2(n_302),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_13),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_13),
.A2(n_301),
.B1(n_403),
.B2(n_407),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_13),
.A2(n_301),
.B1(n_508),
.B2(n_514),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_13),
.A2(n_301),
.B1(n_543),
.B2(n_547),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_14),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_15),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_15),
.A2(n_50),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_15),
.A2(n_50),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_15),
.A2(n_50),
.B1(n_255),
.B2(n_260),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_16),
.Y(n_176)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_16),
.Y(n_184)
);

BUFx4f_ASAP7_75t_L g259 ( 
.A(n_16),
.Y(n_259)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_237),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_235),
.Y(n_20)
);

NAND2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_207),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_22),
.B(n_207),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_141),
.C(n_165),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_23),
.A2(n_141),
.B1(n_142),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_23),
.Y(n_285)
);

XNOR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_64),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_24),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_36),
.B(n_45),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_25),
.A2(n_36),
.B1(n_53),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_25),
.A2(n_53),
.B1(n_297),
.B2(n_361),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_25),
.A2(n_53),
.B1(n_272),
.B2(n_305),
.Y(n_386)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_26),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_26),
.B(n_46),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_26),
.B(n_200),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_26),
.A2(n_52),
.B1(n_296),
.B2(n_304),
.Y(n_295)
);

AO22x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_26)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_27),
.Y(n_473)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_28),
.Y(n_408)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_28),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_29),
.Y(n_228)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_29),
.Y(n_320)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_33),
.Y(n_138)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_39),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_40),
.Y(n_217)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_40),
.Y(n_274)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_40),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_41),
.Y(n_203)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_43),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.Y(n_45)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_53),
.A2(n_199),
.B(n_206),
.Y(n_198)
);

OAI21x1_ASAP7_75t_SL g271 ( 
.A1(n_53),
.A2(n_272),
.B(n_278),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_58),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g309 ( 
.A(n_59),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_99),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_65),
.A2(n_220),
.B1(n_221),
.B2(n_232),
.Y(n_219)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_65),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_65),
.B(n_209),
.C(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_77),
.B(n_88),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_66),
.B(n_156),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_66),
.B(n_266),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_66),
.A2(n_77),
.B1(n_504),
.B2(n_507),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_66),
.A2(n_77),
.B1(n_456),
.B2(n_507),
.Y(n_526)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_67),
.B(n_89),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_67),
.A2(n_189),
.B1(n_195),
.B2(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_67),
.A2(n_195),
.B1(n_455),
.B2(n_462),
.Y(n_454)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B1(n_73),
.B2(n_76),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_70),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_70),
.Y(n_501)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_77),
.B(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_77),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_77),
.A2(n_164),
.B(n_478),
.Y(n_477)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_84),
.B2(n_86),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_80),
.Y(n_490)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_81),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_81),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g494 ( 
.A(n_83),
.Y(n_494)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_86),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_86),
.B(n_335),
.Y(n_495)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_87),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_89),
.A2(n_195),
.B(n_196),
.Y(n_359)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_92),
.Y(n_194)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_97),
.Y(n_442)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_99),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_108),
.B(n_134),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_108),
.B1(n_110),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_103),
.Y(n_370)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_108),
.B(n_136),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_108),
.A2(n_223),
.B(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_109),
.A2(n_145),
.B1(n_224),
.B2(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_109),
.A2(n_224),
.B1(n_313),
.B2(n_366),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_109),
.A2(n_135),
.B(n_225),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_109),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_109),
.A2(n_224),
.B1(n_402),
.B2(n_467),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_121),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_110),
.Y(n_224)
);

AO22x2_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_115),
.B1(n_116),
.B2(n_118),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_117),
.Y(n_269)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_117),
.Y(n_458)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_126),
.B1(n_128),
.B2(n_131),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_136),
.Y(n_281)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_142),
.A2(n_143),
.B(n_153),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_153),
.Y(n_142)
);

INVxp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_148),
.Y(n_334)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_164),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_155),
.B(n_376),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_165),
.A2(n_166),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_186),
.B(n_197),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_167),
.A2(n_168),
.B1(n_197),
.B2(n_198),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_167),
.A2(n_168),
.B1(n_188),
.B2(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2x1_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_173),
.B(n_181),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_171),
.A2(n_173),
.B1(n_335),
.B2(n_542),
.Y(n_541)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_173),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_173),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_173),
.A2(n_518),
.B(n_524),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_173),
.A2(n_532),
.B1(n_542),
.B2(n_555),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_176),
.Y(n_348)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_178),
.B(n_254),
.Y(n_374)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_179),
.Y(n_557)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_181),
.B(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_181),
.Y(n_453)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_182),
.Y(n_352)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_183),
.Y(n_523)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_183),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_184),
.Y(n_357)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_185),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_187),
.B(n_241),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_188),
.Y(n_419)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_195),
.B(n_196),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_192),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_203),
.Y(n_300)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_233),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_219),
.Y(n_210)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_231),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_224),
.Y(n_410)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_226),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_228),
.Y(n_325)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_229),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_230),
.Y(n_371)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_230),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_286),
.B(n_580),
.Y(n_237)
);

NOR2xp67_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_282),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_239),
.B(n_282),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.C(n_244),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_240),
.A2(n_242),
.B1(n_243),
.B2(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_240),
.Y(n_431)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_244),
.B(n_430),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_271),
.C(n_279),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_L g420 ( 
.A(n_245),
.B(n_421),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_264),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_246),
.B(n_264),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_253),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_247),
.Y(n_524)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_250),
.Y(n_398)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_250),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_252),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_253),
.A2(n_342),
.B(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_259),
.Y(n_345)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_259),
.Y(n_521)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_259),
.Y(n_546)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx2_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_271),
.B(n_280),
.Y(n_421)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_273),
.Y(n_337)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_574),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_432),
.Y(n_288)
);

NOR3xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_413),
.C(n_427),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_388),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_377),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_292),
.B(n_377),
.C(n_576),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_358),
.C(n_372),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_293),
.B(n_412),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_321),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_311),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_295),
.B(n_311),
.C(n_321),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_300),
.Y(n_364)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_303),
.A2(n_306),
.B1(n_307),
.B2(n_310),
.Y(n_305)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_306),
.A2(n_310),
.B1(n_367),
.B2(n_371),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_306),
.A2(n_310),
.B1(n_457),
.B2(n_459),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_306),
.A2(n_310),
.B1(n_353),
.B2(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_309),
.Y(n_362)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_318),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_340),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_322),
.B(n_340),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_335),
.B(n_444),
.Y(n_443)
);

OAI21xp33_ASAP7_75t_SL g504 ( 
.A1(n_335),
.A2(n_495),
.B(n_505),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_349),
.B2(n_351),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_341),
.A2(n_351),
.B(n_374),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_341),
.A2(n_374),
.B(n_453),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_341),
.A2(n_531),
.B1(n_535),
.B2(n_536),
.Y(n_530)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_345),
.Y(n_547)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_355),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_358),
.B(n_372),
.Y(n_412)
);

MAJx2_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.C(n_365),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_365),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_366),
.A2(n_402),
.B1(n_409),
.B2(n_410),
.Y(n_401)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_375),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_375),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_381),
.C(n_387),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_381),
.B1(n_382),
.B2(n_387),
.Y(n_379)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_380),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_382),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_383),
.B(n_424),
.C(n_425),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_385),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_386),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_411),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_389),
.B(n_411),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_392),
.C(n_394),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_390),
.B(n_570),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_392),
.A2(n_393),
.B1(n_394),
.B2(n_571),
.Y(n_570)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_394),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_399),
.C(n_401),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_395),
.A2(n_399),
.B1(n_400),
.B2(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_395),
.Y(n_482)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_401),
.B(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g574 ( 
.A1(n_414),
.A2(n_575),
.B(n_577),
.C(n_578),
.D(n_579),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_415),
.B(n_416),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_422),
.B1(n_423),
.B2(n_426),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_417),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_420),
.C(n_422),
.Y(n_428)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_427),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_428),
.B(n_429),
.Y(n_579)
);

OAI21x1_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_568),
.B(n_573),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_484),
.B(n_567),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_474),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_435),
.B(n_474),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_454),
.C(n_466),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_436),
.B(n_565),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_452),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_437),
.B(n_452),
.Y(n_476)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_454),
.B(n_466),
.Y(n_565)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_462),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_463),
.Y(n_506)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_475),
.A2(n_479),
.B1(n_480),
.B2(n_483),
.Y(n_474)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_475),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_476),
.B(n_477),
.C(n_479),
.Y(n_572)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_562),
.B(n_566),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_528),
.B(n_561),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_516),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_487),
.B(n_516),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_502),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_488),
.A2(n_502),
.B1(n_503),
.B2(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_488),
.Y(n_538)
);

OAI32xp33_ASAP7_75t_L g488 ( 
.A1(n_489),
.A2(n_491),
.A3(n_492),
.B1(n_495),
.B2(n_496),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_499),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_525),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_517),
.B(n_526),
.C(n_527),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_518),
.Y(n_535)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_527),
.Y(n_525)
);

OAI21x1_ASAP7_75t_SL g528 ( 
.A1(n_529),
.A2(n_539),
.B(n_560),
.Y(n_528)
);

NOR2x1_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_537),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_530),
.B(n_537),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_540),
.A2(n_553),
.B(n_559),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_548),
.Y(n_540)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_552),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_554),
.B(n_558),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_554),
.B(n_558),
.Y(n_559)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx5_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_564),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_563),
.B(n_564),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_569),
.B(n_572),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_569),
.B(n_572),
.Y(n_573)
);


endmodule