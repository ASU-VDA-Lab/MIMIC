module fake_jpeg_9348_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_29),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g39 ( 
.A1(n_17),
.A2(n_30),
.B(n_26),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_30),
.B(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_28),
.B1(n_23),
.B2(n_21),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_49),
.B1(n_55),
.B2(n_57),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_17),
.B1(n_22),
.B2(n_26),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_68),
.B1(n_31),
.B2(n_24),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_56),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_65),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_34),
.B1(n_17),
.B2(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_34),
.B1(n_26),
.B2(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_69),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_23),
.B1(n_29),
.B2(n_30),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_31),
.B1(n_24),
.B2(n_19),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_24),
.B1(n_19),
.B2(n_33),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_71),
.A2(n_84),
.B1(n_91),
.B2(n_99),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_36),
.C(n_45),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_83),
.C(n_54),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_75),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_77),
.Y(n_114)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_78),
.A2(n_112),
.B1(n_27),
.B2(n_18),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_79),
.A2(n_90),
.B1(n_110),
.B2(n_76),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_44),
.B1(n_43),
.B2(n_32),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_80),
.A2(n_57),
.B1(n_49),
.B2(n_66),
.Y(n_119)
);

CKINVDCx10_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_82),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_36),
.C(n_45),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_31),
.B1(n_33),
.B2(n_11),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_88),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_46),
.A2(n_32),
.B1(n_44),
.B2(n_43),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_48),
.A2(n_12),
.B1(n_11),
.B2(n_13),
.Y(n_91)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_93),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_48),
.A2(n_18),
.B1(n_27),
.B2(n_35),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_59),
.B(n_65),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_25),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_107),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_50),
.A2(n_13),
.B1(n_15),
.B2(n_14),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_25),
.B(n_16),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_25),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_25),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_111),
.Y(n_129)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_55),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_115),
.A2(n_139),
.B(n_101),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_131),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_140),
.B1(n_90),
.B2(n_79),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_106),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_133),
.B(n_81),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_130),
.A2(n_141),
.B1(n_99),
.B2(n_98),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_0),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_45),
.C(n_44),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_138),
.C(n_74),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_45),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_43),
.B1(n_50),
.B2(n_27),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_85),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_144),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_73),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_152),
.B1(n_159),
.B2(n_163),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_108),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_149),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_80),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_150),
.C(n_153),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_93),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_108),
.Y(n_149)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_82),
.B1(n_72),
.B2(n_94),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_134),
.B1(n_113),
.B2(n_136),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_108),
.B1(n_104),
.B2(n_96),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_83),
.C(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_157),
.B(n_25),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_158),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_97),
.B1(n_75),
.B2(n_102),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_162),
.B1(n_121),
.B2(n_123),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_167),
.B(n_35),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_121),
.B1(n_137),
.B2(n_122),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_126),
.A2(n_106),
.B1(n_81),
.B2(n_77),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_166),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_125),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_168),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_95),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_111),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_0),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_170),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_45),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_130),
.A2(n_121),
.B1(n_131),
.B2(n_116),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_134),
.B1(n_136),
.B2(n_113),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_100),
.C(n_27),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_116),
.B(n_117),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_175),
.Y(n_200)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

AOI22x1_ASAP7_75t_R g178 ( 
.A1(n_151),
.A2(n_121),
.B1(n_139),
.B2(n_35),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_178),
.B(n_170),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_201),
.B1(n_171),
.B2(n_167),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_174),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_184),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_172),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_194),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_187),
.A2(n_189),
.B(n_193),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_198),
.Y(n_227)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_207),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_196),
.B(n_205),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_156),
.A2(n_120),
.B1(n_89),
.B2(n_87),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_197),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_165),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_160),
.A2(n_35),
.B1(n_127),
.B2(n_25),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_161),
.B(n_189),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_154),
.B(n_14),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_204),
.B(n_169),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_159),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_152),
.B(n_0),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_147),
.B(n_25),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_219),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_214),
.B(n_220),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_224),
.B1(n_231),
.B2(n_179),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_167),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_192),
.Y(n_237)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_150),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_228),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_180),
.A2(n_158),
.B1(n_173),
.B2(n_155),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_149),
.B(n_146),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_153),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_230),
.C(n_188),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_176),
.B(n_166),
.Y(n_229)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_191),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_173),
.B1(n_16),
.B2(n_2),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_176),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_233),
.Y(n_257)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

BUFx12f_ASAP7_75t_SL g234 ( 
.A(n_182),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_235),
.B1(n_204),
.B2(n_183),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_210),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_241),
.C(n_244),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_191),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_195),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_220),
.Y(n_269)
);

AOI221xp5_ASAP7_75t_L g264 ( 
.A1(n_243),
.A2(n_216),
.B1(n_234),
.B2(n_211),
.C(n_235),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_198),
.C(n_199),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_199),
.C(n_190),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_251),
.C(n_254),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_208),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_246),
.B(n_255),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_201),
.B1(n_185),
.B2(n_193),
.Y(n_250)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_179),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_177),
.C(n_206),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_213),
.A2(n_177),
.B1(n_194),
.B2(n_187),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_216),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_263),
.Y(n_280)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_231),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_264),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_214),
.B(n_227),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_272),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_248),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_275),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_270),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_220),
.Y(n_270)
);

BUFx12f_ASAP7_75t_SL g271 ( 
.A(n_239),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g281 ( 
.A1(n_271),
.A2(n_257),
.B(n_253),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_225),
.C(n_214),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_197),
.C(n_228),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_274),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_16),
.C(n_1),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_16),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_238),
.A2(n_0),
.B(n_1),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_247),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_260),
.B(n_254),
.CI(n_237),
.CON(n_278),
.SN(n_278)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_285),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_251),
.C(n_252),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_290),
.B(n_272),
.Y(n_294)
);

AO21x1_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_4),
.B(n_5),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_256),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_286),
.C(n_267),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_250),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_259),
.A2(n_236),
.B(n_249),
.Y(n_287)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_258),
.C(n_273),
.Y(n_292)
);

XOR2x2_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_2),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_274),
.B(n_4),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_293),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_296),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_303),
.B(n_5),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_267),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_263),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_300),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_280),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_265),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_265),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_302),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_2),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_279),
.B1(n_286),
.B2(n_278),
.Y(n_304)
);

AND5x1_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_311),
.C(n_6),
.D(n_7),
.E(n_8),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_296),
.B(n_277),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_308),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_310),
.C(n_307),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_280),
.Y(n_310)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_299),
.C(n_282),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_316),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_305),
.A2(n_303),
.B(n_282),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_318),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_5),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_311),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_6),
.Y(n_320)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_312),
.A3(n_307),
.B1(n_310),
.B2(n_8),
.C1(n_9),
.C2(n_6),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_316),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_323),
.A2(n_322),
.B(n_319),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_324),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_8),
.Y(n_327)
);


endmodule