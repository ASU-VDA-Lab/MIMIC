module fake_jpeg_12037_n_611 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_611);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_611;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx5_ASAP7_75t_SL g212 ( 
.A(n_62),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_11),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_63),
.B(n_67),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_60),
.Y(n_65)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_66),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_29),
.B(n_10),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_70),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_76),
.Y(n_209)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_60),
.Y(n_77)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_78),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_79),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_80),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_21),
.B(n_10),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_81),
.B(n_84),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_82),
.Y(n_161)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g185 ( 
.A(n_83),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_29),
.B(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_46),
.Y(n_88)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_92),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_93),
.Y(n_190)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_94),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_96),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_20),
.B(n_10),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_30),
.B(n_10),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_103),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_30),
.B(n_12),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_25),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_27),
.Y(n_114)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_34),
.Y(n_115)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

INVx4_ASAP7_75t_SL g119 ( 
.A(n_25),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_119),
.B(n_36),
.Y(n_208)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_43),
.B(n_9),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_28),
.Y(n_126)
);

BUFx2_ASAP7_75t_R g153 ( 
.A(n_126),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_128),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_59),
.B(n_9),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_124),
.B(n_59),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_129),
.B(n_173),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_58),
.B1(n_40),
.B2(n_51),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_131),
.A2(n_152),
.B1(n_161),
.B2(n_159),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_43),
.B1(n_48),
.B2(n_51),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_134),
.A2(n_138),
.B1(n_150),
.B2(n_166),
.Y(n_227)
);

BUFx4f_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_135),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_48),
.B1(n_39),
.B2(n_50),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_83),
.A2(n_31),
.B1(n_55),
.B2(n_58),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_72),
.A2(n_40),
.B1(n_41),
.B2(n_50),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_128),
.B(n_63),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_162),
.B(n_167),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_89),
.A2(n_121),
.B1(n_125),
.B2(n_79),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_99),
.B(n_42),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_104),
.B(n_42),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_71),
.B(n_55),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_176),
.B(n_186),
.Y(n_228)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_88),
.Y(n_184)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_69),
.B(n_31),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_64),
.Y(n_187)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_187),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_65),
.B(n_41),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_191),
.B(n_200),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_119),
.B(n_26),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_66),
.A2(n_70),
.B1(n_95),
.B2(n_93),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_201),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_263)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_74),
.A2(n_56),
.B1(n_26),
.B2(n_35),
.Y(n_204)
);

AO22x1_ASAP7_75t_SL g235 ( 
.A1(n_204),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_107),
.Y(n_205)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_112),
.Y(n_206)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_206),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_208),
.Y(n_244)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_76),
.Y(n_210)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_214),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_145),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_215),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_146),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_216),
.A2(n_218),
.B1(n_225),
.B2(n_230),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_126),
.B(n_36),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_217),
.A2(n_238),
.B(n_255),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_132),
.A2(n_36),
.B1(n_35),
.B2(n_28),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_150),
.A2(n_101),
.B1(n_97),
.B2(n_96),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_220),
.A2(n_245),
.B1(n_247),
.B2(n_271),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_158),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_221),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_35),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_223),
.B(n_243),
.C(n_256),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_155),
.A2(n_28),
.B1(n_82),
.B2(n_14),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_226),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_153),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_229),
.B(n_237),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_155),
.A2(n_8),
.B1(n_17),
.B2(n_16),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_232),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_233),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_201),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_234),
.A2(n_252),
.B1(n_263),
.B2(n_279),
.Y(n_289)
);

OA22x2_ASAP7_75t_L g325 ( 
.A1(n_235),
.A2(n_234),
.B1(n_270),
.B2(n_255),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_189),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_SL g238 ( 
.A(n_191),
.B(n_199),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_197),
.A2(n_181),
.B1(n_130),
.B2(n_204),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_239),
.Y(n_291)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_241),
.Y(n_341)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_195),
.Y(n_242)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_242),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_141),
.B(n_1),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_204),
.A2(n_13),
.B1(n_4),
.B2(n_6),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_246),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_131),
.A2(n_152),
.B1(n_149),
.B2(n_165),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_135),
.Y(n_248)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_248),
.Y(n_300)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_190),
.Y(n_249)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_249),
.Y(n_309)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_137),
.A2(n_2),
.B1(n_18),
.B2(n_6),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_253),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_137),
.B(n_4),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_254),
.B(n_257),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_147),
.A2(n_4),
.B1(n_8),
.B2(n_15),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_141),
.B(n_8),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_160),
.B(n_8),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_179),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_259),
.B(n_281),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_157),
.A2(n_172),
.B1(n_180),
.B2(n_168),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_260),
.A2(n_262),
.B(n_228),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_176),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_265),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

INVx4_ASAP7_75t_SL g314 ( 
.A(n_262),
.Y(n_314)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_185),
.Y(n_264)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_264),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_189),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_142),
.B(n_15),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_266),
.B(n_268),
.C(n_269),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_267),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_144),
.B(n_154),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_164),
.B(n_17),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_212),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_270),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_163),
.A2(n_185),
.B1(n_194),
.B2(n_170),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_194),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_273),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_186),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_192),
.Y(n_276)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_276),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_136),
.B(n_160),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_257),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_178),
.Y(n_278)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_136),
.A2(n_175),
.B1(n_211),
.B2(n_209),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_280),
.A2(n_182),
.B1(n_140),
.B2(n_151),
.Y(n_288)
);

INVx4_ASAP7_75t_SL g281 ( 
.A(n_203),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_188),
.Y(n_282)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_282),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_178),
.Y(n_283)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_283),
.Y(n_342)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_196),
.Y(n_284)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_284),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_175),
.A2(n_174),
.B1(n_177),
.B2(n_156),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_161),
.B1(n_139),
.B2(n_213),
.Y(n_299)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_133),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_286),
.Y(n_307)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_143),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_287),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_288),
.A2(n_313),
.B1(n_317),
.B2(n_215),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_299),
.A2(n_327),
.B1(n_335),
.B2(n_298),
.Y(n_361)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_250),
.A2(n_213),
.B(n_169),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_302),
.B(n_331),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_280),
.A2(n_227),
.B1(n_244),
.B2(n_217),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_222),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_316),
.B(n_322),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_244),
.A2(n_139),
.B1(n_202),
.B2(n_235),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_238),
.B(n_236),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_319),
.B(n_248),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_254),
.B(n_252),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_321),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_268),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_323),
.A2(n_260),
.B(n_269),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_333),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_268),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_326),
.B(n_328),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_270),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_327),
.A2(n_344),
.B(n_219),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_270),
.Y(n_328)
);

OA22x2_ASAP7_75t_L g333 ( 
.A1(n_235),
.A2(n_264),
.B1(n_284),
.B2(n_282),
.Y(n_333)
);

AND2x2_ASAP7_75t_SL g366 ( 
.A(n_333),
.B(n_317),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_281),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_335),
.B(n_338),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g338 ( 
.A(n_256),
.B(n_243),
.CI(n_223),
.CON(n_338),
.SN(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_224),
.B(n_267),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_339),
.B(n_287),
.Y(n_358)
);

MAJx2_ASAP7_75t_L g343 ( 
.A(n_256),
.B(n_243),
.C(n_223),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_266),
.C(n_275),
.Y(n_348)
);

O2A1O1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_269),
.A2(n_266),
.B(n_258),
.C(n_274),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_348),
.B(n_388),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_349),
.B(n_365),
.Y(n_425)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_320),
.Y(n_350)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_350),
.Y(n_401)
);

OAI32xp33_ASAP7_75t_L g351 ( 
.A1(n_292),
.A2(n_246),
.A3(n_241),
.B1(n_226),
.B2(n_240),
.Y(n_351)
);

XOR2x2_ASAP7_75t_L g420 ( 
.A(n_351),
.B(n_300),
.Y(n_420)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_296),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_353),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_308),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_355),
.B(n_358),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_291),
.A2(n_249),
.B1(n_253),
.B2(n_219),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_356),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_357),
.B(n_314),
.Y(n_400)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_320),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_362),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_361),
.A2(n_366),
.B1(n_372),
.B2(n_384),
.Y(n_413)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_340),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_231),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_363),
.B(n_364),
.C(n_373),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_232),
.C(n_286),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_340),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_313),
.A2(n_283),
.B1(n_278),
.B2(n_251),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_367),
.A2(n_369),
.B1(n_374),
.B2(n_390),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_305),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_376),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_312),
.A2(n_221),
.B1(n_233),
.B2(n_276),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_290),
.A2(n_259),
.B(n_242),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_370),
.A2(n_314),
.B(n_332),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_289),
.A2(n_214),
.B1(n_327),
.B2(n_290),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_306),
.B(n_329),
.C(n_326),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_325),
.A2(n_289),
.B1(n_322),
.B2(n_333),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_306),
.B(n_329),
.C(n_323),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_375),
.B(n_379),
.Y(n_419)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_297),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_345),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_377),
.Y(n_424)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_345),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_378),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_292),
.B(n_321),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_325),
.A2(n_333),
.B1(n_328),
.B2(n_298),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_380),
.Y(n_398)
);

OAI21xp33_ASAP7_75t_SL g392 ( 
.A1(n_381),
.A2(n_341),
.B(n_315),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_304),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_382),
.B(n_385),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_321),
.A2(n_325),
.B1(n_318),
.B2(n_344),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_338),
.A2(n_294),
.B1(n_342),
.B2(n_334),
.Y(n_385)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_337),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_386),
.B(n_389),
.Y(n_407)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_295),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_387),
.B(n_350),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_338),
.B(n_304),
.C(n_295),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_307),
.B(n_311),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_307),
.A2(n_311),
.B1(n_342),
.B2(n_334),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_310),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_391),
.B(n_410),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_392),
.A2(n_395),
.B1(n_408),
.B2(n_361),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_374),
.A2(n_330),
.B1(n_310),
.B2(n_315),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_360),
.A2(n_304),
.B(n_314),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_396),
.A2(n_404),
.B(n_421),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_397),
.A2(n_422),
.B(n_382),
.Y(n_431)
);

OAI21xp33_ASAP7_75t_SL g451 ( 
.A1(n_400),
.A2(n_409),
.B(n_411),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_353),
.A2(n_309),
.B(n_337),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_349),
.A2(n_330),
.B1(n_296),
.B2(n_303),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_379),
.B(n_341),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_370),
.A2(n_293),
.B(n_324),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_412),
.A2(n_378),
.B(n_377),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_355),
.B(n_309),
.Y(n_414)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_414),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_368),
.B(n_300),
.Y(n_415)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_415),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_341),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_418),
.B(n_420),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_372),
.A2(n_324),
.B(n_332),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_360),
.A2(n_297),
.B(n_301),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_389),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_423),
.B(n_390),
.Y(n_455)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_427),
.Y(n_433)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_428),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_398),
.A2(n_384),
.B1(n_366),
.B2(n_385),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_429),
.A2(n_436),
.B1(n_448),
.B2(n_421),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_413),
.A2(n_367),
.B1(n_369),
.B2(n_366),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_430),
.A2(n_437),
.B1(n_442),
.B2(n_420),
.Y(n_473)
);

AO21x1_ASAP7_75t_L g462 ( 
.A1(n_431),
.A2(n_451),
.B(n_397),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_398),
.A2(n_346),
.B1(n_371),
.B2(n_357),
.Y(n_432)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_432),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_399),
.A2(n_366),
.B1(n_364),
.B2(n_346),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_413),
.A2(n_375),
.B1(n_373),
.B2(n_388),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_406),
.Y(n_438)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_438),
.Y(n_471)
);

INVx5_ASAP7_75t_L g439 ( 
.A(n_403),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_439),
.B(n_452),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_413),
.A2(n_354),
.B1(n_348),
.B2(n_347),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_363),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_443),
.B(n_446),
.C(n_447),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_407),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_444),
.B(n_445),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_407),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_354),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_417),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_399),
.A2(n_358),
.B1(n_359),
.B2(n_351),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_417),
.B(n_402),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_405),
.Y(n_463)
);

FAx1_ASAP7_75t_SL g450 ( 
.A(n_417),
.B(n_365),
.CI(n_387),
.CON(n_450),
.SN(n_450)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_450),
.B(n_396),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_393),
.Y(n_452)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_403),
.Y(n_454)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_454),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_455),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_456),
.A2(n_397),
.B(n_396),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_402),
.B(n_362),
.C(n_376),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_458),
.C(n_459),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_402),
.B(n_386),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_410),
.B(n_301),
.C(n_336),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_460),
.Y(n_469)
);

OAI32xp33_ASAP7_75t_L g461 ( 
.A1(n_405),
.A2(n_336),
.A3(n_296),
.B1(n_303),
.B2(n_352),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_395),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_462),
.A2(n_466),
.B(n_472),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_463),
.B(n_440),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_477),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_468),
.A2(n_481),
.B1(n_487),
.B2(n_465),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_431),
.A2(n_404),
.B(n_421),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_473),
.A2(n_474),
.B1(n_464),
.B2(n_479),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_430),
.A2(n_420),
.B1(n_392),
.B2(n_423),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_474),
.A2(n_479),
.B1(n_441),
.B2(n_448),
.Y(n_494)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_447),
.B(n_420),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_482),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_434),
.B(n_394),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_435),
.A2(n_412),
.B(n_391),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_478),
.B(n_485),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_455),
.A2(n_425),
.B1(n_391),
.B2(n_395),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_436),
.A2(n_404),
.B1(n_412),
.B2(n_394),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_449),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_453),
.B(n_415),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_422),
.C(n_393),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_486),
.B(n_457),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_429),
.A2(n_425),
.B1(n_416),
.B2(n_414),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_443),
.B(n_422),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_437),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_455),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_441),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_435),
.A2(n_400),
.B(n_425),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_492),
.B(n_456),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_494),
.A2(n_501),
.B1(n_507),
.B2(n_487),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_495),
.B(n_482),
.Y(n_536)
);

OAI21xp33_ASAP7_75t_L g496 ( 
.A1(n_467),
.A2(n_450),
.B(n_438),
.Y(n_496)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_496),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_498),
.B(n_462),
.Y(n_521)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_499),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_500),
.B(n_504),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_464),
.A2(n_428),
.B1(n_440),
.B2(n_433),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_442),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_505),
.B(n_463),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_469),
.B(n_433),
.Y(n_506)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_506),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_508),
.A2(n_513),
.B1(n_514),
.B2(n_473),
.Y(n_526)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_489),
.Y(n_509)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_509),
.Y(n_532)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_471),
.Y(n_510)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_510),
.Y(n_524)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_471),
.Y(n_511)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_511),
.Y(n_529)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_490),
.Y(n_512)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_512),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_468),
.A2(n_425),
.B1(n_408),
.B2(n_450),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_481),
.A2(n_459),
.B1(n_461),
.B2(n_426),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_469),
.B(n_427),
.Y(n_516)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_516),
.Y(n_541)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_484),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_467),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_485),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_518),
.B(n_519),
.Y(n_525)
);

FAx1_ASAP7_75t_SL g519 ( 
.A(n_476),
.B(n_418),
.CI(n_401),
.CON(n_519),
.SN(n_519)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_521),
.B(n_527),
.Y(n_543)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_522),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_526),
.A2(n_528),
.B1(n_494),
.B2(n_501),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_517),
.B(n_506),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_514),
.A2(n_475),
.B1(n_491),
.B2(n_470),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_533),
.A2(n_513),
.B1(n_502),
.B2(n_499),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_495),
.B(n_483),
.C(n_480),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_534),
.B(n_537),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_512),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g557 ( 
.A(n_535),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_536),
.B(n_539),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_500),
.B(n_483),
.C(n_486),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_538),
.B(n_493),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_510),
.B(n_470),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_520),
.A2(n_515),
.B(n_503),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_544),
.B(n_556),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_534),
.B(n_504),
.C(n_493),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_545),
.B(n_551),
.C(n_538),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_540),
.B(n_497),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_546),
.B(n_550),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_525),
.A2(n_515),
.B(n_508),
.Y(n_548)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_548),
.Y(n_565)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_549),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_521),
.B(n_505),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_537),
.B(n_536),
.C(n_530),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_552),
.A2(n_553),
.B1(n_533),
.B2(n_523),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_526),
.A2(n_502),
.B1(n_528),
.B2(n_531),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_554),
.B(n_530),
.Y(n_562)
);

AOI21x1_ASAP7_75t_L g555 ( 
.A1(n_539),
.A2(n_466),
.B(n_478),
.Y(n_555)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_555),
.Y(n_568)
);

INVxp33_ASAP7_75t_SL g556 ( 
.A(n_527),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_531),
.A2(n_472),
.B(n_492),
.Y(n_558)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_558),
.Y(n_573)
);

BUFx24_ASAP7_75t_SL g560 ( 
.A(n_542),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_560),
.B(n_547),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_561),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_562),
.B(n_563),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_543),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_567),
.B(n_570),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_545),
.B(n_532),
.C(n_488),
.Y(n_570)
);

CKINVDCx16_ASAP7_75t_R g571 ( 
.A(n_558),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_571),
.B(n_574),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_547),
.B(n_522),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_572),
.B(n_559),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_551),
.B(n_532),
.C(n_541),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_576),
.B(n_583),
.Y(n_589)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_577),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_569),
.A2(n_548),
.B(n_544),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_578),
.A2(n_581),
.B(n_585),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_570),
.B(n_552),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_580),
.B(n_572),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_569),
.A2(n_565),
.B(n_574),
.Y(n_581)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_566),
.Y(n_583)
);

AOI21x1_ASAP7_75t_L g585 ( 
.A1(n_573),
.A2(n_516),
.B(n_555),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_563),
.B(n_553),
.C(n_549),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_586),
.B(n_573),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_584),
.B(n_557),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_587),
.A2(n_582),
.B(n_580),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_586),
.B(n_561),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_588),
.B(n_595),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_592),
.B(n_593),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_579),
.B(n_550),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_594),
.B(n_575),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_577),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_596),
.B(n_599),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_598),
.A2(n_600),
.B(n_562),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_564),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_590),
.A2(n_568),
.B(n_582),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_601),
.A2(n_587),
.B(n_591),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_602),
.B(n_603),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_597),
.A2(n_592),
.B(n_564),
.Y(n_603)
);

AOI321xp33_ASAP7_75t_L g606 ( 
.A1(n_605),
.A2(n_524),
.A3(n_489),
.B1(n_554),
.B2(n_529),
.C(n_519),
.Y(n_606)
);

AOI21x1_ASAP7_75t_L g608 ( 
.A1(n_606),
.A2(n_604),
.B(n_519),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_608),
.A2(n_607),
.B(n_509),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_609),
.B(n_401),
.C(n_424),
.Y(n_610)
);

OAI321xp33_ASAP7_75t_L g611 ( 
.A1(n_610),
.A2(n_454),
.A3(n_439),
.B1(n_403),
.B2(n_293),
.C(n_303),
.Y(n_611)
);


endmodule