module fake_aes_6159_n_752 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_752);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_752;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g84 ( .A(n_44), .Y(n_84) );
BUFx5_ASAP7_75t_L g85 ( .A(n_48), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_11), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_4), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_40), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_34), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_18), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_61), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_71), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_70), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_5), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_14), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_24), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_39), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_31), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_24), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_50), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_25), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_80), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_11), .B(n_15), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_52), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_25), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_76), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_37), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_3), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_17), .Y(n_109) );
BUFx10_ASAP7_75t_L g110 ( .A(n_21), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_67), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_20), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_33), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_1), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_41), .Y(n_115) );
INVxp33_ASAP7_75t_L g116 ( .A(n_56), .Y(n_116) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_3), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_64), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_43), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_77), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_21), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_63), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_36), .Y(n_124) );
INVxp33_ASAP7_75t_L g125 ( .A(n_45), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_13), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_26), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_2), .Y(n_128) );
INVxp33_ASAP7_75t_SL g129 ( .A(n_62), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_10), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_0), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_19), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_28), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_8), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_133), .B(n_92), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_133), .B(n_1), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_85), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_115), .B(n_42), .Y(n_139) );
INVxp67_ASAP7_75t_L g140 ( .A(n_95), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_85), .Y(n_141) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_92), .A2(n_38), .B(n_82), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_95), .B(n_2), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_97), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_85), .B(n_4), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_85), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_97), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_100), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_100), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_116), .B(n_5), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g153 ( .A(n_93), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_85), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_115), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_85), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_85), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_99), .B(n_6), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_91), .Y(n_160) );
INVx5_ASAP7_75t_L g161 ( .A(n_110), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_104), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_111), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_109), .B(n_6), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_109), .B(n_7), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_113), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_117), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_118), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_125), .B(n_119), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_134), .B(n_9), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_120), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_122), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_124), .Y(n_174) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_127), .A2(n_10), .B(n_12), .Y(n_175) );
NAND2xp33_ASAP7_75t_L g176 ( .A(n_106), .B(n_51), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_87), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_90), .B(n_12), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_101), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_105), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_159), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_159), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_140), .A2(n_107), .B1(n_102), .B2(n_129), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_161), .B(n_94), .Y(n_185) );
INVx5_ASAP7_75t_L g186 ( .A(n_139), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_140), .A2(n_129), .B1(n_131), .B2(n_94), .Y(n_187) );
NAND3x1_ASAP7_75t_L g188 ( .A(n_168), .B(n_103), .C(n_114), .Y(n_188) );
BUFx8_ASAP7_75t_SL g189 ( .A(n_144), .Y(n_189) );
OR2x2_ASAP7_75t_L g190 ( .A(n_153), .B(n_131), .Y(n_190) );
AND2x6_ASAP7_75t_L g191 ( .A(n_159), .B(n_128), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_135), .B(n_123), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_135), .B(n_108), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_161), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_177), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_161), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_135), .B(n_132), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_161), .B(n_106), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_161), .B(n_110), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_161), .B(n_110), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_153), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_161), .B(n_121), .Y(n_203) );
INVx4_ASAP7_75t_L g204 ( .A(n_161), .Y(n_204) );
OAI22xp33_ASAP7_75t_SL g205 ( .A1(n_168), .A2(n_96), .B1(n_112), .B2(n_126), .Y(n_205) );
AND2x6_ASAP7_75t_L g206 ( .A(n_159), .B(n_89), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_135), .B(n_98), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_150), .B(n_89), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_159), .Y(n_209) );
NAND2xp33_ASAP7_75t_L g210 ( .A(n_139), .B(n_55), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_159), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_177), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_135), .B(n_130), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_177), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_155), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_150), .A2(n_130), .B1(n_126), .B2(n_86), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_165), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_177), .Y(n_221) );
BUFx4f_ASAP7_75t_L g222 ( .A(n_139), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_165), .Y(n_223) );
NAND2x1p5_ASAP7_75t_L g224 ( .A(n_144), .B(n_86), .Y(n_224) );
NOR2xp33_ASAP7_75t_SL g225 ( .A(n_139), .B(n_53), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_177), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_177), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_177), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_163), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_177), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_163), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_144), .Y(n_233) );
INVx4_ASAP7_75t_L g234 ( .A(n_139), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_163), .Y(n_235) );
INVx1_ASAP7_75t_SL g236 ( .A(n_151), .Y(n_236) );
AO22x2_ASAP7_75t_L g237 ( .A1(n_135), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_170), .B(n_16), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_170), .B(n_16), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_156), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_152), .B(n_17), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_156), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_148), .Y(n_243) );
INVx1_ASAP7_75t_SL g244 ( .A(n_151), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_142), .Y(n_245) );
AO22x2_ASAP7_75t_L g246 ( .A1(n_146), .A2(n_18), .B1(n_19), .B2(n_20), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_148), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_148), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_148), .Y(n_249) );
INVx4_ASAP7_75t_L g250 ( .A(n_139), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_198), .B(n_151), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_220), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_198), .B(n_137), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_241), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_236), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_244), .B(n_137), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_218), .Y(n_257) );
BUFx2_ASAP7_75t_L g258 ( .A(n_206), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_245), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_192), .B(n_178), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_233), .A2(n_166), .B1(n_171), .B2(n_150), .Y(n_261) );
INVx1_ASAP7_75t_SL g262 ( .A(n_202), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_218), .Y(n_263) );
NOR2x1_ASAP7_75t_R g264 ( .A(n_238), .B(n_166), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_220), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_220), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_191), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_215), .A2(n_171), .B1(n_152), .B2(n_164), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_191), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_191), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_198), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_215), .A2(n_176), .B1(n_167), .B2(n_169), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_238), .A2(n_160), .B1(n_164), .B2(n_167), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_238), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_192), .B(n_136), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_193), .B(n_136), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_239), .B(n_173), .Y(n_277) );
BUFx12f_ASAP7_75t_L g278 ( .A(n_239), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_206), .A2(n_176), .B1(n_169), .B2(n_173), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_239), .A2(n_160), .B1(n_174), .B2(n_175), .Y(n_280) );
OR2x6_ASAP7_75t_L g281 ( .A(n_237), .B(n_179), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_193), .B(n_149), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_243), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_247), .Y(n_284) );
BUFx8_ASAP7_75t_L g285 ( .A(n_206), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_207), .B(n_149), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_248), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_191), .B(n_174), .Y(n_288) );
NAND3xp33_ASAP7_75t_L g289 ( .A(n_187), .B(n_146), .C(n_179), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_234), .B(n_156), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_249), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_182), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_201), .B(n_143), .Y(n_293) );
AND2x6_ASAP7_75t_L g294 ( .A(n_183), .B(n_148), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_209), .B(n_211), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_212), .B(n_180), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_190), .B(n_184), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_185), .B(n_143), .Y(n_298) );
INVx4_ASAP7_75t_L g299 ( .A(n_204), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_214), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_200), .B(n_145), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_191), .B(n_145), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_189), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_206), .A2(n_160), .B1(n_178), .B2(n_180), .Y(n_304) );
NOR2xp67_ASAP7_75t_L g305 ( .A(n_208), .B(n_158), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_217), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_230), .B(n_180), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_232), .B(n_160), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_223), .A2(n_172), .B1(n_162), .B2(n_181), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_194), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_226), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_195), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_235), .B(n_155), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_206), .B(n_142), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_208), .B(n_142), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_199), .B(n_203), .Y(n_316) );
AND2x6_ASAP7_75t_SL g317 ( .A(n_205), .B(n_22), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_240), .B(n_155), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_204), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_237), .A2(n_175), .B1(n_156), .B2(n_158), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_240), .B(n_155), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_242), .B(n_155), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_242), .B(n_162), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_195), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_237), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_255), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_266), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_294), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_266), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_297), .A2(n_188), .B1(n_224), .B2(n_246), .Y(n_330) );
NAND2x1p5_ASAP7_75t_L g331 ( .A(n_270), .B(n_204), .Y(n_331) );
NAND3xp33_ASAP7_75t_L g332 ( .A(n_320), .B(n_219), .C(n_210), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_273), .A2(n_224), .B1(n_219), .B2(n_188), .Y(n_333) );
INVx4_ASAP7_75t_L g334 ( .A(n_270), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_290), .A2(n_222), .B(n_245), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_253), .B(n_181), .Y(n_336) );
NOR2x1_ASAP7_75t_L g337 ( .A(n_289), .B(n_162), .Y(n_337) );
INVx5_ASAP7_75t_L g338 ( .A(n_294), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_299), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_253), .B(n_246), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_262), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_281), .A2(n_246), .B1(n_222), .B2(n_245), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_259), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_271), .Y(n_344) );
BUFx10_ASAP7_75t_L g345 ( .A(n_288), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_310), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_296), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_259), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_290), .A2(n_222), .B(n_245), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_296), .Y(n_350) );
OR2x6_ASAP7_75t_L g351 ( .A(n_278), .B(n_250), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_256), .B(n_189), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_253), .B(n_181), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_251), .B(n_175), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_252), .Y(n_355) );
NAND2x1p5_ASAP7_75t_L g356 ( .A(n_267), .B(n_197), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_252), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_252), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_278), .A2(n_250), .B1(n_234), .B2(n_210), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_301), .A2(n_250), .B(n_234), .Y(n_360) );
BUFx2_ASAP7_75t_R g361 ( .A(n_303), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_259), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_251), .B(n_181), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_251), .B(n_196), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_294), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_307), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_288), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_281), .A2(n_175), .B1(n_156), .B2(n_158), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_288), .Y(n_369) );
NOR2xp67_ASAP7_75t_SL g370 ( .A(n_259), .B(n_186), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_310), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_265), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_277), .B(n_175), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_277), .Y(n_374) );
INVx6_ASAP7_75t_L g375 ( .A(n_285), .Y(n_375) );
INVx4_ASAP7_75t_SL g376 ( .A(n_294), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_261), .B(n_197), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_295), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_281), .B(n_175), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_277), .A2(n_162), .B1(n_172), .B2(n_194), .Y(n_380) );
BUFx3_ASAP7_75t_L g381 ( .A(n_285), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_268), .A2(n_225), .B1(n_172), .B2(n_139), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_260), .B(n_158), .Y(n_383) );
INVx1_ASAP7_75t_SL g384 ( .A(n_303), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_376), .B(n_254), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_338), .B(n_365), .Y(n_386) );
INVx6_ASAP7_75t_L g387 ( .A(n_345), .Y(n_387) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_373), .A2(n_314), .B(n_315), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_333), .A2(n_281), .B1(n_325), .B2(n_274), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_366), .A2(n_304), .B1(n_272), .B2(n_279), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_345), .Y(n_391) );
OR2x6_ASAP7_75t_L g392 ( .A(n_375), .B(n_267), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_378), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_335), .A2(n_259), .B(n_298), .Y(n_394) );
CKINVDCx11_ASAP7_75t_R g395 ( .A(n_341), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_347), .A2(n_282), .B1(n_276), .B2(n_275), .C(n_309), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_372), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_372), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_374), .A2(n_280), .B1(n_293), .B2(n_286), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_343), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_340), .A2(n_292), .B1(n_300), .B2(n_306), .Y(n_401) );
AOI21xp33_ASAP7_75t_L g402 ( .A1(n_352), .A2(n_264), .B(n_332), .Y(n_402) );
OR2x6_ASAP7_75t_L g403 ( .A(n_375), .B(n_267), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_330), .A2(n_305), .B1(n_294), .B2(n_285), .Y(n_404) );
BUFx8_ASAP7_75t_L g405 ( .A(n_381), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_345), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_327), .Y(n_407) );
OAI222xp33_ASAP7_75t_L g408 ( .A1(n_342), .A2(n_258), .B1(n_314), .B2(n_315), .C1(n_317), .C2(n_292), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_327), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_329), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_352), .A2(n_258), .B1(n_302), .B2(n_269), .Y(n_411) );
AOI222xp33_ASAP7_75t_L g412 ( .A1(n_350), .A2(n_295), .B1(n_306), .B2(n_311), .C1(n_300), .C2(n_315), .Y(n_412) );
INVx4_ASAP7_75t_L g413 ( .A(n_376), .Y(n_413) );
BUFx12f_ASAP7_75t_L g414 ( .A(n_375), .Y(n_414) );
BUFx10_ASAP7_75t_L g415 ( .A(n_375), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_329), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_326), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_336), .Y(n_418) );
O2A1O1Ixp33_ASAP7_75t_L g419 ( .A1(n_363), .A2(n_311), .B(n_172), .C(n_265), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_344), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_376), .B(n_269), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_385), .B(n_376), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_402), .A2(n_340), .B1(n_381), .B2(n_314), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_397), .B(n_383), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_393), .A2(n_384), .B1(n_353), .B2(n_380), .C(n_354), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_417), .A2(n_379), .B1(n_338), .B2(n_351), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_397), .B(n_379), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_389), .A2(n_351), .B1(n_383), .B2(n_354), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_395), .A2(n_351), .B1(n_337), .B2(n_369), .Y(n_429) );
NAND2x1_ASAP7_75t_L g430 ( .A(n_413), .B(n_343), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_399), .A2(n_382), .B1(n_368), .B2(n_365), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g432 ( .A1(n_405), .A2(n_338), .B1(n_373), .B2(n_328), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_398), .B(n_367), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_398), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_420), .B(n_355), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_396), .A2(n_377), .B1(n_364), .B2(n_359), .C(n_351), .Y(n_436) );
INVx8_ASAP7_75t_L g437 ( .A(n_414), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_395), .A2(n_294), .B1(n_358), .B2(n_357), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g439 ( .A1(n_390), .A2(n_349), .B(n_360), .Y(n_439) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_408), .A2(n_291), .B1(n_283), .B2(n_357), .C1(n_323), .C2(n_139), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_L g441 ( .A1(n_419), .A2(n_316), .B(n_339), .C(n_328), .Y(n_441) );
OAI211xp5_ASAP7_75t_L g442 ( .A1(n_404), .A2(n_313), .B(n_158), .C(n_339), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g443 ( .A1(n_401), .A2(n_291), .B1(n_283), .B2(n_339), .C(n_308), .Y(n_443) );
A2O1A1Ixp33_ASAP7_75t_L g444 ( .A1(n_418), .A2(n_338), .B(n_269), .C(n_284), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_405), .A2(n_338), .B1(n_139), .B2(n_371), .Y(n_445) );
CKINVDCx11_ASAP7_75t_R g446 ( .A(n_414), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_412), .A2(n_346), .B1(n_371), .B2(n_334), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_388), .A2(n_346), .B1(n_334), .B2(n_343), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_405), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_407), .Y(n_450) );
OAI211xp5_ASAP7_75t_SL g451 ( .A1(n_420), .A2(n_147), .B(n_141), .C(n_154), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_407), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_440), .B(n_138), .C(n_141), .Y(n_453) );
AOI22xp33_ASAP7_75t_SL g454 ( .A1(n_437), .A2(n_449), .B1(n_422), .B2(n_436), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_434), .B(n_409), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_423), .A2(n_391), .B1(n_406), .B2(n_403), .C(n_392), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_428), .A2(n_411), .B1(n_385), .B2(n_403), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_422), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_446), .Y(n_459) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_430), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_440), .B(n_138), .C(n_141), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g462 ( .A1(n_425), .A2(n_406), .B1(n_391), .B2(n_392), .C(n_403), .Y(n_462) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_439), .B(n_394), .C(n_416), .Y(n_463) );
AOI33xp33_ASAP7_75t_L g464 ( .A1(n_429), .A2(n_138), .A3(n_141), .B1(n_154), .B2(n_147), .B3(n_157), .Y(n_464) );
OAI33xp33_ASAP7_75t_L g465 ( .A1(n_426), .A2(n_138), .A3(n_147), .B1(n_154), .B2(n_157), .B3(n_221), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_450), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_450), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_430), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_435), .A2(n_424), .B1(n_439), .B2(n_443), .C(n_431), .Y(n_469) );
OAI222xp33_ASAP7_75t_L g470 ( .A1(n_432), .A2(n_413), .B1(n_392), .B2(n_403), .C1(n_386), .C2(n_385), .Y(n_470) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_441), .A2(n_416), .B(n_410), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_446), .A2(n_392), .B1(n_387), .B2(n_415), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_437), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_427), .A2(n_409), .B1(n_410), .B2(n_387), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_427), .A2(n_387), .B1(n_386), .B2(n_413), .Y(n_475) );
INVxp67_ASAP7_75t_SL g476 ( .A(n_452), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_434), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_447), .A2(n_387), .B1(n_386), .B2(n_361), .Y(n_478) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_448), .A2(n_318), .B(n_322), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_424), .Y(n_480) );
OAI211xp5_ASAP7_75t_SL g481 ( .A1(n_438), .A2(n_154), .B(n_157), .C(n_147), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_422), .Y(n_482) );
OR2x6_ASAP7_75t_L g483 ( .A(n_437), .B(n_400), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_437), .A2(n_415), .B1(n_139), .B2(n_421), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_433), .A2(n_157), .B1(n_321), .B2(n_287), .C(n_284), .Y(n_485) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_442), .A2(n_415), .B1(n_421), .B2(n_400), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_433), .B(n_400), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_451), .Y(n_488) );
NAND2xp33_ASAP7_75t_L g489 ( .A(n_444), .B(n_400), .Y(n_489) );
AOI33xp33_ASAP7_75t_L g490 ( .A1(n_454), .A2(n_445), .A3(n_221), .B1(n_22), .B2(n_23), .B3(n_287), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_477), .B(n_23), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_477), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_455), .B(n_400), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_466), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_460), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_466), .B(n_139), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_467), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_455), .B(n_27), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_467), .Y(n_499) );
AOI33xp33_ASAP7_75t_L g500 ( .A1(n_480), .A2(n_421), .A3(n_263), .B1(n_257), .B2(n_324), .B3(n_312), .Y(n_500) );
AOI221x1_ASAP7_75t_L g501 ( .A1(n_463), .A2(n_213), .B1(n_216), .B2(n_227), .C(n_228), .Y(n_501) );
INVx4_ASAP7_75t_L g502 ( .A(n_483), .Y(n_502) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_474), .Y(n_503) );
INVx3_ASAP7_75t_L g504 ( .A(n_460), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_480), .B(n_487), .Y(n_505) );
AOI211xp5_ASAP7_75t_L g506 ( .A1(n_478), .A2(n_213), .B(n_216), .C(n_227), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_469), .B(n_257), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_471), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_487), .B(n_29), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_471), .B(n_30), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_473), .B(n_334), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_471), .B(n_32), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_476), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_457), .A2(n_362), .B1(n_348), .B2(n_343), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_463), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_471), .B(n_479), .Y(n_516) );
AOI211xp5_ASAP7_75t_L g517 ( .A1(n_470), .A2(n_229), .B(n_216), .C(n_227), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_479), .B(n_35), .Y(n_518) );
INVxp67_ASAP7_75t_L g519 ( .A(n_479), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_460), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_458), .B(n_46), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g522 ( .A1(n_462), .A2(n_263), .B1(n_331), .B2(n_356), .C(n_227), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_486), .B(n_362), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_458), .B(n_362), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_458), .B(n_47), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_482), .B(n_49), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_460), .B(n_54), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_483), .Y(n_528) );
OAI31xp33_ASAP7_75t_L g529 ( .A1(n_456), .A2(n_331), .A3(n_356), .B(n_319), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_460), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_482), .B(n_348), .Y(n_531) );
OAI221xp5_ASAP7_75t_L g532 ( .A1(n_472), .A2(n_331), .B1(n_356), .B2(n_213), .C(n_216), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_468), .Y(n_533) );
OAI33xp33_ASAP7_75t_L g534 ( .A1(n_459), .A2(n_57), .A3(n_58), .B1(n_59), .B2(n_60), .B3(n_65), .Y(n_534) );
OAI221xp5_ASAP7_75t_L g535 ( .A1(n_488), .A2(n_213), .B1(n_228), .B2(n_229), .C(n_299), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_468), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_482), .B(n_66), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_468), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_468), .B(n_68), .Y(n_539) );
NOR2xp33_ASAP7_75t_R g540 ( .A(n_459), .B(n_468), .Y(n_540) );
NAND3xp33_ASAP7_75t_L g541 ( .A(n_464), .B(n_228), .C(n_229), .Y(n_541) );
INVxp67_ASAP7_75t_L g542 ( .A(n_513), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_505), .B(n_475), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_517), .A2(n_489), .B(n_465), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_505), .B(n_488), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_494), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_513), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_494), .B(n_483), .Y(n_548) );
OAI33xp33_ASAP7_75t_L g549 ( .A1(n_491), .A2(n_481), .A3(n_453), .B1(n_461), .B2(n_484), .B3(n_75), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_497), .B(n_483), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_492), .B(n_489), .Y(n_551) );
OR2x6_ASAP7_75t_L g552 ( .A(n_502), .B(n_362), .Y(n_552) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_541), .B(n_362), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_492), .B(n_485), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_516), .B(n_69), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_497), .B(n_72), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_516), .B(n_73), .Y(n_557) );
NOR3xp33_ASAP7_75t_L g558 ( .A(n_490), .B(n_231), .C(n_324), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_502), .B(n_74), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_495), .B(n_78), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_516), .B(n_79), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_493), .B(n_81), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_499), .B(n_83), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_499), .B(n_228), .Y(n_564) );
NAND3x2_ASAP7_75t_L g565 ( .A(n_518), .B(n_229), .C(n_186), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_493), .B(n_348), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_502), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_518), .B(n_231), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_503), .B(n_231), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_509), .Y(n_570) );
INVx4_ASAP7_75t_L g571 ( .A(n_502), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_509), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_528), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_518), .B(n_348), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_528), .Y(n_575) );
OAI322xp33_ASAP7_75t_L g576 ( .A1(n_519), .A2(n_312), .A3(n_299), .B1(n_348), .B2(n_343), .C1(n_319), .C2(n_186), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_503), .B(n_319), .Y(n_577) );
INVxp67_ASAP7_75t_L g578 ( .A(n_498), .Y(n_578) );
BUFx3_ASAP7_75t_L g579 ( .A(n_511), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_517), .A2(n_186), .B1(n_370), .B2(n_196), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_498), .B(n_370), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_520), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_530), .B(n_524), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_533), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_533), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_515), .B(n_530), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_536), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_495), .B(n_504), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_507), .B(n_500), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_536), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_507), .B(n_522), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_515), .B(n_538), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_522), .B(n_534), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_538), .B(n_519), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_536), .B(n_495), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_529), .B(n_540), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_495), .B(n_504), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_504), .B(n_508), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_508), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_529), .B(n_506), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_504), .B(n_508), .Y(n_601) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_542), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_599), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_547), .B(n_510), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_586), .B(n_510), .Y(n_605) );
OAI21xp33_ASAP7_75t_SL g606 ( .A1(n_600), .A2(n_523), .B(n_512), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_545), .B(n_512), .Y(n_607) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_579), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_586), .B(n_598), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_545), .B(n_512), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_598), .B(n_514), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_583), .B(n_514), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_594), .B(n_539), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_592), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_579), .B(n_537), .Y(n_615) );
AOI21xp33_ASAP7_75t_SL g616 ( .A1(n_596), .A2(n_532), .B(n_541), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_543), .B(n_506), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_594), .B(n_539), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_551), .B(n_595), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_551), .B(n_527), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_595), .B(n_527), .Y(n_621) );
NOR2xp67_ASAP7_75t_L g622 ( .A(n_571), .B(n_532), .Y(n_622) );
OAI22xp33_ASAP7_75t_SL g623 ( .A1(n_571), .A2(n_535), .B1(n_527), .B2(n_531), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_571), .B(n_527), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_591), .B(n_546), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_591), .B(n_526), .Y(n_626) );
AOI21xp33_ASAP7_75t_L g627 ( .A1(n_567), .A2(n_526), .B(n_537), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_546), .B(n_525), .Y(n_628) );
NOR2x1_ASAP7_75t_L g629 ( .A(n_553), .B(n_535), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_573), .B(n_575), .Y(n_630) );
OAI31xp33_ASAP7_75t_L g631 ( .A1(n_593), .A2(n_521), .A3(n_525), .B(n_496), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_593), .A2(n_534), .B1(n_521), .B2(n_496), .C(n_524), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_548), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_597), .B(n_531), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_597), .B(n_496), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_592), .Y(n_636) );
AOI21x1_ASAP7_75t_L g637 ( .A1(n_544), .A2(n_501), .B(n_589), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_550), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g639 ( .A(n_559), .B(n_501), .C(n_580), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_587), .B(n_590), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_587), .B(n_590), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_601), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_601), .B(n_582), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_584), .B(n_585), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_588), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_576), .A2(n_549), .B(n_552), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_588), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_588), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_578), .B(n_570), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_555), .B(n_561), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_555), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_557), .B(n_561), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_572), .B(n_557), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_559), .B(n_554), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_568), .B(n_577), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_608), .B(n_562), .Y(n_656) );
XNOR2xp5_ASAP7_75t_L g657 ( .A(n_650), .B(n_565), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_609), .B(n_574), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_625), .B(n_568), .Y(n_659) );
BUFx2_ASAP7_75t_L g660 ( .A(n_606), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_614), .B(n_569), .Y(n_661) );
NAND3xp33_ASAP7_75t_L g662 ( .A(n_616), .B(n_569), .C(n_562), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_609), .B(n_574), .Y(n_663) );
AOI211xp5_ASAP7_75t_L g664 ( .A1(n_606), .A2(n_581), .B(n_560), .C(n_558), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g665 ( .A(n_602), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_614), .B(n_566), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_644), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_642), .B(n_564), .Y(n_668) );
NAND3xp33_ASAP7_75t_SL g669 ( .A(n_646), .B(n_556), .C(n_563), .Y(n_669) );
AOI21x1_ASAP7_75t_SL g670 ( .A1(n_617), .A2(n_560), .B(n_552), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_644), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_636), .B(n_560), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_654), .A2(n_552), .B1(n_626), .B2(n_649), .Y(n_673) );
NOR2x1_ASAP7_75t_L g674 ( .A(n_622), .B(n_552), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_619), .B(n_634), .Y(n_675) );
INVx1_ASAP7_75t_SL g676 ( .A(n_633), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_633), .Y(n_677) );
INVx1_ASAP7_75t_SL g678 ( .A(n_643), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_636), .Y(n_679) );
INVx2_ASAP7_75t_SL g680 ( .A(n_647), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_643), .B(n_638), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_615), .A2(n_655), .B1(n_651), .B2(n_650), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_630), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_638), .B(n_642), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_642), .B(n_619), .Y(n_685) );
AND2x2_ASAP7_75t_SL g686 ( .A(n_652), .B(n_651), .Y(n_686) );
INVx3_ASAP7_75t_L g687 ( .A(n_603), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_616), .B(n_631), .C(n_632), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_611), .B(n_605), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_623), .B(n_622), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_652), .A2(n_653), .B1(n_611), .B2(n_635), .Y(n_691) );
XOR2x2_ASAP7_75t_L g692 ( .A(n_624), .B(n_623), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_640), .B(n_641), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_631), .A2(n_648), .B1(n_645), .B2(n_605), .C(n_610), .Y(n_694) );
AOI31xp33_ASAP7_75t_L g695 ( .A1(n_629), .A2(n_627), .A3(n_639), .B(n_647), .Y(n_695) );
OR2x2_ASAP7_75t_L g696 ( .A(n_612), .B(n_607), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_645), .B(n_635), .Y(n_697) );
XNOR2xp5_ASAP7_75t_L g698 ( .A(n_613), .B(n_618), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_604), .B(n_612), .Y(n_699) );
NOR2x1_ASAP7_75t_L g700 ( .A(n_629), .B(n_639), .Y(n_700) );
NOR2x1_ASAP7_75t_L g701 ( .A(n_628), .B(n_620), .Y(n_701) );
NOR3x1_ASAP7_75t_L g702 ( .A(n_637), .B(n_620), .C(n_621), .Y(n_702) );
XNOR2x1_ASAP7_75t_L g703 ( .A(n_621), .B(n_637), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_608), .B(n_654), .Y(n_704) );
NOR3x1_ASAP7_75t_L g705 ( .A(n_626), .B(n_596), .C(n_625), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_644), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_614), .B(n_636), .Y(n_707) );
XOR2x2_ASAP7_75t_L g708 ( .A(n_608), .B(n_449), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_644), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_608), .B(n_654), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_654), .A2(n_625), .B1(n_649), .B2(n_606), .C(n_602), .Y(n_711) );
OAI21xp5_ASAP7_75t_L g712 ( .A1(n_700), .A2(n_660), .B(n_688), .Y(n_712) );
OA22x2_ASAP7_75t_L g713 ( .A1(n_660), .A2(n_690), .B1(n_665), .B2(n_677), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_665), .B(n_704), .Y(n_714) );
OAI221xp5_ASAP7_75t_L g715 ( .A1(n_711), .A2(n_695), .B1(n_692), .B2(n_673), .C(n_703), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_669), .A2(n_694), .B1(n_710), .B2(n_686), .Y(n_716) );
AOI211xp5_ASAP7_75t_L g717 ( .A1(n_664), .A2(n_662), .B(n_657), .C(n_656), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_708), .Y(n_718) );
NOR2x1_ASAP7_75t_SL g719 ( .A(n_680), .B(n_675), .Y(n_719) );
BUFx2_ASAP7_75t_L g720 ( .A(n_677), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_702), .B(n_686), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_674), .A2(n_657), .B(n_707), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_699), .A2(n_659), .B1(n_701), .B2(n_696), .Y(n_723) );
OA22x2_ASAP7_75t_L g724 ( .A1(n_691), .A2(n_682), .B1(n_698), .B2(n_676), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_683), .A2(n_667), .B1(n_706), .B2(n_671), .C(n_709), .Y(n_725) );
NAND5xp2_ASAP7_75t_L g726 ( .A(n_670), .B(n_672), .C(n_705), .D(n_661), .E(n_689), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_687), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_724), .A2(n_680), .B1(n_679), .B2(n_707), .Y(n_728) );
INVx1_ASAP7_75t_SL g729 ( .A(n_720), .Y(n_729) );
XNOR2xp5_ASAP7_75t_L g730 ( .A(n_717), .B(n_678), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g731 ( .A(n_713), .B(n_687), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_715), .A2(n_689), .B1(n_666), .B2(n_684), .Y(n_732) );
OAI21xp33_ASAP7_75t_L g733 ( .A1(n_713), .A2(n_697), .B(n_681), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_717), .A2(n_697), .B1(n_663), .B2(n_658), .Y(n_734) );
XOR2xp5_ASAP7_75t_L g735 ( .A(n_718), .B(n_668), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_725), .B(n_675), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_729), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_735), .B(n_714), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_736), .B(n_712), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g740 ( .A1(n_728), .A2(n_712), .B(n_722), .C(n_721), .Y(n_740) );
NAND3x1_ASAP7_75t_L g741 ( .A(n_732), .B(n_716), .C(n_719), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_737), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_739), .B(n_730), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_741), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_742), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_743), .A2(n_738), .B(n_740), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_746), .B(n_744), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_745), .Y(n_748) );
AOI222xp33_ASAP7_75t_SL g749 ( .A1(n_748), .A2(n_744), .B1(n_726), .B2(n_733), .C1(n_731), .C2(n_734), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_747), .Y(n_750) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_750), .A2(n_727), .B1(n_685), .B2(n_693), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_751), .A2(n_749), .B(n_723), .Y(n_752) );
endmodule