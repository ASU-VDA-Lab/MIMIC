module fake_jpeg_15577_n_200 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_200);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

OR2x2_ASAP7_75t_L g13 ( 
.A(n_12),
.B(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_17),
.B1(n_18),
.B2(n_26),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_20),
.B1(n_17),
.B2(n_26),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_17),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_28),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_20),
.B1(n_26),
.B2(n_16),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_20),
.B1(n_36),
.B2(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_14),
.B1(n_15),
.B2(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_28),
.A2(n_22),
.B1(n_15),
.B2(n_23),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_30),
.B(n_22),
.Y(n_84)
);

AOI22x1_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_41),
.B1(n_43),
.B2(n_32),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_41),
.B1(n_38),
.B2(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_13),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_65),
.Y(n_77)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_68),
.Y(n_81)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_13),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_35),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_35),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_72),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_99)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_48),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_75),
.B(n_78),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_48),
.B(n_37),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_58),
.B1(n_59),
.B2(n_57),
.Y(n_89)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_43),
.B1(n_32),
.B2(n_40),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_0),
.Y(n_83)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_59),
.C(n_54),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_68),
.B(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_41),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_112)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_77),
.B(n_71),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_93),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_67),
.Y(n_92)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_101),
.B(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_54),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_91),
.B(n_101),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_63),
.B(n_15),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_85),
.B(n_82),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_40),
.B1(n_25),
.B2(n_21),
.Y(n_100)
);

OA21x2_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_40),
.B(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_19),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_117),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_101),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_95),
.B(n_96),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_94),
.B(n_92),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_77),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_94),
.C(n_100),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_118),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_114),
.B(n_115),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_73),
.B1(n_85),
.B2(n_82),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_119),
.B1(n_88),
.B2(n_103),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_92),
.B(n_25),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_87),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_76),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_19),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_133),
.Y(n_147)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_123),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_128),
.B1(n_106),
.B2(n_112),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_132),
.C(n_135),
.Y(n_142)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_19),
.B(n_1),
.C(n_3),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_89),
.C(n_99),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_80),
.B1(n_24),
.B2(n_21),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_72),
.C(n_80),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_19),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_105),
.C(n_115),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_134),
.C(n_128),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_116),
.B(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_150),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_149),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_133),
.B(n_19),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_132),
.C(n_124),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_130),
.C(n_125),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_154),
.C(n_161),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_130),
.C(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_163),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_123),
.C(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_0),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_147),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_172),
.C(n_160),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_156),
.A2(n_145),
.B(n_137),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_158),
.B(n_4),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_141),
.B1(n_143),
.B2(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_162),
.B(n_12),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_171),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_141),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_141),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_168),
.A2(n_155),
.B(n_160),
.C(n_159),
.Y(n_174)
);

OAI22x1_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_179),
.B1(n_180),
.B2(n_1),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_153),
.B(n_161),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_176),
.C(n_169),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_163),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_178),
.B(n_6),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_158),
.B1(n_4),
.B2(n_5),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_165),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_182),
.B(n_183),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_181),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_164),
.C(n_19),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_186),
.B(n_187),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_52),
.B(n_10),
.Y(n_193)
);

OAI21x1_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_190),
.B(n_9),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_186),
.A2(n_8),
.B(n_9),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_193),
.B(n_195),
.Y(n_196)
);

AOI31xp67_ASAP7_75t_SL g197 ( 
.A1(n_194),
.A2(n_190),
.A3(n_192),
.B(n_10),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_10),
.B(n_11),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_196),
.C(n_11),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_11),
.Y(n_200)
);


endmodule