module fake_ariane_1424_n_162 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_41, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_40, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_162);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_41;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_162;

wire n_83;
wire n_56;
wire n_60;
wire n_160;
wire n_64;
wire n_124;
wire n_119;
wire n_90;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_158;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_152;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_43;
wire n_81;
wire n_87;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_54;

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

INVxp33_ASAP7_75t_SL g54 ( 
.A(n_29),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVxp33_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_1),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_21),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_0),
.Y(n_71)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_1),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_2),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_3),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_57),
.B(n_6),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_23),
.Y(n_88)
);

AO21x2_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_26),
.B(n_30),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_31),
.B1(n_39),
.B2(n_40),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_64),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_56),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_53),
.B(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_55),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_66),
.C(n_57),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_66),
.B(n_61),
.Y(n_103)
);

NOR2xp67_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_104),
.B(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_88),
.B(n_90),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_71),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_75),
.B(n_88),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_81),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_SL g115 ( 
.A1(n_103),
.A2(n_90),
.B(n_87),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_89),
.B(n_87),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_76),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_84),
.B1(n_75),
.B2(n_76),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_80),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

AO21x2_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_89),
.B(n_98),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

OAI21x1_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_81),
.B(n_77),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_119),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_112),
.B(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_108),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_121),
.B(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_108),
.Y(n_138)
);

OAI221xp5_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_108),
.B1(n_107),
.B2(n_105),
.C(n_81),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_107),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_107),
.B(n_130),
.Y(n_141)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_126),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_126),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_107),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_135),
.B1(n_138),
.B2(n_127),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_144),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_146),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_148),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_143),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_151),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_145),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_157)
);

AND2x4_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_155),
.Y(n_158)
);

NOR5xp2_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_139),
.C(n_125),
.D(n_147),
.E(n_128),
.Y(n_159)
);

OAI21x1_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_158),
.B(n_136),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_139),
.B(n_125),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_160),
.B1(n_125),
.B2(n_127),
.Y(n_162)
);


endmodule