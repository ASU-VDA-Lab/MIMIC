module fake_jpeg_19233_n_174 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_6),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_38),
.Y(n_52)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_18),
.B1(n_22),
.B2(n_26),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_47),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_46),
.B1(n_33),
.B2(n_35),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_16),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_49),
.C(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_26),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_37),
.B1(n_39),
.B2(n_32),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_32),
.B(n_37),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_57),
.B(n_71),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_65),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_64),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_35),
.B1(n_38),
.B2(n_33),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_72),
.B1(n_46),
.B2(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_28),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_17),
.Y(n_85)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_55),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

AOI32xp33_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_51),
.A3(n_43),
.B1(n_50),
.B2(n_23),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_81),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_75),
.A2(n_50),
.B1(n_55),
.B2(n_40),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_29),
.B(n_17),
.C(n_2),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_63),
.A3(n_72),
.B1(n_66),
.B2(n_3),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_40),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_95),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_55),
.B1(n_30),
.B2(n_27),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_8),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_30),
.C(n_27),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_65),
.C(n_68),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_106),
.C(n_80),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_67),
.B(n_64),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_107),
.B(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_103),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_109),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_58),
.C(n_56),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_56),
.B(n_1),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_15),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_10),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_15),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_113),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_77),
.B1(n_82),
.B2(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_120),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_86),
.B1(n_92),
.B2(n_96),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_124),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_94),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_126),
.C(n_110),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_88),
.B1(n_84),
.B2(n_93),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_114),
.B1(n_107),
.B2(n_5),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_84),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_129),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_100),
.B(n_103),
.C(n_108),
.D(n_101),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_123),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_99),
.C(n_110),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_129),
.C(n_120),
.Y(n_145)
);

AO221x1_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.C(n_5),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_141),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_121),
.B1(n_127),
.B2(n_5),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_145),
.C(n_148),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_130),
.B(n_123),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_146),
.A2(n_134),
.B(n_132),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_140),
.A2(n_122),
.B1(n_119),
.B2(n_116),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_7),
.Y(n_151)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_139),
.B1(n_140),
.B2(n_138),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_142),
.B1(n_132),
.B2(n_136),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_147),
.B(n_136),
.C(n_133),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_159),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_144),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_162),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_151),
.B1(n_11),
.B2(n_13),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_163),
.Y(n_168)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_170),
.B(n_14),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_160),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_166),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_167),
.A2(n_10),
.B(n_11),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_173),
.B(n_172),
.Y(n_174)
);


endmodule