module fake_jpeg_1465_n_21 (n_3, n_2, n_1, n_0, n_4, n_5, n_21);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_21;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_1),
.A2(n_2),
.B1(n_5),
.B2(n_4),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_1),
.Y(n_9)
);

AOI22xp33_ASAP7_75t_SL g10 ( 
.A1(n_0),
.A2(n_5),
.B1(n_3),
.B2(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_6),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g12 ( 
.A1(n_7),
.A2(n_0),
.B1(n_2),
.B2(n_9),
.Y(n_12)
);

A2O1A1Ixp33_ASAP7_75t_SL g17 ( 
.A1(n_12),
.A2(n_14),
.B(n_7),
.C(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_13),
.B(n_8),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_10),
.A2(n_0),
.B1(n_9),
.B2(n_6),
.Y(n_14)
);

AOI21x1_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_16),
.B(n_17),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_12),
.B(n_14),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_19),
.C(n_11),
.Y(n_21)
);


endmodule