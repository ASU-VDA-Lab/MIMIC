module real_aes_885_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_782, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_782;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g241 ( .A(n_0), .B(n_178), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_1), .B(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_2), .B(n_154), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_3), .B(n_176), .Y(n_491) );
INVx1_ASAP7_75t_L g150 ( .A(n_4), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_5), .B(n_154), .Y(n_199) );
NAND2xp33_ASAP7_75t_SL g261 ( .A(n_6), .B(n_160), .Y(n_261) );
INVx1_ASAP7_75t_L g253 ( .A(n_7), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_8), .A2(n_58), .B1(n_771), .B2(n_772), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_8), .Y(n_771) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_9), .Y(n_111) );
AND2x2_ASAP7_75t_L g197 ( .A(n_10), .B(n_183), .Y(n_197) );
AND2x2_ASAP7_75t_L g484 ( .A(n_11), .B(n_259), .Y(n_484) );
AND2x2_ASAP7_75t_L g493 ( .A(n_12), .B(n_140), .Y(n_493) );
INVx2_ASAP7_75t_L g142 ( .A(n_13), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_14), .B(n_176), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_15), .Y(n_113) );
AOI221x1_ASAP7_75t_L g256 ( .A1(n_16), .A2(n_162), .B1(n_257), .B2(n_259), .C(n_260), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_17), .B(n_154), .Y(n_221) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_18), .A2(n_70), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_18), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_19), .B(n_154), .Y(n_533) );
NOR2xp33_ASAP7_75t_SL g107 ( .A(n_20), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g131 ( .A(n_20), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_21), .A2(n_769), .B1(n_773), .B2(n_774), .Y(n_768) );
INVx1_ASAP7_75t_L g773 ( .A(n_21), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_22), .A2(n_92), .B1(n_145), .B2(n_154), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_23), .A2(n_162), .B(n_201), .Y(n_200) );
AOI221xp5_ASAP7_75t_SL g230 ( .A1(n_24), .A2(n_37), .B1(n_154), .B2(n_162), .C(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_25), .B(n_178), .Y(n_202) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_26), .A2(n_91), .B(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g184 ( .A(n_26), .B(n_91), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_27), .B(n_176), .Y(n_225) );
INVxp67_ASAP7_75t_L g255 ( .A(n_28), .Y(n_255) );
AND2x2_ASAP7_75t_L g194 ( .A(n_29), .B(n_182), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_30), .A2(n_162), .B(n_240), .Y(n_239) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_31), .A2(n_259), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_32), .B(n_176), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_33), .A2(n_162), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_34), .B(n_176), .Y(n_547) );
AND2x2_ASAP7_75t_L g152 ( .A(n_35), .B(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g160 ( .A(n_35), .B(n_150), .Y(n_160) );
INVx1_ASAP7_75t_L g166 ( .A(n_35), .Y(n_166) );
NOR3xp33_ASAP7_75t_L g109 ( .A(n_36), .B(n_110), .C(n_112), .Y(n_109) );
OR2x6_ASAP7_75t_L g129 ( .A(n_36), .B(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_38), .B(n_154), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g161 ( .A1(n_39), .A2(n_82), .B1(n_162), .B2(n_164), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_40), .B(n_176), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_41), .B(n_154), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_42), .B(n_178), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_43), .A2(n_162), .B(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g244 ( .A(n_44), .B(n_182), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_45), .B(n_178), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_46), .B(n_182), .Y(n_234) );
AOI22xp5_ASAP7_75t_SL g120 ( .A1(n_47), .A2(n_121), .B1(n_122), .B2(n_123), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_47), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_48), .B(n_154), .Y(n_515) );
INVx1_ASAP7_75t_L g148 ( .A(n_49), .Y(n_148) );
INVx1_ASAP7_75t_L g157 ( .A(n_49), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_50), .B(n_176), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_51), .Y(n_779) );
AND2x2_ASAP7_75t_L g523 ( .A(n_52), .B(n_182), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_53), .B(n_154), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_54), .B(n_178), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_55), .B(n_178), .Y(n_546) );
AND2x2_ASAP7_75t_L g185 ( .A(n_56), .B(n_182), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_57), .B(n_154), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_58), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_59), .B(n_176), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_60), .B(n_154), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_61), .A2(n_162), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_62), .B(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_SL g226 ( .A(n_63), .B(n_183), .Y(n_226) );
AND2x2_ASAP7_75t_L g539 ( .A(n_64), .B(n_183), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_65), .A2(n_162), .B(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_66), .B(n_176), .Y(n_203) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_67), .B(n_140), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_68), .B(n_178), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_69), .B(n_178), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_70), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_71), .A2(n_94), .B1(n_162), .B2(n_164), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_72), .B(n_176), .Y(n_536) );
INVx1_ASAP7_75t_L g153 ( .A(n_73), .Y(n_153) );
INVx1_ASAP7_75t_L g159 ( .A(n_73), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_74), .B(n_178), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_75), .A2(n_162), .B(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_76), .A2(n_162), .B(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_77), .A2(n_162), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g549 ( .A(n_78), .B(n_183), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_79), .B(n_182), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_80), .A2(n_85), .B1(n_145), .B2(n_154), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_81), .B(n_154), .Y(n_180) );
INVx1_ASAP7_75t_L g108 ( .A(n_83), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_84), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_86), .B(n_178), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_87), .B(n_178), .Y(n_233) );
AND2x2_ASAP7_75t_L g505 ( .A(n_88), .B(n_140), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_89), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_90), .A2(n_162), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_93), .B(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_95), .A2(n_162), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_96), .B(n_176), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_97), .B(n_154), .Y(n_243) );
INVxp67_ASAP7_75t_L g258 ( .A(n_98), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_99), .B(n_176), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_100), .A2(n_162), .B(n_223), .Y(n_222) );
BUFx2_ASAP7_75t_L g538 ( .A(n_101), .Y(n_538) );
BUFx2_ASAP7_75t_L g117 ( .A(n_102), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_114), .B(n_778), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g780 ( .A(n_105), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
AND2x4_ASAP7_75t_SL g106 ( .A(n_107), .B(n_109), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_108), .B(n_131), .Y(n_130) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
AND2x6_ASAP7_75t_SL g128 ( .A(n_113), .B(n_129), .Y(n_128) );
OR2x6_ASAP7_75t_SL g756 ( .A(n_113), .B(n_757), .Y(n_756) );
OR2x2_ASAP7_75t_L g760 ( .A(n_113), .B(n_129), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_113), .B(n_757), .Y(n_767) );
AO221x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_118), .B1(n_765), .B2(n_768), .C(n_775), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
NOR2x1_ASAP7_75t_R g765 ( .A(n_117), .B(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_761), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_126), .B(n_758), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_120), .Y(n_762) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_132), .B1(n_461), .B2(n_754), .Y(n_126) );
INVx3_ASAP7_75t_SL g764 ( .A(n_127), .Y(n_764) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g757 ( .A(n_129), .Y(n_757) );
AO22x1_ASAP7_75t_L g763 ( .A1(n_132), .A2(n_461), .B1(n_755), .B2(n_764), .Y(n_763) );
XNOR2x1_ASAP7_75t_L g769 ( .A(n_132), .B(n_770), .Y(n_769) );
AND3x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_332), .C(n_406), .Y(n_132) );
NOR3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_274), .C(n_305), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_207), .B(n_216), .C(n_245), .Y(n_134) );
AOI21x1_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_186), .B(n_205), .Y(n_135) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_136), .A2(n_308), .B1(n_314), .B2(n_317), .Y(n_307) );
AND2x2_ASAP7_75t_L g441 ( .A(n_136), .B(n_209), .Y(n_441) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_170), .Y(n_136) );
BUFx2_ASAP7_75t_L g212 ( .A(n_137), .Y(n_212) );
AND2x2_ASAP7_75t_L g300 ( .A(n_137), .B(n_171), .Y(n_300) );
AND2x2_ASAP7_75t_L g371 ( .A(n_137), .B(n_215), .Y(n_371) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_138), .Y(n_265) );
AOI21x1_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_143), .B(n_169), .Y(n_138) );
INVx2_ASAP7_75t_SL g139 ( .A(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_140), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_140), .A2(n_533), .B(n_534), .Y(n_532) );
BUFx4f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx3_ASAP7_75t_L g237 ( .A(n_141), .Y(n_237) );
AND2x2_ASAP7_75t_SL g183 ( .A(n_142), .B(n_184), .Y(n_183) );
AND2x4_ASAP7_75t_L g204 ( .A(n_142), .B(n_184), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_161), .Y(n_143) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_145), .A2(n_164), .B1(n_252), .B2(n_254), .Y(n_251) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_151), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g163 ( .A(n_148), .B(n_150), .Y(n_163) );
AND2x4_ASAP7_75t_L g176 ( .A(n_148), .B(n_158), .Y(n_176) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x6_ASAP7_75t_L g162 ( .A(n_152), .B(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g168 ( .A(n_153), .Y(n_168) );
AND2x6_ASAP7_75t_L g178 ( .A(n_153), .B(n_156), .Y(n_178) );
AND2x4_ASAP7_75t_L g154 ( .A(n_155), .B(n_160), .Y(n_154) );
INVx1_ASAP7_75t_L g262 ( .A(n_155), .Y(n_262) );
AND2x4_ASAP7_75t_L g155 ( .A(n_156), .B(n_158), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx5_ASAP7_75t_L g179 ( .A(n_160), .Y(n_179) );
AND2x4_ASAP7_75t_L g164 ( .A(n_163), .B(n_165), .Y(n_164) );
NOR2x1p5_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g264 ( .A(n_170), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g206 ( .A(n_171), .B(n_196), .Y(n_206) );
OR2x2_ASAP7_75t_L g214 ( .A(n_171), .B(n_215), .Y(n_214) );
AND2x4_ASAP7_75t_L g269 ( .A(n_171), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g316 ( .A(n_171), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_171), .B(n_215), .Y(n_324) );
AND2x2_ASAP7_75t_L g361 ( .A(n_171), .B(n_265), .Y(n_361) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_171), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_171), .B(n_195), .Y(n_402) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_181), .B(n_185), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_180), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_177), .B(n_179), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_178), .B(n_538), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_179), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_179), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_179), .A2(n_224), .B(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_179), .A2(n_232), .B(n_233), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_179), .A2(n_241), .B(n_242), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_179), .A2(n_481), .B(n_482), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_179), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_179), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_179), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_179), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_179), .A2(n_536), .B(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_179), .A2(n_546), .B(n_547), .Y(n_545) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_181), .A2(n_188), .B(n_194), .Y(n_187) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_181), .A2(n_188), .B(n_194), .Y(n_215) );
AOI21x1_ASAP7_75t_L g486 ( .A1(n_181), .A2(n_487), .B(n_493), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_182), .A2(n_230), .B(n_234), .Y(n_229) );
AO21x2_ASAP7_75t_L g471 ( .A1(n_182), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_182), .A2(n_500), .B(n_501), .Y(n_499) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g303 ( .A(n_186), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_186), .B(n_264), .Y(n_359) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_186), .Y(n_460) );
AND2x4_ASAP7_75t_L g186 ( .A(n_187), .B(n_195), .Y(n_186) );
AND2x2_ASAP7_75t_L g205 ( .A(n_187), .B(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g285 ( .A(n_187), .B(n_196), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_187), .B(n_316), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_193), .Y(n_188) );
AND2x2_ASAP7_75t_L g352 ( .A(n_195), .B(n_269), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_195), .B(n_264), .Y(n_408) );
INVx5_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g210 ( .A(n_196), .Y(n_210) );
AND2x2_ASAP7_75t_L g279 ( .A(n_196), .B(n_270), .Y(n_279) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_196), .Y(n_299) );
AND2x4_ASAP7_75t_L g306 ( .A(n_196), .B(n_215), .Y(n_306) );
AND2x2_ASAP7_75t_SL g453 ( .A(n_196), .B(n_265), .Y(n_453) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_204), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_204), .B(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_204), .B(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_204), .B(n_258), .Y(n_257) );
NOR3xp33_ASAP7_75t_L g260 ( .A(n_204), .B(n_261), .C(n_262), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_204), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_204), .A2(n_525), .B(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g432 ( .A(n_205), .Y(n_432) );
INVx1_ASAP7_75t_L g374 ( .A(n_206), .Y(n_374) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_211), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g296 ( .A(n_210), .B(n_214), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_210), .B(n_265), .Y(n_389) );
AND2x2_ASAP7_75t_L g391 ( .A(n_210), .B(n_213), .Y(n_391) );
AOI32xp33_ASAP7_75t_L g457 ( .A1(n_210), .A2(n_273), .A3(n_428), .B1(n_458), .B2(n_460), .Y(n_457) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
AND2x2_ASAP7_75t_L g283 ( .A(n_212), .B(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g401 ( .A(n_212), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g424 ( .A(n_212), .B(n_285), .Y(n_424) );
AND2x2_ASAP7_75t_L g451 ( .A(n_212), .B(n_352), .Y(n_451) );
AND2x2_ASAP7_75t_L g377 ( .A(n_213), .B(n_265), .Y(n_377) );
AND2x2_ASAP7_75t_L g452 ( .A(n_213), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g270 ( .A(n_215), .Y(n_270) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_227), .Y(n_217) );
NOR2x1p5_ASAP7_75t_L g310 ( .A(n_218), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g328 ( .A(n_218), .Y(n_328) );
OR2x2_ASAP7_75t_L g356 ( .A(n_218), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x4_ASAP7_75t_SL g273 ( .A(n_219), .B(n_250), .Y(n_273) );
AND2x4_ASAP7_75t_L g289 ( .A(n_219), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g292 ( .A(n_219), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g320 ( .A(n_219), .B(n_229), .Y(n_320) );
OR2x2_ASAP7_75t_L g345 ( .A(n_219), .B(n_294), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_219), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_219), .B(n_229), .Y(n_380) );
INVx2_ASAP7_75t_L g396 ( .A(n_219), .Y(n_396) );
AND2x2_ASAP7_75t_L g411 ( .A(n_219), .B(n_249), .Y(n_411) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_219), .Y(n_435) );
INVx1_ASAP7_75t_L g440 ( .A(n_219), .Y(n_440) );
OR2x6_ASAP7_75t_L g219 ( .A(n_220), .B(n_226), .Y(n_219) );
AND2x2_ASAP7_75t_L g304 ( .A(n_227), .B(n_289), .Y(n_304) );
AND2x2_ASAP7_75t_L g325 ( .A(n_227), .B(n_273), .Y(n_325) );
INVx1_ASAP7_75t_L g357 ( .A(n_227), .Y(n_357) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_235), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g248 ( .A(n_229), .Y(n_248) );
INVx2_ASAP7_75t_L g294 ( .A(n_229), .Y(n_294) );
BUFx3_ASAP7_75t_L g311 ( .A(n_229), .Y(n_311) );
AND2x2_ASAP7_75t_L g350 ( .A(n_229), .B(n_235), .Y(n_350) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_229), .Y(n_448) );
INVx2_ASAP7_75t_L g263 ( .A(n_235), .Y(n_263) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_235), .Y(n_272) );
INVx1_ASAP7_75t_L g288 ( .A(n_235), .Y(n_288) );
OR2x2_ASAP7_75t_L g293 ( .A(n_235), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g313 ( .A(n_235), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_235), .B(n_290), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_235), .B(n_396), .Y(n_395) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AOI21x1_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_244), .Y(n_236) );
INVx4_ASAP7_75t_L g259 ( .A(n_237), .Y(n_259) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_237), .A2(n_478), .B(n_484), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_243), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_264), .B(n_266), .Y(n_245) );
AND2x2_ASAP7_75t_SL g246 ( .A(n_247), .B(n_249), .Y(n_246) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_247), .Y(n_456) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVxp67_ASAP7_75t_SL g282 ( .A(n_248), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_248), .B(n_288), .Y(n_330) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_248), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_249), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g335 ( .A(n_249), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g386 ( .A(n_249), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_249), .A2(n_391), .B1(n_392), .B2(n_397), .C(n_400), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_249), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g249 ( .A(n_250), .B(n_263), .Y(n_249) );
INVx3_ASAP7_75t_L g290 ( .A(n_250), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_250), .B(n_294), .Y(n_394) );
AND2x2_ASAP7_75t_L g423 ( .A(n_250), .B(n_396), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_250), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
INVx3_ASAP7_75t_L g542 ( .A(n_259), .Y(n_542) );
AND2x2_ASAP7_75t_L g331 ( .A(n_264), .B(n_306), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_264), .A2(n_284), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g268 ( .A(n_265), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g277 ( .A(n_265), .Y(n_277) );
OR2x2_ASAP7_75t_L g323 ( .A(n_265), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_265), .B(n_306), .Y(n_415) );
OR2x2_ASAP7_75t_L g447 ( .A(n_265), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g459 ( .A(n_265), .B(n_365), .Y(n_459) );
INVxp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
INVx2_ASAP7_75t_L g337 ( .A(n_268), .Y(n_337) );
INVx3_ASAP7_75t_SL g403 ( .A(n_269), .Y(n_403) );
INVxp67_ASAP7_75t_L g353 ( .A(n_271), .Y(n_353) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
AOI322xp5_ASAP7_75t_L g275 ( .A1(n_273), .A2(n_276), .A3(n_280), .B1(n_283), .B2(n_286), .C1(n_291), .C2(n_295), .Y(n_275) );
INVx1_ASAP7_75t_SL g364 ( .A(n_273), .Y(n_364) );
AND2x4_ASAP7_75t_L g449 ( .A(n_273), .B(n_336), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_297), .Y(n_274) );
NOR2x1_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OR2x2_ASAP7_75t_L g302 ( .A(n_277), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g398 ( .A(n_277), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g426 ( .A(n_277), .B(n_279), .Y(n_426) );
AOI32xp33_ASAP7_75t_L g427 ( .A1(n_277), .A2(n_278), .A3(n_428), .B1(n_430), .B2(n_433), .Y(n_427) );
OR2x2_ASAP7_75t_L g431 ( .A(n_277), .B(n_324), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g387 ( .A(n_278), .B(n_303), .C(n_388), .Y(n_387) );
OAI22xp33_ASAP7_75t_SL g407 ( .A1(n_278), .A2(n_344), .B1(n_408), .B2(n_409), .Y(n_407) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g410 ( .A(n_281), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_285), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
OAI322xp33_ASAP7_75t_L g333 ( .A1(n_289), .A2(n_293), .A3(n_302), .B1(n_334), .B2(n_337), .C1(n_338), .C2(n_339), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_289), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_289), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g312 ( .A(n_290), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g344 ( .A(n_290), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_290), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g405 ( .A(n_293), .Y(n_405) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_294), .Y(n_336) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_301), .B(n_304), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_300), .B(n_348), .Y(n_347) );
AOI322xp5_ASAP7_75t_SL g442 ( .A1(n_300), .A2(n_306), .A3(n_423), .B1(n_441), .B2(n_443), .C1(n_446), .C2(n_449), .Y(n_442) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI21xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B(n_321), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_306), .B(n_316), .Y(n_338) );
INVx2_ASAP7_75t_SL g348 ( .A(n_306), .Y(n_348) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_SL g373 ( .A(n_312), .Y(n_373) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_313), .Y(n_343) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g418 ( .A(n_319), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g372 ( .A(n_320), .B(n_373), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_325), .B1(n_326), .B2(n_331), .Y(n_321) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NOR4xp75_ASAP7_75t_L g332 ( .A(n_333), .B(n_346), .C(n_366), .D(n_382), .Y(n_332) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g340 ( .A(n_341), .B(n_344), .Y(n_340) );
INVxp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_344), .A2(n_421), .B1(n_424), .B2(n_425), .Y(n_420) );
OR2x2_ASAP7_75t_L g385 ( .A(n_345), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g429 ( .A(n_345), .Y(n_429) );
OAI221xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B1(n_351), .B2(n_353), .C(n_354), .Y(n_346) );
INVx2_ASAP7_75t_L g365 ( .A(n_350), .Y(n_365) );
AND2x2_ASAP7_75t_L g422 ( .A(n_350), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B1(n_360), .B2(n_362), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g417 ( .A(n_361), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_362), .A2(n_368), .B1(n_384), .B2(n_387), .Y(n_383) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
OAI221xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_372), .B1(n_374), .B2(n_375), .C(n_782), .Y(n_366) );
AND2x2_ASAP7_75t_SL g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g434 ( .A(n_373), .B(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g419 ( .A(n_381), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_390), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B(n_404), .Y(n_400) );
NOR3xp33_ASAP7_75t_SL g406 ( .A(n_407), .B(n_412), .C(n_436), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_427), .Y(n_412) );
O2A1O1Ixp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B(n_418), .C(n_420), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g428 ( .A(n_419), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
NAND4xp25_ASAP7_75t_SL g436 ( .A(n_437), .B(n_442), .C(n_450), .D(n_457), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
OAI21xp5_ASAP7_75t_SL g450 ( .A1(n_451), .A2(n_452), .B(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_679), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_615), .C(n_662), .Y(n_462) );
NAND4xp25_ASAP7_75t_SL g463 ( .A(n_464), .B(n_550), .C(n_568), .D(n_594), .Y(n_463) );
OAI21xp33_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_509), .B(n_510), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_466), .B(n_494), .Y(n_465) );
INVx1_ASAP7_75t_L g730 ( .A(n_466), .Y(n_730) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_474), .Y(n_466) );
INVx2_ASAP7_75t_L g554 ( .A(n_467), .Y(n_554) );
AND2x2_ASAP7_75t_L g574 ( .A(n_467), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g676 ( .A(n_467), .B(n_496), .Y(n_676) );
AND2x2_ASAP7_75t_L g736 ( .A(n_467), .B(n_555), .Y(n_736) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_468), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g620 ( .A(n_469), .B(n_477), .Y(n_620) );
BUFx3_ASAP7_75t_L g630 ( .A(n_469), .Y(n_630) );
AND2x2_ASAP7_75t_L g693 ( .A(n_469), .B(n_694), .Y(n_693) );
AND2x4_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
AND2x4_ASAP7_75t_L g508 ( .A(n_470), .B(n_471), .Y(n_508) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g739 ( .A(n_475), .Y(n_739) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
AND2x2_ASAP7_75t_L g507 ( .A(n_476), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g694 ( .A(n_476), .Y(n_694) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g509 ( .A(n_477), .B(n_498), .Y(n_509) );
AND2x2_ASAP7_75t_L g571 ( .A(n_477), .B(n_485), .Y(n_571) );
INVx2_ASAP7_75t_L g576 ( .A(n_477), .Y(n_576) );
AND2x2_ASAP7_75t_L g578 ( .A(n_477), .B(n_486), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_483), .Y(n_478) );
INVx1_ASAP7_75t_L g556 ( .A(n_485), .Y(n_556) );
INVx2_ASAP7_75t_L g560 ( .A(n_485), .Y(n_560) );
AND2x4_ASAP7_75t_SL g591 ( .A(n_485), .B(n_498), .Y(n_591) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_485), .Y(n_623) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_486), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_492), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_507), .Y(n_494) );
AND2x2_ASAP7_75t_L g657 ( .A(n_495), .B(n_602), .Y(n_657) );
INVx2_ASAP7_75t_SL g745 ( .A(n_495), .Y(n_745) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_506), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g558 ( .A(n_497), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g665 ( .A(n_497), .B(n_578), .Y(n_665) );
INVx4_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g553 ( .A(n_498), .Y(n_553) );
AND2x4_ASAP7_75t_L g555 ( .A(n_498), .B(n_556), .Y(n_555) );
NOR2x1_ASAP7_75t_L g575 ( .A(n_498), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g648 ( .A(n_498), .Y(n_648) );
AND2x2_ASAP7_75t_L g667 ( .A(n_498), .B(n_606), .Y(n_667) );
AND2x2_ASAP7_75t_L g698 ( .A(n_498), .B(n_607), .Y(n_698) );
OR2x6_ASAP7_75t_L g498 ( .A(n_499), .B(n_505), .Y(n_498) );
AND2x2_ASAP7_75t_L g637 ( .A(n_507), .B(n_591), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_507), .B(n_648), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_507), .A2(n_748), .B1(n_750), .B2(n_751), .Y(n_747) );
AND2x2_ASAP7_75t_L g750 ( .A(n_507), .B(n_557), .Y(n_750) );
INVx3_ASAP7_75t_L g603 ( .A(n_508), .Y(n_603) );
AND2x2_ASAP7_75t_L g606 ( .A(n_508), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g622 ( .A(n_509), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g631 ( .A(n_509), .Y(n_631) );
AND2x4_ASAP7_75t_SL g510 ( .A(n_511), .B(n_520), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_511), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g682 ( .A(n_511), .B(n_683), .Y(n_682) );
NOR3xp33_ASAP7_75t_L g734 ( .A(n_511), .B(n_644), .C(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_L g752 ( .A(n_511), .B(n_646), .Y(n_752) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g567 ( .A(n_513), .B(n_531), .Y(n_567) );
INVx1_ASAP7_75t_L g584 ( .A(n_513), .Y(n_584) );
INVx2_ASAP7_75t_L g597 ( .A(n_513), .Y(n_597) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_513), .Y(n_612) );
AND2x2_ASAP7_75t_L g626 ( .A(n_513), .B(n_599), .Y(n_626) );
AND2x2_ASAP7_75t_L g705 ( .A(n_513), .B(n_522), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_520), .A2(n_569), .B1(n_572), .B2(n_579), .C(n_585), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_520), .A2(n_698), .B1(n_699), .B2(n_700), .C(n_701), .Y(n_697) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
INVx2_ASAP7_75t_L g639 ( .A(n_521), .Y(n_639) );
AND2x2_ASAP7_75t_L g699 ( .A(n_521), .B(n_583), .Y(n_699) );
AND2x2_ASAP7_75t_L g709 ( .A(n_521), .B(n_595), .Y(n_709) );
OR2x2_ASAP7_75t_L g749 ( .A(n_521), .B(n_633), .Y(n_749) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_SL g566 ( .A(n_522), .B(n_567), .Y(n_566) );
NAND2x1_ASAP7_75t_L g582 ( .A(n_522), .B(n_531), .Y(n_582) );
INVx4_ASAP7_75t_L g611 ( .A(n_522), .Y(n_611) );
OR2x2_ASAP7_75t_L g653 ( .A(n_522), .B(n_540), .Y(n_653) );
OR2x6_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
AND2x2_ASAP7_75t_L g704 ( .A(n_530), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_540), .Y(n_530) );
INVx2_ASAP7_75t_SL g592 ( .A(n_531), .Y(n_592) );
NOR2x1_ASAP7_75t_SL g598 ( .A(n_531), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g613 ( .A(n_531), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g644 ( .A(n_531), .B(n_611), .Y(n_644) );
AND2x2_ASAP7_75t_L g651 ( .A(n_531), .B(n_597), .Y(n_651) );
BUFx2_ASAP7_75t_L g685 ( .A(n_531), .Y(n_685) );
AND2x2_ASAP7_75t_L g696 ( .A(n_531), .B(n_611), .Y(n_696) );
OR2x6_ASAP7_75t_L g531 ( .A(n_532), .B(n_539), .Y(n_531) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_540), .Y(n_564) );
AND2x2_ASAP7_75t_L g583 ( .A(n_540), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g614 ( .A(n_540), .Y(n_614) );
AND2x2_ASAP7_75t_L g640 ( .A(n_540), .B(n_596), .Y(n_640) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_549), .Y(n_541) );
AO21x1_ASAP7_75t_SL g599 ( .A1(n_542), .A2(n_543), .B(n_549), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_548), .Y(n_543) );
OAI31xp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_555), .A3(n_557), .B(n_561), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx2_ASAP7_75t_L g659 ( .A(n_553), .Y(n_659) );
NOR2xp67_ASAP7_75t_L g569 ( .A(n_554), .B(n_570), .Y(n_569) );
AOI322xp5_ASAP7_75t_L g649 ( .A1(n_554), .A2(n_643), .A3(n_650), .B1(n_654), .B2(n_655), .C1(n_657), .C2(n_658), .Y(n_649) );
AND2x2_ASAP7_75t_L g721 ( .A(n_554), .B(n_698), .Y(n_721) );
AOI221xp5_ASAP7_75t_SL g634 ( .A1(n_555), .A2(n_635), .B1(n_637), .B2(n_638), .C(n_641), .Y(n_634) );
INVx2_ASAP7_75t_L g654 ( .A(n_555), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_557), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_557), .B(n_650), .Y(n_753) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g628 ( .A(n_558), .B(n_603), .Y(n_628) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g607 ( .A(n_560), .B(n_576), .Y(n_607) );
AND2x4_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g678 ( .A(n_564), .Y(n_678) );
O2A1O1Ixp5_ASAP7_75t_L g669 ( .A1(n_565), .A2(n_670), .B(n_672), .C(n_674), .Y(n_669) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_566), .A2(n_702), .B1(n_703), .B2(n_706), .Y(n_701) );
OR2x2_ASAP7_75t_L g656 ( .A(n_567), .B(n_653), .Y(n_656) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_573), .B(n_577), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g589 ( .A(n_576), .Y(n_589) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_578), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g632 ( .A(n_582), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_582), .B(n_583), .Y(n_675) );
OR2x2_ASAP7_75t_L g677 ( .A(n_582), .B(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_582), .B(n_726), .Y(n_725) );
BUFx2_ASAP7_75t_L g593 ( .A(n_584), .Y(n_593) );
NOR4xp25_ASAP7_75t_L g585 ( .A(n_586), .B(n_590), .C(n_592), .D(n_593), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g713 ( .A(n_587), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g741 ( .A(n_587), .B(n_590), .Y(n_741) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g671 ( .A(n_589), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_590), .B(n_619), .Y(n_706) );
AOI321xp33_ASAP7_75t_L g708 ( .A1(n_590), .A2(n_709), .A3(n_710), .B1(n_711), .B2(n_713), .C(n_716), .Y(n_708) );
INVx2_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_SL g670 ( .A(n_591), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_591), .B(n_630), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_592), .B(n_614), .Y(n_719) );
OR2x2_ASAP7_75t_L g746 ( .A(n_593), .B(n_630), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_600), .B(n_604), .Y(n_594) );
AND2x2_ASAP7_75t_L g635 ( .A(n_595), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g661 ( .A(n_597), .B(n_599), .Y(n_661) );
INVx2_ASAP7_75t_L g646 ( .A(n_598), .Y(n_646) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_601), .B(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g702 ( .A(n_602), .B(n_654), .Y(n_702) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g660 ( .A(n_603), .B(n_661), .Y(n_660) );
NOR2x1_ASAP7_75t_L g738 ( .A(n_603), .B(n_739), .Y(n_738) );
NOR2xp67_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g689 ( .A(n_607), .Y(n_689) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_613), .Y(n_609) );
NOR2xp67_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_611), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g636 ( .A(n_611), .Y(n_636) );
BUFx2_ASAP7_75t_L g718 ( .A(n_611), .Y(n_718) );
INVxp67_ASAP7_75t_L g726 ( .A(n_614), .Y(n_726) );
NAND3xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_634), .C(n_649), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_624), .B(n_627), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_621), .Y(n_617) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g647 ( .A(n_620), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g700 ( .A(n_621), .Y(n_700) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g715 ( .A(n_623), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_624), .A2(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_SL g633 ( .A(n_626), .Y(n_633) );
AND2x2_ASAP7_75t_L g695 ( .A(n_626), .B(n_696), .Y(n_695) );
AOI21xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B(n_632), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_628), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_674) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g664 ( .A(n_630), .Y(n_664) );
OR2x2_ASAP7_75t_L g712 ( .A(n_633), .B(n_644), .Y(n_712) );
NOR4xp25_ASAP7_75t_L g744 ( .A(n_636), .B(n_685), .C(n_745), .D(n_746), .Y(n_744) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
OR2x2_ASAP7_75t_L g645 ( .A(n_639), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_639), .B(n_661), .Y(n_743) );
AOI21xp33_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_645), .B(n_647), .Y(n_641) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g732 ( .A(n_644), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g740 ( .A(n_646), .Y(n_740) );
AND2x4_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVxp67_ASAP7_75t_L g668 ( .A(n_651), .Y(n_668) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g684 ( .A(n_653), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
AND2x2_ASAP7_75t_L g687 ( .A(n_659), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g733 ( .A(n_661), .Y(n_733) );
A2O1A1Ixp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_666), .B(n_668), .C(n_669), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g723 ( .A(n_665), .Y(n_723) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_L g727 ( .A(n_670), .Y(n_727) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_707), .C(n_728), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_686), .B(n_690), .C(n_697), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI21xp5_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_693), .B(n_695), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
O2A1O1Ixp33_ASAP7_75t_L g729 ( .A1(n_693), .A2(n_730), .B(n_731), .C(n_734), .Y(n_729) );
BUFx2_ASAP7_75t_L g710 ( .A(n_694), .Y(n_710) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_720), .Y(n_707) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_717), .A2(n_723), .B1(n_724), .B2(n_727), .Y(n_722) );
OR2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND4xp25_ASAP7_75t_L g728 ( .A(n_729), .B(n_737), .C(n_747), .D(n_753), .Y(n_728) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_740), .B1(n_741), .B2(n_742), .C(n_744), .Y(n_737) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
CKINVDCx11_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
INVxp67_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
BUFx3_ASAP7_75t_L g777 ( .A(n_767), .Y(n_777) );
INVx2_ASAP7_75t_L g774 ( .A(n_769), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
endmodule