module fake_jpeg_9503_n_278 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_40),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_58),
.C(n_15),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_25),
.B1(n_31),
.B2(n_24),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_49),
.B1(n_56),
.B2(n_60),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_25),
.B1(n_20),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_57),
.B1(n_59),
.B2(n_15),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_25),
.B1(n_31),
.B2(n_24),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_55),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_25),
.B1(n_31),
.B2(n_20),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_27),
.B1(n_19),
.B2(n_30),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_20),
.B(n_23),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_15),
.B1(n_30),
.B2(n_19),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_30),
.B1(n_17),
.B2(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_18),
.B1(n_19),
.B2(n_17),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_63),
.B1(n_15),
.B2(n_26),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_17),
.B1(n_18),
.B2(n_27),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_73),
.A2(n_79),
.B1(n_85),
.B2(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_50),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_53),
.B1(n_43),
.B2(n_64),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_63),
.B1(n_62),
.B2(n_60),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_16),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_39),
.B1(n_34),
.B2(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_16),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_81),
.B(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_38),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_38),
.Y(n_84)
);

AO22x1_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_38),
.B1(n_35),
.B2(n_32),
.Y(n_85)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_44),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_104),
.B(n_101),
.C(n_97),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_99),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_58),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_92),
.C(n_65),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_49),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_70),
.A2(n_46),
.B1(n_45),
.B2(n_50),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_82),
.B1(n_80),
.B2(n_53),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_96),
.B(n_106),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_97),
.A2(n_28),
.B(n_26),
.Y(n_126)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_11),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_73),
.B1(n_75),
.B2(n_78),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_72),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_85),
.B1(n_69),
.B2(n_68),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_113),
.B1(n_119),
.B2(n_123),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_88),
.C(n_97),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_84),
.B(n_68),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_112),
.B(n_32),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_79),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_66),
.B1(n_100),
.B2(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_116),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_89),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_52),
.B1(n_43),
.B2(n_64),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_120),
.B1(n_128),
.B2(n_122),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_86),
.A2(n_52),
.B1(n_43),
.B2(n_64),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_51),
.B1(n_72),
.B2(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_127),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_51),
.B1(n_72),
.B2(n_66),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_87),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_130),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_77),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_136),
.B1(n_145),
.B2(n_152),
.Y(n_157)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_134),
.B(n_139),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_110),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_128),
.A2(n_86),
.B1(n_104),
.B2(n_88),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_151),
.C(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_153),
.Y(n_162)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_95),
.B1(n_102),
.B2(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_108),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_95),
.B1(n_102),
.B2(n_51),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_115),
.B1(n_118),
.B2(n_116),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_149),
.B(n_120),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_66),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_109),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_131),
.Y(n_163)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_179),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_168),
.Y(n_189)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_111),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_166),
.C(n_171),
.Y(n_183)
);

XOR2x1_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_175),
.B1(n_28),
.B2(n_32),
.Y(n_195)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_172),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_112),
.C(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_103),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_125),
.B1(n_112),
.B2(n_114),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_177),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_147),
.B(n_124),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_124),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_187),
.C(n_200),
.Y(n_202)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_23),
.B(n_61),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_146),
.B1(n_144),
.B2(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_149),
.C(n_136),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_138),
.B(n_126),
.C(n_130),
.D(n_48),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_173),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_140),
.B1(n_100),
.B2(n_27),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_194),
.B1(n_196),
.B2(n_201),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_157),
.A2(n_28),
.B1(n_109),
.B2(n_29),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_198),
.B1(n_174),
.B2(n_156),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_167),
.B1(n_175),
.B2(n_168),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_177),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_167),
.A2(n_48),
.B1(n_61),
.B2(n_71),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_48),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_178),
.B1(n_159),
.B2(n_170),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_180),
.C(n_200),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_208),
.C(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_156),
.B1(n_158),
.B2(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_171),
.C(n_160),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_184),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_215),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_219),
.Y(n_232)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_29),
.A3(n_22),
.B1(n_23),
.B2(n_35),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_213),
.B1(n_23),
.B2(n_29),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_61),
.C(n_71),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_71),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_188),
.A3(n_190),
.B1(n_191),
.B2(n_195),
.C1(n_189),
.C2(n_193),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_0),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_217),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_218),
.B(n_198),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

MAJx2_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_190),
.C(n_199),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_229),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_189),
.B1(n_181),
.B2(n_193),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_217),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_214),
.A2(n_71),
.B1(n_14),
.B2(n_13),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_203),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_35),
.C(n_29),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_233),
.C(n_0),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_29),
.C(n_22),
.Y(n_233)
);

AOI31xp67_ASAP7_75t_SL g235 ( 
.A1(n_217),
.A2(n_22),
.A3(n_14),
.B(n_13),
.Y(n_235)
);

OAI211xp5_ASAP7_75t_L g236 ( 
.A1(n_235),
.A2(n_221),
.B(n_218),
.C(n_14),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_226),
.Y(n_237)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_223),
.B(n_204),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_241),
.Y(n_249)
);

AND2x6_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_219),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_12),
.B(n_11),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_232),
.B(n_206),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_218),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_243),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_228),
.B1(n_220),
.B2(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_12),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_1),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_233),
.B(n_12),
.Y(n_253)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_1),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_11),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_242),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_262),
.B(n_251),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_248),
.Y(n_262)
);

AO21x1_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_255),
.B(n_239),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_265),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_240),
.Y(n_264)
);

OAI221xp5_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_266),
.B1(n_240),
.B2(n_250),
.C(n_3),
.Y(n_269)
);

OAI33xp33_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_269),
.A3(n_270),
.B1(n_271),
.B2(n_10),
.B3(n_7),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_253),
.B(n_252),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_268),
.A2(n_260),
.B1(n_6),
.B2(n_7),
.Y(n_272)
);

AOI322xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_273),
.C(n_274),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_4),
.C(n_8),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_8),
.C(n_9),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_276),
.A2(n_275),
.B1(n_8),
.B2(n_9),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_9),
.Y(n_278)
);


endmodule