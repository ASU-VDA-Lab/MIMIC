module fake_netlist_5_1088_n_107 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_107);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_107;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_1),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_34),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_2),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_23),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_27),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

AO22x2_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

AO22x2_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_20),
.B1(n_26),
.B2(n_31),
.Y(n_52)
);

NAND2x1p5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_39),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_43),
.B1(n_28),
.B2(n_21),
.Y(n_60)
);

AND2x4_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_52),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_56),
.B(n_46),
.C(n_39),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_41),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_44),
.B(n_37),
.C(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_53),
.Y(n_69)
);

OAI211xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_44),
.B(n_60),
.C(n_37),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_58),
.B(n_59),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_52),
.Y(n_72)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_62),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_69),
.B1(n_66),
.B2(n_68),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_77),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_71),
.B(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_82),
.A2(n_53),
.B(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_81),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_84),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_67),
.B1(n_72),
.B2(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_92),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_91),
.A2(n_88),
.B(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_50),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_72),
.C(n_71),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_85),
.B(n_50),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_9),
.Y(n_101)
);

OAI221xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_97),
.B1(n_93),
.B2(n_28),
.C(n_74),
.Y(n_102)
);

NAND4xp25_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_99),
.C(n_101),
.D(n_74),
.Y(n_103)
);

AOI211xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_98),
.B(n_10),
.C(n_9),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_10),
.B1(n_51),
.B2(n_14),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);


endmodule