module fake_netlist_6_4922_n_107 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_19, n_107);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;
input n_19;

output n_107;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVxp33_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_R g44 ( 
.A(n_30),
.B(n_3),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_32),
.Y(n_53)
);

OAI221xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_35),
.B1(n_26),
.B2(n_29),
.C(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_31),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_22),
.B(n_4),
.C(n_5),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_43),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_39),
.B(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_14),
.Y(n_60)
);

OAI21x1_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_16),
.B(n_17),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_44),
.Y(n_63)
);

AND2x4_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_57),
.Y(n_64)
);

NAND2x1p5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_56),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NAND2x1p5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_54),
.Y(n_68)
);

OAI21x1_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_52),
.B(n_4),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_67),
.B(n_52),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_58),
.Y(n_71)
);

INVxp67_ASAP7_75t_SL g72 ( 
.A(n_67),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_36),
.B1(n_37),
.B2(n_47),
.Y(n_74)
);

AOI31xp33_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_44),
.A3(n_8),
.B(n_7),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_68),
.C(n_64),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_64),
.Y(n_77)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_65),
.B(n_69),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_74),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_76),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_64),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_66),
.C(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_88),
.B1(n_83),
.B2(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_90),
.B(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

AO21x1_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_85),
.B(n_65),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_85),
.B1(n_66),
.B2(n_84),
.C(n_65),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_78),
.B(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_101),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_R g104 ( 
.A(n_103),
.B(n_93),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_100),
.B1(n_94),
.B2(n_97),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_99),
.B1(n_66),
.B2(n_78),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_78),
.B(n_66),
.Y(n_107)
);


endmodule