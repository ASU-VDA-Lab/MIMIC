module fake_netlist_1_10653_n_669 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_669);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_669;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_23), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_2), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_69), .Y(n_79) );
BUFx3_ASAP7_75t_L g80 ( .A(n_30), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_48), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_26), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_3), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_62), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_44), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_21), .Y(n_86) );
BUFx3_ASAP7_75t_L g87 ( .A(n_59), .Y(n_87) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_28), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_24), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_10), .Y(n_90) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_4), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_4), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_50), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_17), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_34), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_35), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_1), .Y(n_97) );
BUFx5_ASAP7_75t_L g98 ( .A(n_67), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_18), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_51), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_13), .Y(n_101) );
BUFx2_ASAP7_75t_L g102 ( .A(n_43), .Y(n_102) );
CKINVDCx14_ASAP7_75t_R g103 ( .A(n_38), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_9), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_37), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_29), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_49), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_1), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_55), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_14), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_61), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_70), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_60), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_32), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_41), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_12), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_57), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_11), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_25), .Y(n_121) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_101), .A2(n_0), .B1(n_3), .B2(n_5), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_102), .B(n_103), .Y(n_123) );
OA21x2_ASAP7_75t_L g124 ( .A1(n_77), .A2(n_40), .B(n_75), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_91), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_98), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_98), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_98), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_119), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_119), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_79), .B(n_0), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_98), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_103), .B(n_5), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_81), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_98), .B(n_6), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_119), .Y(n_137) );
NAND2xp33_ASAP7_75t_R g138 ( .A(n_82), .B(n_42), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_119), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_101), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_98), .Y(n_141) );
NAND2xp33_ASAP7_75t_L g142 ( .A(n_98), .B(n_45), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_78), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_119), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_80), .B(n_7), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_80), .B(n_9), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_95), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_83), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_109), .B(n_10), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_87), .B(n_11), .Y(n_151) );
OAI22xp5_ASAP7_75t_SL g152 ( .A1(n_109), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_87), .B(n_53), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_117), .B(n_90), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_92), .B(n_15), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_88), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_99), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_100), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_88), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_107), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_110), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_150), .A2(n_114), .B1(n_120), .B2(n_118), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_123), .B(n_134), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_123), .B(n_105), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_153), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_129), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_126), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_134), .B(n_121), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_155), .B(n_82), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_133), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_129), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_125), .B(n_105), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_129), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_155), .B(n_84), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_126), .Y(n_179) );
BUFx4f_ASAP7_75t_L g180 ( .A(n_153), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_136), .B(n_116), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_147), .B(n_84), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_147), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_136), .B(n_85), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_129), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_145), .B(n_148), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_129), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_127), .Y(n_190) );
NOR2xp33_ASAP7_75t_SL g191 ( .A(n_133), .B(n_114), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_127), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_147), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_150), .B(n_85), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_145), .B(n_112), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_128), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_151), .B(n_94), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_148), .B(n_112), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_143), .B(n_94), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_130), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_151), .A2(n_104), .B1(n_113), .B2(n_111), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_151), .A2(n_108), .B1(n_97), .B2(n_93), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_128), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_132), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_149), .B(n_115), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_158), .B(n_162), .Y(n_206) );
NOR2x1p5_ASAP7_75t_L g207 ( .A(n_156), .B(n_88), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_158), .B(n_106), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_130), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_132), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_159), .B(n_96), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_141), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_171), .B(n_162), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_204), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_177), .B(n_161), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_170), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_164), .B(n_161), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_194), .A2(n_122), .B1(n_131), .B2(n_140), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_170), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_186), .B(n_159), .Y(n_220) );
INVx5_ASAP7_75t_L g221 ( .A(n_170), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_204), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_180), .A2(n_142), .B(n_124), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_195), .B(n_153), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_198), .B(n_153), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_193), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_194), .B(n_154), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_193), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_199), .B(n_154), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_211), .B(n_141), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_180), .A2(n_142), .B(n_124), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_206), .Y(n_232) );
NAND2x1p5_ASAP7_75t_L g233 ( .A(n_184), .B(n_135), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_201), .A2(n_152), .B1(n_124), .B2(n_88), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_170), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_207), .B(n_15), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_165), .B(n_124), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_172), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_204), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_184), .B(n_144), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_184), .B(n_144), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_204), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_188), .B(n_160), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_205), .B(n_160), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_207), .B(n_16), .Y(n_245) );
OR2x6_ASAP7_75t_L g246 ( .A(n_183), .B(n_138), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_172), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_172), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_172), .A2(n_160), .B1(n_157), .B2(n_144), .Y(n_249) );
AO22x1_ASAP7_75t_L g250 ( .A1(n_173), .A2(n_16), .B1(n_160), .B2(n_157), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_212), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_202), .B(n_160), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_182), .A2(n_157), .B1(n_144), .B2(n_139), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_197), .B(n_157), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_182), .B(n_157), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_182), .A2(n_144), .B1(n_139), .B2(n_137), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_184), .B(n_137), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_182), .B(n_139), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_185), .B(n_139), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_185), .B(n_139), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_208), .B(n_137), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_163), .A2(n_137), .B1(n_130), .B2(n_22), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_163), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_180), .B(n_130), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_185), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_166), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_175), .B(n_137), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_185), .A2(n_130), .B1(n_20), .B2(n_27), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_180), .A2(n_19), .B1(n_31), .B2(n_33), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_212), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_212), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_SL g272 ( .A1(n_237), .A2(n_169), .B(n_181), .C(n_212), .Y(n_272) );
NOR3xp33_ASAP7_75t_L g273 ( .A(n_263), .B(n_191), .C(n_179), .Y(n_273) );
OR2x4_ASAP7_75t_L g274 ( .A(n_217), .B(n_210), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_219), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_218), .B(n_210), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_266), .B(n_166), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_237), .A2(n_166), .B(n_178), .C(n_192), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_236), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_219), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_223), .A2(n_178), .B(n_192), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_219), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_213), .B(n_179), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_267), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_221), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_266), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_216), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_221), .B(n_178), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_231), .A2(n_190), .B(n_203), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_246), .A2(n_190), .B1(n_203), .B2(n_168), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_215), .B(n_196), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_221), .B(n_196), .Y(n_292) );
BUFx12f_ASAP7_75t_L g293 ( .A(n_236), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g294 ( .A1(n_227), .A2(n_168), .B1(n_167), .B2(n_187), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_232), .B(n_36), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_224), .A2(n_187), .B(n_176), .Y(n_296) );
NAND3xp33_ASAP7_75t_SL g297 ( .A(n_262), .B(n_187), .C(n_176), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_216), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_246), .A2(n_176), .B1(n_174), .B2(n_167), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_220), .A2(n_174), .B1(n_167), .B2(n_189), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_225), .A2(n_174), .B(n_200), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_238), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_L g303 ( .A1(n_234), .A2(n_39), .B(n_46), .C(n_47), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_240), .A2(n_200), .B(n_189), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g305 ( .A1(n_252), .A2(n_52), .B(n_54), .C(n_56), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_246), .B(n_58), .Y(n_306) );
O2A1O1Ixp5_ASAP7_75t_L g307 ( .A1(n_264), .A2(n_209), .B(n_200), .C(n_189), .Y(n_307) );
AND2x4_ASAP7_75t_SL g308 ( .A(n_236), .B(n_209), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_238), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_245), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_240), .A2(n_200), .B(n_189), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_247), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_230), .B(n_63), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_247), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_226), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_267), .B(n_64), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_229), .B(n_65), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_241), .A2(n_209), .B(n_200), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_267), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_241), .A2(n_209), .B(n_200), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_228), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_275), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_276), .B(n_221), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_315), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_285), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_281), .A2(n_257), .B(n_264), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_289), .A2(n_257), .B(n_259), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_293), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_274), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_273), .A2(n_245), .B1(n_265), .B2(n_248), .Y(n_330) );
INVx4_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_274), .B(n_235), .Y(n_332) );
AO31x2_ASAP7_75t_L g333 ( .A1(n_289), .A2(n_269), .A3(n_243), .B(n_260), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_280), .Y(n_334) );
AO31x2_ASAP7_75t_L g335 ( .A1(n_278), .A2(n_258), .A3(n_255), .B(n_244), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_283), .B(n_245), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_SL g337 ( .A1(n_272), .A2(n_268), .B(n_254), .C(n_271), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g338 ( .A1(n_281), .A2(n_233), .B(n_271), .Y(n_338) );
OR2x6_ASAP7_75t_L g339 ( .A(n_310), .B(n_250), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_321), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_279), .A2(n_261), .B(n_233), .C(n_270), .Y(n_341) );
AO31x2_ASAP7_75t_L g342 ( .A1(n_301), .A2(n_214), .A3(n_251), .B(n_242), .Y(n_342) );
BUFx12f_ASAP7_75t_L g343 ( .A(n_319), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_286), .Y(n_344) );
AO21x1_ASAP7_75t_L g345 ( .A1(n_303), .A2(n_261), .B(n_270), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_291), .B(n_261), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_284), .A2(n_242), .B1(n_222), .B2(n_251), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_306), .A2(n_239), .B1(n_222), .B2(n_214), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_305), .A2(n_239), .B(n_249), .C(n_253), .Y(n_349) );
A2O1A1Ixp33_ASAP7_75t_L g350 ( .A1(n_295), .A2(n_249), .B(n_253), .C(n_256), .Y(n_350) );
O2A1O1Ixp33_ASAP7_75t_L g351 ( .A1(n_317), .A2(n_256), .B(n_68), .C(n_71), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_287), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_298), .B(n_66), .Y(n_353) );
A2O1A1Ixp33_ASAP7_75t_L g354 ( .A1(n_316), .A2(n_189), .B(n_209), .C(n_74), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_324), .B(n_314), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_336), .B(n_286), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_323), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_344), .Y(n_358) );
OAI211xp5_ASAP7_75t_SL g359 ( .A1(n_329), .A2(n_299), .B(n_290), .C(n_292), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_339), .Y(n_360) );
AOI21xp33_ASAP7_75t_L g361 ( .A1(n_341), .A2(n_313), .B(n_294), .Y(n_361) );
NOR2xp67_ASAP7_75t_L g362 ( .A(n_331), .B(n_302), .Y(n_362) );
OAI22x1_ASAP7_75t_L g363 ( .A1(n_353), .A2(n_312), .B1(n_309), .B2(n_282), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_330), .A2(n_323), .B1(n_343), .B2(n_339), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_331), .B(n_286), .Y(n_365) );
OA21x2_ASAP7_75t_L g366 ( .A1(n_354), .A2(n_301), .B(n_307), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_344), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_337), .A2(n_318), .B(n_311), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_337), .A2(n_318), .B(n_311), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_340), .Y(n_370) );
NAND2x1p5_ASAP7_75t_L g371 ( .A(n_344), .B(n_288), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_322), .Y(n_372) );
OAI21x1_ASAP7_75t_L g373 ( .A1(n_338), .A2(n_320), .B(n_304), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_322), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_334), .Y(n_375) );
OA21x2_ASAP7_75t_L g376 ( .A1(n_354), .A2(n_320), .B(n_304), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_326), .A2(n_296), .B(n_297), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_342), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_327), .A2(n_296), .B(n_300), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_349), .A2(n_277), .B(n_308), .Y(n_380) );
INVx2_ASAP7_75t_SL g381 ( .A(n_344), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_368), .A2(n_349), .B(n_345), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_372), .B(n_335), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_380), .A2(n_330), .B(n_346), .Y(n_384) );
AOI21xp5_ASAP7_75t_SL g385 ( .A1(n_363), .A2(n_339), .B(n_353), .Y(n_385) );
CKINVDCx16_ASAP7_75t_R g386 ( .A(n_360), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_378), .Y(n_387) );
AO21x2_ASAP7_75t_L g388 ( .A1(n_369), .A2(n_348), .B(n_350), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_358), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_372), .B(n_335), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_374), .B(n_335), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_374), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_378), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g394 ( .A1(n_364), .A2(n_332), .B1(n_352), .B2(n_347), .C(n_351), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_357), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_373), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_375), .B(n_335), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_375), .B(n_342), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_373), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g400 ( .A1(n_377), .A2(n_350), .B(n_347), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_379), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_370), .A2(n_328), .B1(n_325), .B2(n_334), .C(n_189), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_370), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_360), .B(n_333), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_363), .A2(n_325), .B1(n_333), .B2(n_342), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_358), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_358), .B(n_342), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_355), .B(n_356), .Y(n_409) );
OA21x2_ASAP7_75t_L g410 ( .A1(n_361), .A2(n_333), .B(n_209), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_359), .A2(n_333), .B1(n_73), .B2(n_76), .Y(n_411) );
OA21x2_ASAP7_75t_L g412 ( .A1(n_367), .A2(n_72), .B(n_381), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_358), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_398), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_404), .B(n_365), .Y(n_415) );
AND2x2_ASAP7_75t_SL g416 ( .A(n_412), .B(n_365), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_398), .B(n_367), .Y(n_417) );
INVxp67_ASAP7_75t_L g418 ( .A(n_404), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_398), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_387), .B(n_381), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_383), .B(n_376), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_412), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_383), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_383), .B(n_376), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_397), .B(n_376), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_397), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_395), .B(n_365), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_390), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_390), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_394), .A2(n_365), .B1(n_362), .B2(n_376), .Y(n_431) );
INVx4_ASAP7_75t_L g432 ( .A(n_412), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_387), .B(n_371), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_412), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_408), .B(n_366), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_408), .B(n_362), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_392), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_392), .Y(n_438) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_401), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_408), .B(n_371), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_409), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_389), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_409), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_393), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_393), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_386), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_409), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_393), .B(n_390), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_405), .B(n_371), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_391), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_391), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_405), .B(n_366), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_413), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_386), .B(n_366), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_400), .B(n_366), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_413), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_400), .B(n_388), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_395), .A2(n_412), .B1(n_394), .B2(n_385), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_414), .B(n_399), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_437), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_444), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_414), .B(n_399), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_420), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_438), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_420), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_441), .B(n_384), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_423), .B(n_399), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_423), .B(n_396), .Y(n_468) );
INVx2_ASAP7_75t_SL g469 ( .A(n_436), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_444), .Y(n_470) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_432), .B(n_412), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_426), .B(n_396), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_453), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_419), .B(n_396), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_426), .B(n_427), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_446), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_417), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_427), .B(n_410), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_453), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_436), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_443), .B(n_384), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_447), .B(n_406), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_417), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_421), .B(n_410), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_418), .B(n_406), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_421), .B(n_402), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_436), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_424), .B(n_410), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_456), .Y(n_489) );
NOR2xp33_ASAP7_75t_SL g490 ( .A(n_416), .B(n_432), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_424), .B(n_410), .Y(n_491) );
INVxp33_ASAP7_75t_L g492 ( .A(n_428), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_425), .B(n_410), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_445), .Y(n_494) );
AND2x6_ASAP7_75t_SL g495 ( .A(n_415), .B(n_403), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_456), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_433), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_425), .B(n_402), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_429), .B(n_389), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_435), .B(n_402), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_445), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_433), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_429), .B(n_382), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_435), .B(n_401), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_430), .B(n_448), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_450), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_448), .B(n_401), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_430), .B(n_389), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_439), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_451), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_457), .B(n_382), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_451), .B(n_457), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_449), .B(n_382), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_460), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_465), .B(n_449), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_460), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_512), .B(n_452), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_492), .B(n_454), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_465), .B(n_440), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_464), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_464), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_477), .B(n_440), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_483), .B(n_440), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_473), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_473), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_505), .B(n_452), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_463), .B(n_455), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_479), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_512), .B(n_455), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_500), .B(n_432), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_461), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_461), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_461), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_469), .B(n_434), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_469), .B(n_434), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_463), .B(n_442), .Y(n_537) );
INVx4_ASAP7_75t_L g538 ( .A(n_495), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_513), .B(n_442), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_497), .B(n_422), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_476), .A2(n_458), .B1(n_416), .B2(n_431), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_495), .B(n_434), .Y(n_542) );
NAND2x1_ASAP7_75t_L g543 ( .A(n_471), .B(n_422), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_475), .B(n_422), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_475), .B(n_388), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_502), .B(n_389), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_497), .B(n_389), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_480), .B(n_407), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_498), .B(n_382), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_500), .B(n_439), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_479), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_504), .B(n_439), .Y(n_552) );
OAI221xp5_ASAP7_75t_L g553 ( .A1(n_485), .A2(n_411), .B1(n_403), .B2(n_407), .C(n_439), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_504), .B(n_439), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_484), .B(n_382), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_498), .B(n_388), .Y(n_556) );
OR3x2_ASAP7_75t_L g557 ( .A(n_514), .B(n_411), .C(n_388), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_506), .B(n_388), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_470), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_506), .B(n_407), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_474), .B(n_407), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_470), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_489), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_474), .B(n_407), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_480), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_484), .B(n_493), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_488), .B(n_491), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_488), .B(n_491), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_566), .B(n_567), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_566), .B(n_493), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_515), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_567), .B(n_487), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_568), .B(n_487), .Y(n_573) );
NAND2x1_ASAP7_75t_L g574 ( .A(n_565), .B(n_471), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_535), .B(n_486), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_527), .B(n_514), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_530), .B(n_482), .Y(n_577) );
INVxp67_ASAP7_75t_L g578 ( .A(n_542), .Y(n_578) );
A2O1A1Ixp33_ASAP7_75t_L g579 ( .A1(n_542), .A2(n_490), .B(n_511), .C(n_507), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_538), .A2(n_511), .B1(n_507), .B2(n_466), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_517), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_538), .B(n_481), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_521), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_568), .B(n_486), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_518), .B(n_503), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_522), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_532), .Y(n_587) );
INVx2_ASAP7_75t_SL g588 ( .A(n_565), .Y(n_588) );
OAI21xp33_ASAP7_75t_L g589 ( .A1(n_541), .A2(n_490), .B(n_503), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_538), .B(n_478), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_530), .B(n_489), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_525), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_555), .B(n_486), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_518), .B(n_486), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_555), .B(n_496), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_519), .B(n_496), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_531), .B(n_508), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_541), .A2(n_478), .B1(n_509), .B2(n_499), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_526), .Y(n_599) );
NAND2xp33_ASAP7_75t_L g600 ( .A(n_531), .B(n_508), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_529), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_544), .B(n_459), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_535), .B(n_470), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_516), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_519), .B(n_459), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_545), .B(n_462), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_551), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_578), .B(n_539), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_582), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_571), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_604), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_569), .Y(n_612) );
AOI211xp5_ASAP7_75t_L g613 ( .A1(n_589), .A2(n_553), .B(n_524), .C(n_523), .Y(n_613) );
OAI211xp5_ASAP7_75t_SL g614 ( .A1(n_582), .A2(n_537), .B(n_549), .C(n_558), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_598), .A2(n_543), .B(n_560), .C(n_563), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_600), .A2(n_536), .B1(n_535), .B2(n_557), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_580), .A2(n_557), .B1(n_536), .B2(n_528), .C(n_546), .Y(n_617) );
XOR2x2_ASAP7_75t_L g618 ( .A(n_590), .B(n_520), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_581), .Y(n_619) );
A2O1A1Ixp33_ASAP7_75t_SL g620 ( .A1(n_596), .A2(n_533), .B(n_532), .C(n_534), .Y(n_620) );
OAI211xp5_ASAP7_75t_L g621 ( .A1(n_590), .A2(n_556), .B(n_540), .C(n_548), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_579), .A2(n_536), .B(n_559), .Y(n_622) );
BUFx4f_ASAP7_75t_SL g623 ( .A(n_588), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_569), .B(n_554), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_583), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_579), .A2(n_559), .B(n_561), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_570), .B(n_554), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_596), .B(n_552), .Y(n_628) );
OAI31xp33_ASAP7_75t_L g629 ( .A1(n_603), .A2(n_552), .A3(n_550), .B(n_547), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_577), .B(n_550), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_570), .B(n_564), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_610), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_617), .A2(n_600), .B1(n_605), .B2(n_575), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_613), .B(n_595), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_609), .A2(n_575), .B1(n_576), .B2(n_593), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_611), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_615), .B(n_574), .C(n_603), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_623), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_623), .A2(n_575), .B1(n_588), .B2(n_585), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_619), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_625), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_630), .Y(n_642) );
NOR2x1_ASAP7_75t_L g643 ( .A(n_621), .B(n_622), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_612), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_628), .Y(n_645) );
AOI222xp33_ASAP7_75t_L g646 ( .A1(n_643), .A2(n_618), .B1(n_614), .B2(n_608), .C1(n_620), .C2(n_586), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_638), .B(n_608), .Y(n_647) );
AOI211x1_ASAP7_75t_L g648 ( .A1(n_639), .A2(n_626), .B(n_624), .C(n_618), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g649 ( .A1(n_633), .A2(n_616), .B1(n_629), .B2(n_620), .C(n_591), .Y(n_649) );
NAND4xp25_ASAP7_75t_L g650 ( .A(n_636), .B(n_572), .C(n_573), .D(n_606), .Y(n_650) );
AOI222xp33_ASAP7_75t_L g651 ( .A1(n_634), .A2(n_599), .B1(n_607), .B2(n_592), .C1(n_601), .C2(n_593), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_637), .A2(n_584), .B(n_627), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_639), .A2(n_594), .B(n_631), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_646), .B(n_635), .C(n_644), .D(n_645), .Y(n_654) );
NAND5xp2_ASAP7_75t_L g655 ( .A(n_652), .B(n_642), .C(n_641), .D(n_640), .E(n_632), .Y(n_655) );
OAI211xp5_ASAP7_75t_L g656 ( .A1(n_648), .A2(n_651), .B(n_647), .C(n_649), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_650), .B(n_587), .C(n_562), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_653), .A2(n_602), .B1(n_597), .B2(n_587), .C(n_472), .Y(n_658) );
NAND4xp75_ASAP7_75t_L g659 ( .A(n_656), .B(n_602), .C(n_467), .D(n_468), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_658), .B(n_562), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_657), .B(n_462), .Y(n_661) );
AOI22x1_ASAP7_75t_L g662 ( .A1(n_659), .A2(n_654), .B1(n_655), .B2(n_534), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g663 ( .A(n_660), .B(n_533), .C(n_510), .Y(n_663) );
XNOR2x1_ASAP7_75t_L g664 ( .A(n_662), .B(n_661), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_664), .Y(n_665) );
AOI222xp33_ASAP7_75t_L g666 ( .A1(n_665), .A2(n_663), .B1(n_510), .B2(n_472), .C1(n_468), .C2(n_467), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_666), .B(n_510), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_667), .A2(n_494), .B(n_501), .C(n_665), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_494), .B1(n_501), .B2(n_665), .Y(n_669) );
endmodule