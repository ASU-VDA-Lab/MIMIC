module real_jpeg_30134_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_315, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_315;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_0),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_0),
.A2(n_56),
.B1(n_62),
.B2(n_63),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_1),
.Y(n_92)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_1),
.Y(n_95)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_1),
.Y(n_242)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_3),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_69),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_69),
.Y(n_110)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_5),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_5),
.A2(n_32),
.B(n_36),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_5),
.B(n_34),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_5),
.A2(n_53),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_5),
.B(n_53),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_5),
.B(n_57),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_5),
.A2(n_90),
.B1(n_238),
.B2(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_5),
.A2(n_35),
.B(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_6),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_158),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_158),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_158),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_7),
.A2(n_40),
.B1(n_53),
.B2(n_54),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_7),
.A2(n_40),
.B1(n_62),
.B2(n_63),
.Y(n_163)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_9),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_101),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_101),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_101),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_10),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_10),
.A2(n_29),
.B1(n_53),
.B2(n_54),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_10),
.A2(n_29),
.B1(n_62),
.B2(n_63),
.Y(n_171)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_12),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_135),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_135),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_135),
.Y(n_258)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_14),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_14),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_15),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_147),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_15),
.A2(n_53),
.B1(n_54),
.B2(n_147),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_147),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_16),
.A2(n_35),
.B1(n_36),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_16),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_16),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_16),
.A2(n_46),
.B1(n_62),
.B2(n_63),
.Y(n_164)
);

INVx11_ASAP7_75t_SL g65 ( 
.A(n_17),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_115),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_102),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_22),
.B(n_102),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_73),
.C(n_79),
.Y(n_22)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_23),
.B(n_73),
.CI(n_79),
.CON(n_136),
.SN(n_136)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_72),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_24),
.A2(n_25),
.B1(n_104),
.B2(n_112),
.Y(n_103)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_25),
.B(n_43),
.C(n_71),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_39),
.B2(n_41),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_26),
.A2(n_30),
.B1(n_41),
.B2(n_99),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_32),
.Y(n_33)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_28),
.A2(n_38),
.B(n_156),
.C(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_30),
.A2(n_41),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_31),
.A2(n_34),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_31),
.A2(n_34),
.B1(n_100),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_31),
.A2(n_34),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_31),
.A2(n_34),
.B1(n_134),
.B2(n_186),
.Y(n_200)
);

AO22x1_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_49),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g262 ( 
.A1(n_35),
.A2(n_54),
.A3(n_255),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_36),
.B(n_156),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_39),
.Y(n_106)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_58),
.B1(n_70),
.B2(n_71),
.Y(n_42)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_55),
.B2(n_57),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_48),
.B1(n_52),
.B2(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_47),
.A2(n_55),
.B1(n_57),
.B2(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_47),
.A2(n_57),
.B1(n_76),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_47),
.A2(n_57),
.B1(n_146),
.B2(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_47),
.A2(n_57),
.B1(n_132),
.B2(n_189),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_48),
.A2(n_52),
.B1(n_145),
.B2(n_148),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_48),
.A2(n_52),
.B1(n_148),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_48),
.A2(n_52),
.B1(n_169),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_54),
.B1(n_60),
.B2(n_61),
.Y(n_67)
);

OAI32xp33_ASAP7_75t_L g215 ( 
.A1(n_53),
.A2(n_60),
.A3(n_63),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_53),
.B(n_266),
.Y(n_265)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_58),
.A2(n_71),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_66),
.B(n_68),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_66),
.B1(n_68),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_59),
.A2(n_66),
.B1(n_85),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_59),
.A2(n_66),
.B1(n_130),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_59),
.A2(n_66),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_59),
.A2(n_66),
.B1(n_213),
.B2(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_59),
.B(n_156),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_59),
.A2(n_66),
.B1(n_152),
.B2(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_61),
.B(n_62),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_62),
.B(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_74),
.B(n_77),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_97),
.B(n_98),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_81),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_89),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_82),
.A2(n_83),
.B1(n_89),
.B2(n_97),
.Y(n_295)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_86),
.A2(n_88),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_86),
.A2(n_88),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_97),
.B1(n_98),
.B2(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B(n_96),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_96),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_90),
.A2(n_127),
.B1(n_128),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_90),
.A2(n_128),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_90),
.A2(n_128),
.B1(n_232),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_90),
.A2(n_128),
.B1(n_227),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_91),
.A2(n_94),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_91),
.A2(n_94),
.B1(n_163),
.B2(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_91),
.A2(n_94),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

INVx5_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_95),
.B(n_156),
.Y(n_244)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_113),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_109),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_137),
.B(n_311),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_136),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_117),
.B(n_136),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_123),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_118),
.B(n_122),
.Y(n_299)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_123),
.A2(n_124),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_131),
.C(n_133),
.Y(n_124)
);

FAx1_ASAP7_75t_L g294 ( 
.A(n_125),
.B(n_131),
.CI(n_133),
.CON(n_294),
.SN(n_294)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_126),
.B(n_129),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_136),
.Y(n_313)
);

AOI321xp33_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_292),
.A3(n_300),
.B1(n_305),
.B2(n_310),
.C(n_315),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_191),
.C(n_203),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_173),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_140),
.B(n_173),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_159),
.C(n_165),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_141),
.B(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_154),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_149),
.B2(n_150),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_150),
.C(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_157),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_159),
.A2(n_165),
.B1(n_166),
.B2(n_290),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_159),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_162),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_172),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_167),
.B(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_170),
.B(n_172),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_171),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_181),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_180),
.C(n_181),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_178),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_190),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_187),
.C(n_190),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g306 ( 
.A1(n_192),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_193),
.B(n_194),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_196),
.B(n_197),
.C(n_202),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_198),
.B(n_200),
.C(n_201),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_286),
.B(n_291),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_272),
.B(n_285),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_248),
.B(n_271),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_228),
.B(n_247),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_218),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_208),
.B(n_218),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_214),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_210),
.B1(n_214),
.B2(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_225),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_223),
.C(n_225),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_224),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_226),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_235),
.B(n_246),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_234),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_240),
.B(n_245),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_237),
.B(n_239),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_249),
.B(n_250),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_261),
.B1(n_269),
.B2(n_270),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_251)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_256),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_260),
.C(n_270),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_258),
.Y(n_282)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_267),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_267),
.Y(n_280)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_273),
.B(n_274),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_281),
.C(n_283),
.Y(n_287)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_280),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_281),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_297),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_297),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.C(n_296),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_295),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_294),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_301),
.A2(n_306),
.B(n_309),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_303),
.Y(n_309)
);


endmodule