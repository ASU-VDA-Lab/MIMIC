module fake_jpeg_20861_n_179 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_127;
wire n_76;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_4),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

INVx11_ASAP7_75t_SL g73 ( 
.A(n_14),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_7),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_0),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_75),
.Y(n_93)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_95),
.Y(n_103)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_100),
.Y(n_109)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_60),
.Y(n_125)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_110),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_73),
.B(n_51),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_67),
.B(n_57),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_114),
.B(n_70),
.CI(n_59),
.CON(n_116),
.SN(n_116)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_66),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_81),
.B(n_68),
.C(n_64),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_131),
.B(n_55),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_126),
.B(n_56),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_52),
.B1(n_54),
.B2(n_62),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_80),
.B1(n_76),
.B2(n_69),
.Y(n_136)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_53),
.B1(n_65),
.B2(n_74),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_129),
.A2(n_69),
.B1(n_56),
.B2(n_2),
.Y(n_137)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_137),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_130),
.B1(n_115),
.B2(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_139),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_79),
.C(n_61),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_141),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_77),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_28),
.B(n_50),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_144),
.A2(n_146),
.B(n_134),
.C(n_138),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_1),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_157),
.B1(n_8),
.B2(n_17),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_18),
.C(n_19),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_135),
.A2(n_123),
.B1(n_3),
.B2(n_4),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_142),
.B1(n_6),
.B2(n_7),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_160),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_149),
.A2(n_142),
.B1(n_10),
.B2(n_12),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_162),
.C(n_163),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_156),
.C(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_160),
.C(n_153),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_149),
.B(n_164),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_148),
.Y(n_169)
);

AND2x4_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_165),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_22),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_48),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_25),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_42),
.Y(n_175)
);

AOI21x1_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_27),
.B(n_29),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_32),
.C(n_34),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_35),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_36),
.Y(n_179)
);


endmodule