module real_aes_1216_n_15 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_15);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_15;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_51;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_27;
wire n_23;
wire n_38;
wire n_50;
wire n_29;
wire n_20;
wire n_52;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
CKINVDCx20_ASAP7_75t_R g28 ( .A(n_0), .Y(n_28) );
NOR3xp33_ASAP7_75t_SL g26 ( .A(n_1), .B(n_6), .C(n_27), .Y(n_26) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_2), .Y(n_27) );
BUFx2_ASAP7_75t_L g52 ( .A(n_3), .Y(n_52) );
NAND3xp33_ASAP7_75t_SL g19 ( .A(n_4), .B(n_20), .C(n_21), .Y(n_19) );
NOR2xp33_ASAP7_75t_R g42 ( .A(n_4), .B(n_25), .Y(n_42) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_5), .Y(n_22) );
NOR2xp33_ASAP7_75t_R g48 ( .A(n_5), .B(n_9), .Y(n_48) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_7), .Y(n_30) );
CKINVDCx20_ASAP7_75t_R g20 ( .A(n_8), .Y(n_20) );
NOR2xp33_ASAP7_75t_R g46 ( .A(n_8), .B(n_47), .Y(n_46) );
CKINVDCx20_ASAP7_75t_R g29 ( .A(n_9), .Y(n_29) );
NAND2xp33_ASAP7_75t_SL g31 ( .A(n_9), .B(n_18), .Y(n_31) );
AOI322xp5_ASAP7_75t_SL g32 ( .A1(n_9), .A2(n_10), .A3(n_11), .B1(n_33), .B2(n_37), .C1(n_38), .C2(n_49), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g37 ( .A(n_9), .B(n_34), .Y(n_37) );
NAND2xp33_ASAP7_75t_SL g23 ( .A(n_12), .B(n_24), .Y(n_23) );
CKINVDCx20_ASAP7_75t_R g36 ( .A(n_12), .Y(n_36) );
NOR2xp33_ASAP7_75t_R g21 ( .A(n_13), .B(n_22), .Y(n_21) );
CKINVDCx20_ASAP7_75t_R g44 ( .A(n_13), .Y(n_44) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_14), .Y(n_16) );
OAI221xp5_ASAP7_75t_R g15 ( .A1(n_16), .A2(n_17), .B1(n_30), .B2(n_31), .C(n_32), .Y(n_15) );
NAND2xp33_ASAP7_75t_SL g17 ( .A(n_18), .B(n_29), .Y(n_17) );
NOR2xp33_ASAP7_75t_R g18 ( .A(n_19), .B(n_23), .Y(n_18) );
OR2x2_ASAP7_75t_L g34 ( .A(n_19), .B(n_35), .Y(n_34) );
NAND2xp33_ASAP7_75t_SL g35 ( .A(n_24), .B(n_36), .Y(n_35) );
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_25), .Y(n_24) );
NAND2xp33_ASAP7_75t_SL g25 ( .A(n_26), .B(n_28), .Y(n_25) );
CKINVDCx20_ASAP7_75t_R g33 ( .A(n_34), .Y(n_33) );
NAND2xp33_ASAP7_75t_SL g41 ( .A(n_36), .B(n_42), .Y(n_41) );
CKINVDCx20_ASAP7_75t_R g38 ( .A(n_39), .Y(n_38) );
NAND2xp33_ASAP7_75t_SL g39 ( .A(n_40), .B(n_43), .Y(n_39) );
CKINVDCx20_ASAP7_75t_R g40 ( .A(n_41), .Y(n_40) );
NOR2xp33_ASAP7_75t_R g43 ( .A(n_44), .B(n_45), .Y(n_43) );
CKINVDCx20_ASAP7_75t_R g45 ( .A(n_46), .Y(n_45) );
CKINVDCx14_ASAP7_75t_R g47 ( .A(n_48), .Y(n_47) );
CKINVDCx11_ASAP7_75t_R g49 ( .A(n_50), .Y(n_49) );
CKINVDCx20_ASAP7_75t_R g50 ( .A(n_51), .Y(n_50) );
HB1xp67_ASAP7_75t_L g51 ( .A(n_52), .Y(n_51) );
endmodule