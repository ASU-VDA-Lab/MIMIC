module fake_aes_9543_n_655 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_655);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_655;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g75 ( .A(n_52), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_59), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_55), .Y(n_77) );
BUFx3_ASAP7_75t_L g78 ( .A(n_60), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_37), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_61), .Y(n_80) );
INVx2_ASAP7_75t_SL g81 ( .A(n_5), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_26), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_72), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_62), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_15), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_46), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_36), .Y(n_87) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_14), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_5), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_1), .Y(n_90) );
BUFx2_ASAP7_75t_SL g91 ( .A(n_19), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_35), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_41), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_10), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_64), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_9), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_65), .Y(n_97) );
INVx1_ASAP7_75t_SL g98 ( .A(n_8), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_53), .Y(n_99) );
INVxp33_ASAP7_75t_L g100 ( .A(n_34), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_48), .Y(n_101) );
INVx2_ASAP7_75t_SL g102 ( .A(n_40), .Y(n_102) );
CKINVDCx14_ASAP7_75t_R g103 ( .A(n_31), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_28), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_25), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_69), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_27), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_3), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_50), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_70), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_30), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_1), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_7), .Y(n_114) );
INVxp33_ASAP7_75t_L g115 ( .A(n_16), .Y(n_115) );
NOR2xp67_ASAP7_75t_L g116 ( .A(n_73), .B(n_17), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_54), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_32), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_12), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_13), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_109), .B(n_0), .Y(n_121) );
AND2x6_ASAP7_75t_L g122 ( .A(n_78), .B(n_29), .Y(n_122) );
NOR2x1_ASAP7_75t_L g123 ( .A(n_109), .B(n_33), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_113), .Y(n_124) );
BUFx3_ASAP7_75t_L g125 ( .A(n_78), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_113), .B(n_0), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_113), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_81), .B(n_2), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_79), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_100), .B(n_115), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_76), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_78), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_81), .B(n_3), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_105), .Y(n_135) );
OAI22x1_ASAP7_75t_L g136 ( .A1(n_89), .A2(n_4), .B1(n_6), .B2(n_7), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_76), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_83), .Y(n_139) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_82), .A2(n_39), .B(n_71), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_108), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_120), .B(n_4), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_105), .Y(n_145) );
AOI22xp5_ASAP7_75t_L g146 ( .A1(n_89), .A2(n_6), .B1(n_8), .B2(n_9), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_112), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_112), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_102), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g150 ( .A1(n_94), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_118), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_118), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_88), .Y(n_153) );
BUFx2_ASAP7_75t_L g154 ( .A(n_90), .Y(n_154) );
INVx5_ASAP7_75t_L g155 ( .A(n_102), .Y(n_155) );
OAI22xp5_ASAP7_75t_SL g156 ( .A1(n_94), .A2(n_11), .B1(n_13), .B2(n_14), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_82), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_108), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_88), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_85), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_131), .B(n_103), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_124), .B(n_120), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_131), .B(n_96), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_154), .Y(n_164) );
INVx6_ASAP7_75t_L g165 ( .A(n_155), .Y(n_165) );
NAND3xp33_ASAP7_75t_L g166 ( .A(n_121), .B(n_119), .C(n_88), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_155), .Y(n_167) );
OR2x2_ASAP7_75t_L g168 ( .A(n_154), .B(n_98), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_143), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_143), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_133), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_127), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_133), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_132), .B(n_114), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
OR2x2_ASAP7_75t_L g176 ( .A(n_132), .B(n_119), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_155), .B(n_117), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_133), .Y(n_178) );
AND2x2_ASAP7_75t_SL g179 ( .A(n_143), .B(n_117), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_137), .B(n_75), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_155), .B(n_95), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_137), .B(n_114), .Y(n_184) );
INVx1_ASAP7_75t_SL g185 ( .A(n_126), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_122), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_126), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_155), .B(n_95), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_125), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_122), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_149), .B(n_85), .Y(n_191) );
INVx1_ASAP7_75t_SL g192 ( .A(n_126), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_160), .B(n_77), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_127), .Y(n_194) );
BUFx8_ASAP7_75t_SL g195 ( .A(n_129), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_122), .Y(n_196) );
NAND2xp33_ASAP7_75t_SL g197 ( .A(n_136), .B(n_88), .Y(n_197) );
INVx8_ASAP7_75t_L g198 ( .A(n_122), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_149), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_160), .B(n_80), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_128), .Y(n_201) );
NAND2x1p5_ASAP7_75t_L g202 ( .A(n_123), .B(n_99), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_125), .Y(n_203) );
INVxp67_ASAP7_75t_SL g204 ( .A(n_157), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_134), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_135), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_157), .B(n_92), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_122), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_128), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_130), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_122), .A2(n_111), .B1(n_88), .B2(n_91), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_141), .B(n_101), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_135), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_130), .Y(n_214) );
BUFx10_ASAP7_75t_L g215 ( .A(n_135), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_205), .B(n_141), .Y(n_216) );
OR2x2_ASAP7_75t_L g217 ( .A(n_168), .B(n_164), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_169), .A2(n_138), .B(n_139), .C(n_142), .Y(n_218) );
INVxp67_ASAP7_75t_L g219 ( .A(n_168), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_203), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_179), .A2(n_156), .B1(n_150), .B2(n_146), .Y(n_221) );
AND2x6_ASAP7_75t_SL g222 ( .A(n_163), .B(n_136), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_179), .A2(n_138), .B1(n_139), .B2(n_142), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_203), .Y(n_224) );
NAND3xp33_ASAP7_75t_L g225 ( .A(n_211), .B(n_135), .C(n_152), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_186), .B(n_93), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_182), .B(n_141), .Y(n_227) );
CKINVDCx11_ASAP7_75t_R g228 ( .A(n_162), .Y(n_228) );
BUFx8_ASAP7_75t_L g229 ( .A(n_162), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_161), .B(n_158), .Y(n_230) );
BUFx12f_ASAP7_75t_L g231 ( .A(n_164), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_204), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_199), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_162), .A2(n_111), .B1(n_144), .B2(n_147), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_161), .B(n_158), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_200), .B(n_158), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_215), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_185), .B(n_104), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_215), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_186), .B(n_110), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_197), .A2(n_144), .B1(n_148), .B2(n_147), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_174), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_193), .B(n_148), .Y(n_243) );
OR2x6_ASAP7_75t_L g244 ( .A(n_198), .B(n_91), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_174), .Y(n_245) );
INVxp67_ASAP7_75t_L g246 ( .A(n_207), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_192), .B(n_86), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_176), .B(n_86), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_184), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_195), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_170), .B(n_87), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_176), .B(n_184), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_215), .Y(n_253) );
BUFx4f_ASAP7_75t_L g254 ( .A(n_202), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_189), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_209), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_212), .B(n_87), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_197), .A2(n_152), .B1(n_151), .B2(n_145), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_187), .B(n_97), .Y(n_259) );
OR2x2_ASAP7_75t_SL g260 ( .A(n_195), .B(n_140), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_187), .B(n_97), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_214), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_186), .B(n_99), .Y(n_263) );
NOR2x2_ASAP7_75t_L g264 ( .A(n_202), .B(n_140), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_190), .Y(n_265) );
INVx8_ASAP7_75t_L g266 ( .A(n_198), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_187), .A2(n_145), .B1(n_151), .B2(n_152), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_209), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_202), .B(n_106), .Y(n_269) );
INVxp67_ASAP7_75t_L g270 ( .A(n_210), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_190), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_189), .B(n_106), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_213), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_191), .B(n_107), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_219), .A2(n_166), .B1(n_198), .B2(n_194), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_263), .A2(n_208), .B(n_198), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_262), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_219), .B(n_196), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_252), .B(n_210), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_246), .B(n_201), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_217), .B(n_201), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_223), .A2(n_196), .B1(n_172), .B2(n_194), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_265), .B(n_190), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_259), .A2(n_208), .B(n_167), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_246), .B(n_201), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_266), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_261), .A2(n_167), .B(n_172), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_270), .A2(n_177), .B(n_188), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_273), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_266), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_242), .A2(n_183), .B1(n_107), .B2(n_145), .C(n_151), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_270), .A2(n_140), .B(n_178), .Y(n_292) );
NAND3xp33_ASAP7_75t_SL g293 ( .A(n_250), .B(n_213), .C(n_206), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_226), .A2(n_140), .B(n_178), .Y(n_294) );
INVx4_ASAP7_75t_L g295 ( .A(n_228), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_245), .B(n_116), .Y(n_296) );
NOR3xp33_ASAP7_75t_SL g297 ( .A(n_227), .B(n_116), .C(n_20), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_240), .A2(n_171), .B(n_180), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_223), .B(n_213), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_229), .Y(n_300) );
BUFx4f_ASAP7_75t_SL g301 ( .A(n_231), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_249), .A2(n_145), .B1(n_151), .B2(n_152), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_SL g303 ( .A1(n_218), .A2(n_180), .B(n_175), .C(n_173), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_229), .B(n_165), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_254), .B(n_165), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g306 ( .A1(n_216), .A2(n_175), .B(n_173), .C(n_171), .Y(n_306) );
AO22x1_ASAP7_75t_L g307 ( .A1(n_254), .A2(n_152), .B1(n_151), .B2(n_145), .Y(n_307) );
INVx5_ASAP7_75t_L g308 ( .A(n_244), .Y(n_308) );
AO21x2_ASAP7_75t_L g309 ( .A1(n_269), .A2(n_206), .B(n_181), .Y(n_309) );
NOR2xp33_ASAP7_75t_SL g310 ( .A(n_266), .B(n_181), .Y(n_310) );
NAND2x1_ASAP7_75t_L g311 ( .A(n_244), .B(n_165), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_256), .B(n_165), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_265), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_232), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_233), .Y(n_315) );
OAI21xp5_ASAP7_75t_L g316 ( .A1(n_225), .A2(n_159), .B(n_153), .Y(n_316) );
OR2x6_ASAP7_75t_L g317 ( .A(n_244), .B(n_159), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_230), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_235), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_265), .B(n_159), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_278), .A2(n_221), .B1(n_238), .B2(n_234), .Y(n_321) );
OAI22xp33_ASAP7_75t_L g322 ( .A1(n_295), .A2(n_248), .B1(n_247), .B2(n_236), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_318), .B(n_251), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_284), .A2(n_257), .B(n_265), .Y(n_324) );
AOI31xp67_ASAP7_75t_L g325 ( .A1(n_320), .A2(n_264), .A3(n_260), .B(n_255), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_294), .A2(n_271), .B(n_268), .Y(n_326) );
AO31x2_ASAP7_75t_L g327 ( .A1(n_292), .A2(n_272), .A3(n_251), .B(n_274), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_300), .Y(n_328) );
OAI22xp5_ASAP7_75t_SL g329 ( .A1(n_295), .A2(n_241), .B1(n_222), .B2(n_258), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_288), .A2(n_271), .B(n_272), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_319), .B(n_227), .Y(n_331) );
OAI21x1_ASAP7_75t_L g332 ( .A1(n_316), .A2(n_267), .B(n_220), .Y(n_332) );
A2O1A1Ixp33_ASAP7_75t_L g333 ( .A1(n_297), .A2(n_287), .B(n_315), .C(n_243), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_281), .B(n_241), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_279), .A2(n_224), .B1(n_253), .B2(n_239), .Y(n_335) );
NOR2xp67_ASAP7_75t_SL g336 ( .A(n_308), .B(n_237), .Y(n_336) );
OAI21xp5_ASAP7_75t_L g337 ( .A1(n_299), .A2(n_267), .B(n_258), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_286), .Y(n_338) );
NAND3xp33_ASAP7_75t_L g339 ( .A(n_302), .B(n_153), .C(n_159), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_303), .A2(n_159), .B(n_153), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_286), .Y(n_341) );
AOI22xp33_ASAP7_75t_SL g342 ( .A1(n_308), .A2(n_153), .B1(n_21), .B2(n_22), .Y(n_342) );
INVx5_ASAP7_75t_SL g343 ( .A(n_286), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_280), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_282), .A2(n_153), .B(n_23), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_282), .A2(n_18), .B(n_24), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_285), .B(n_38), .Y(n_347) );
O2A1O1Ixp5_ASAP7_75t_L g348 ( .A1(n_311), .A2(n_42), .B(n_43), .C(n_44), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_314), .B(n_45), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_SL g350 ( .A1(n_293), .A2(n_47), .B(n_49), .C(n_51), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_333), .A2(n_306), .B(n_298), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_338), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_321), .B(n_296), .Y(n_353) );
OAI21xp5_ASAP7_75t_L g354 ( .A1(n_330), .A2(n_316), .B(n_312), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_338), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_326), .A2(n_317), .B(n_312), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_327), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_344), .B(n_277), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_323), .B(n_296), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_327), .Y(n_360) );
A2O1A1Ixp33_ASAP7_75t_L g361 ( .A1(n_331), .A2(n_291), .B(n_308), .C(n_305), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_349), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_329), .A2(n_317), .B1(n_301), .B2(n_304), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_328), .Y(n_364) );
A2O1A1Ixp33_ASAP7_75t_L g365 ( .A1(n_346), .A2(n_275), .B(n_289), .C(n_276), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_322), .B(n_290), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_334), .B(n_290), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_327), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_347), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_343), .B(n_290), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_343), .B(n_309), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_341), .B(n_309), .Y(n_372) );
AO21x2_ASAP7_75t_L g373 ( .A1(n_340), .A2(n_283), .B(n_307), .Y(n_373) );
AO21x2_ASAP7_75t_L g374 ( .A1(n_345), .A2(n_313), .B(n_310), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_348), .A2(n_310), .B(n_313), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_341), .B(n_317), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_353), .B(n_329), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_359), .B(n_338), .Y(n_378) );
AO21x2_ASAP7_75t_L g379 ( .A1(n_368), .A2(n_350), .B(n_337), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_357), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_359), .B(n_332), .Y(n_381) );
OAI211xp5_ASAP7_75t_L g382 ( .A1(n_363), .A2(n_342), .B(n_324), .C(n_339), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_357), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_357), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_360), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_360), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_368), .B(n_313), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_360), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_367), .B(n_336), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_364), .B(n_335), .Y(n_390) );
OA21x2_ASAP7_75t_L g391 ( .A1(n_375), .A2(n_339), .B(n_325), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_358), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_372), .Y(n_393) );
AO21x2_ASAP7_75t_L g394 ( .A1(n_351), .A2(n_56), .B(n_57), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_358), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_371), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_362), .B(n_58), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_362), .B(n_63), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_371), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_364), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_352), .Y(n_401) );
AO21x1_ASAP7_75t_SL g402 ( .A1(n_366), .A2(n_66), .B(n_67), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_352), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_352), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_352), .Y(n_405) );
OA21x2_ASAP7_75t_L g406 ( .A1(n_375), .A2(n_68), .B(n_74), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_369), .B(n_354), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_376), .B(n_355), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_352), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_396), .B(n_355), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_393), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_392), .B(n_369), .Y(n_412) );
OR2x6_ASAP7_75t_L g413 ( .A(n_386), .B(n_356), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_400), .B(n_370), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_381), .B(n_355), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_395), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_380), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_377), .B(n_361), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_381), .B(n_354), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_380), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_393), .Y(n_422) );
BUFx3_ASAP7_75t_L g423 ( .A(n_380), .Y(n_423) );
BUFx3_ASAP7_75t_L g424 ( .A(n_383), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_383), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_383), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_384), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_377), .B(n_376), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_384), .Y(n_429) );
INVx5_ASAP7_75t_SL g430 ( .A(n_394), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_378), .B(n_365), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_396), .B(n_374), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_378), .B(n_373), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_399), .B(n_374), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_399), .B(n_374), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_387), .B(n_373), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_384), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_385), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_385), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_387), .B(n_373), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_385), .Y(n_441) );
INVx5_ASAP7_75t_SL g442 ( .A(n_394), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_388), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_407), .B(n_388), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_388), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_407), .Y(n_446) );
INVx2_ASAP7_75t_SL g447 ( .A(n_408), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_404), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_390), .B(n_389), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_408), .B(n_405), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_404), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_405), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_389), .B(n_398), .Y(n_453) );
INVx4_ASAP7_75t_L g454 ( .A(n_401), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_401), .B(n_409), .Y(n_455) );
NAND4xp25_ASAP7_75t_SL g456 ( .A(n_382), .B(n_398), .C(n_397), .D(n_402), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_453), .A2(n_397), .B1(n_382), .B2(n_409), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_419), .B(n_379), .Y(n_458) );
AND2x4_ASAP7_75t_SL g459 ( .A(n_415), .B(n_409), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_419), .B(n_379), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_436), .B(n_379), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_411), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_416), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_411), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_436), .B(n_379), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_440), .B(n_401), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_412), .B(n_403), .Y(n_467) );
NAND2x1_ASAP7_75t_L g468 ( .A(n_441), .B(n_406), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_415), .B(n_403), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_440), .B(n_403), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_422), .B(n_394), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_422), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_448), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_432), .B(n_434), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_448), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_447), .B(n_394), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_432), .B(n_391), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_425), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_447), .B(n_391), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_425), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_421), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_441), .Y(n_482) );
INVx3_ASAP7_75t_L g483 ( .A(n_423), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_451), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_434), .B(n_391), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_421), .Y(n_486) );
NAND2xp33_ASAP7_75t_R g487 ( .A(n_449), .B(n_406), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_435), .B(n_391), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_441), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_423), .Y(n_490) );
AND2x4_ASAP7_75t_SL g491 ( .A(n_450), .B(n_402), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_429), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_435), .B(n_406), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_423), .B(n_406), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_441), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_428), .B(n_450), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_424), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_418), .B(n_446), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_424), .B(n_426), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_417), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_451), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_444), .B(n_433), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_417), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_444), .B(n_446), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_424), .B(n_426), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_429), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_414), .B(n_410), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_452), .B(n_454), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_420), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_439), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_439), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_443), .B(n_445), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_463), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_496), .B(n_443), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_474), .B(n_455), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_502), .B(n_445), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_474), .B(n_455), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_466), .B(n_426), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_466), .B(n_437), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_498), .B(n_452), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_457), .A2(n_456), .B1(n_431), .B2(n_410), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_462), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_508), .B(n_413), .Y(n_523) );
NOR2xp33_ASAP7_75t_SL g524 ( .A(n_491), .B(n_454), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_462), .Y(n_525) );
INVxp67_ASAP7_75t_SL g526 ( .A(n_497), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_508), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_486), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_491), .A2(n_454), .B1(n_413), .B2(n_427), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_502), .B(n_437), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_459), .B(n_454), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_504), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_470), .B(n_420), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_504), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_473), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_507), .B(n_427), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_459), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_475), .Y(n_538) );
INVxp67_ASAP7_75t_SL g539 ( .A(n_490), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_470), .B(n_438), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_484), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_512), .B(n_438), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_477), .B(n_413), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_458), .A2(n_413), .B1(n_430), .B2(n_442), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_512), .B(n_413), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_500), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_508), .B(n_430), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_477), .B(n_430), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_485), .B(n_430), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_481), .B(n_442), .Y(n_550) );
INVxp67_ASAP7_75t_SL g551 ( .A(n_490), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_464), .B(n_442), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_472), .B(n_442), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_501), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_467), .B(n_458), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_481), .B(n_460), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_500), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g558 ( .A(n_487), .B(n_471), .C(n_476), .Y(n_558) );
BUFx2_ASAP7_75t_L g559 ( .A(n_483), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_485), .B(n_488), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_499), .Y(n_561) );
NOR2xp67_ASAP7_75t_L g562 ( .A(n_483), .B(n_479), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_517), .B(n_488), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_532), .B(n_461), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_536), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_534), .B(n_461), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_513), .B(n_465), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_516), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_527), .Y(n_569) );
XNOR2x1_ASAP7_75t_L g570 ( .A(n_521), .B(n_469), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_535), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_556), .A2(n_465), .B1(n_511), .B2(n_510), .C(n_506), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_546), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_517), .B(n_469), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_515), .B(n_469), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_560), .B(n_460), .Y(n_576) );
XOR2x2_ASAP7_75t_L g577 ( .A(n_537), .B(n_505), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_555), .B(n_511), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_561), .B(n_505), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_556), .B(n_510), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_528), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_538), .Y(n_582) );
AOI32xp33_ASAP7_75t_L g583 ( .A1(n_524), .A2(n_543), .A3(n_526), .B1(n_539), .B2(n_551), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_528), .B(n_478), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_543), .B(n_499), .Y(n_585) );
INVxp33_ASAP7_75t_L g586 ( .A(n_562), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_558), .A2(n_492), .B1(n_478), .B2(n_480), .C(n_506), .Y(n_587) );
OAI32xp33_ASAP7_75t_L g588 ( .A1(n_545), .A2(n_514), .A3(n_547), .B1(n_530), .B2(n_550), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_541), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_529), .B(n_483), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_520), .B(n_480), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_546), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_519), .B(n_492), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_519), .B(n_493), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_518), .B(n_493), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_559), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_554), .Y(n_597) );
CKINVDCx14_ASAP7_75t_R g598 ( .A(n_577), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_584), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_563), .B(n_549), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_573), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_573), .Y(n_602) );
OAI222xp33_ASAP7_75t_L g603 ( .A1(n_583), .A2(n_544), .B1(n_523), .B2(n_549), .C1(n_548), .C2(n_531), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_572), .B(n_540), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_577), .Y(n_605) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_581), .Y(n_606) );
OAI21xp33_ASAP7_75t_L g607 ( .A1(n_586), .A2(n_548), .B(n_544), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_569), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_597), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_569), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_587), .B(n_540), .Y(n_611) );
INVx2_ASAP7_75t_SL g612 ( .A(n_574), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_570), .A2(n_523), .B1(n_518), .B2(n_547), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_568), .B(n_522), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_571), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_575), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_576), .B(n_542), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_592), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_563), .B(n_533), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_598), .A2(n_570), .B1(n_565), .B2(n_591), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_611), .B(n_591), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_606), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_605), .B(n_586), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_617), .Y(n_624) );
NAND2x1_ASAP7_75t_L g625 ( .A(n_600), .B(n_619), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_604), .B(n_580), .Y(n_626) );
OR3x1_ASAP7_75t_L g627 ( .A(n_598), .B(n_588), .C(n_550), .Y(n_627) );
A2O1A1Ixp33_ASAP7_75t_L g628 ( .A1(n_607), .A2(n_596), .B(n_590), .C(n_523), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_613), .A2(n_590), .B1(n_567), .B2(n_566), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_603), .A2(n_589), .B1(n_582), .B2(n_564), .C(n_593), .Y(n_630) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_608), .A2(n_578), .B(n_594), .C(n_552), .Y(n_631) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_610), .A2(n_553), .B(n_525), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_624), .Y(n_633) );
NAND3xp33_ASAP7_75t_SL g634 ( .A(n_630), .B(n_616), .C(n_600), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g635 ( .A1(n_623), .A2(n_599), .B(n_614), .C(n_615), .Y(n_635) );
NOR4xp25_ASAP7_75t_L g636 ( .A(n_628), .B(n_609), .C(n_612), .D(n_619), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_620), .A2(n_612), .B1(n_579), .B2(n_585), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_625), .A2(n_617), .B(n_602), .C(n_618), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_627), .A2(n_602), .B1(n_595), .B2(n_601), .C(n_618), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_621), .A2(n_585), .B1(n_595), .B2(n_601), .Y(n_640) );
NOR5xp2_ASAP7_75t_L g641 ( .A(n_638), .B(n_622), .C(n_631), .D(n_632), .E(n_629), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_633), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_634), .B(n_626), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_636), .B(n_592), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_642), .Y(n_645) );
NOR3xp33_ASAP7_75t_L g646 ( .A(n_643), .B(n_639), .C(n_635), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_644), .B(n_637), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_646), .B(n_641), .C(n_640), .Y(n_648) );
INVxp33_ASAP7_75t_SL g649 ( .A(n_645), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_648), .A2(n_647), .B1(n_533), .B2(n_468), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_650), .A2(n_649), .B1(n_557), .B2(n_489), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_651), .A2(n_557), .B1(n_468), .B2(n_494), .C(n_489), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_652), .A2(n_482), .B(n_495), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_653), .A2(n_494), .B1(n_482), .B2(n_495), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_654), .A2(n_503), .B1(n_509), .B2(n_649), .C(n_648), .Y(n_655) );
endmodule