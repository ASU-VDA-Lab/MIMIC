module fake_ariane_1598_n_241 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_32, n_28, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_241);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_32;
input n_28;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_241;

wire n_83;
wire n_233;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_124;
wire n_119;
wire n_167;
wire n_90;
wire n_195;
wire n_38;
wire n_213;
wire n_47;
wire n_110;
wire n_153;
wire n_221;
wire n_197;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_237;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_236;
wire n_205;
wire n_71;
wire n_109;
wire n_208;
wire n_96;
wire n_156;
wire n_209;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_210;
wire n_147;
wire n_204;
wire n_225;
wire n_235;
wire n_200;
wire n_51;
wire n_166;
wire n_76;
wire n_218;
wire n_103;
wire n_79;
wire n_226;
wire n_46;
wire n_220;
wire n_84;
wire n_199;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_224;
wire n_44;
wire n_240;
wire n_82;
wire n_178;
wire n_217;
wire n_42;
wire n_57;
wire n_131;
wire n_201;
wire n_229;
wire n_70;
wire n_222;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_214;
wire n_227;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_188;
wire n_185;
wire n_58;
wire n_37;
wire n_65;
wire n_123;
wire n_212;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_198;
wire n_148;
wire n_232;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_228;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_206;
wire n_207;
wire n_238;
wire n_41;
wire n_219;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_231;
wire n_192;
wire n_80;
wire n_146;
wire n_234;
wire n_230;
wire n_211;
wire n_194;
wire n_97;
wire n_154;
wire n_215;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_78;
wire n_193;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_216;
wire n_155;
wire n_127;
wire n_239;
wire n_223;
wire n_54;

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_0),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_7),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_17),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

AND2x4_ASAP7_75t_L g90 ( 
.A(n_37),
.B(n_18),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_19),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_62),
.B(n_24),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_48),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_67),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_83),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_47),
.B1(n_61),
.B2(n_56),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_56),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_86),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_64),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_61),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_32),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_94),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_73),
.B(n_87),
.C(n_81),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_87),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_79),
.A2(n_84),
.B(n_82),
.C(n_80),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_88),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_94),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

NOR2xp67_ASAP7_75t_L g132 ( 
.A(n_76),
.B(n_97),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_134),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_93),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_99),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_111),
.B(n_103),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_107),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_112),
.A2(n_125),
.B1(n_115),
.B2(n_122),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_113),
.Y(n_148)
);

AND3x1_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_110),
.C(n_126),
.Y(n_149)
);

AND3x1_ASAP7_75t_SL g150 ( 
.A(n_119),
.B(n_131),
.C(n_128),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_132),
.Y(n_151)
);

BUFx4f_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

NOR2x1p5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_145),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_136),
.B1(n_148),
.B2(n_149),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_155),
.C(n_154),
.Y(n_166)
);

NOR2xp67_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_161),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_144),
.B(n_156),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

OR2x6_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_161),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_147),
.Y(n_172)
);

NAND2x1p5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_151),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

AND2x4_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_158),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_129),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_136),
.A2(n_137),
.B(n_145),
.C(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_146),
.A2(n_111),
.B1(n_112),
.B2(n_136),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_164),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

OAI221xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_163),
.B1(n_165),
.B2(n_178),
.C(n_183),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_163),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_187),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_204),
.Y(n_211)
);

AND2x4_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_174),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_183),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_196),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_173),
.Y(n_217)
);

OAI211xp5_ASAP7_75t_SL g218 ( 
.A1(n_201),
.A2(n_184),
.B(n_176),
.C(n_167),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_192),
.B1(n_191),
.B2(n_203),
.Y(n_221)
);

AO21x2_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_202),
.B(n_200),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_189),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_216),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_216),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_210),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_220),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_227),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

AND3x1_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_226),
.C(n_213),
.Y(n_232)
);

NOR3xp33_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_218),
.C(n_229),
.Y(n_233)
);

NAND4xp75_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_232),
.C(n_226),
.D(n_231),
.Y(n_234)
);

O2A1O1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_215),
.B(n_203),
.C(n_173),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_235),
.Y(n_236)
);

AOI221xp5_ASAP7_75t_L g237 ( 
.A1(n_236),
.A2(n_221),
.B1(n_194),
.B2(n_222),
.C(n_206),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_237),
.A2(n_222),
.B1(n_197),
.B2(n_192),
.Y(n_238)
);

AOI222xp33_ASAP7_75t_L g239 ( 
.A1(n_238),
.A2(n_189),
.B1(n_212),
.B2(n_205),
.C1(n_208),
.C2(n_214),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_212),
.Y(n_240)
);

AOI221xp5_ASAP7_75t_L g241 ( 
.A1(n_240),
.A2(n_217),
.B1(n_211),
.B2(n_214),
.C(n_171),
.Y(n_241)
);


endmodule