module fake_jpeg_25648_n_37 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_0),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_19),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_18),
.B1(n_7),
.B2(n_8),
.Y(n_20)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_4),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_22),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_18),
.A2(n_16),
.B1(n_8),
.B2(n_17),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_18),
.C(n_16),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_22),
.B1(n_24),
.B2(n_8),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_17),
.B1(n_14),
.B2(n_26),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_12),
.B(n_9),
.C(n_13),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_15),
.B(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_33),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_9),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_29),
.A3(n_9),
.B1(n_13),
.B2(n_10),
.C1(n_14),
.C2(n_3),
.Y(n_36)
);

AO221x1_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_3),
.B1(n_13),
.B2(n_34),
.C(n_31),
.Y(n_37)
);


endmodule