module real_jpeg_30422_n_21 (n_17, n_8, n_0, n_157, n_2, n_10, n_9, n_12, n_154, n_156, n_152, n_6, n_159, n_153, n_161, n_162, n_11, n_14, n_160, n_7, n_18, n_3, n_5, n_4, n_1, n_20, n_19, n_158, n_16, n_15, n_13, n_155, n_21);

input n_17;
input n_8;
input n_0;
input n_157;
input n_2;
input n_10;
input n_9;
input n_12;
input n_154;
input n_156;
input n_152;
input n_6;
input n_159;
input n_153;
input n_161;
input n_162;
input n_11;
input n_14;
input n_160;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_158;
input n_16;
input n_15;
input n_13;
input n_155;

output n_21;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_80;
wire n_30;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_0),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_0),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_1),
.B(n_88),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_2),
.B(n_24),
.Y(n_144)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_4),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_5),
.Y(n_105)
);

AOI221xp5_ASAP7_75t_L g85 ( 
.A1(n_6),
.A2(n_17),
.B1(n_86),
.B2(n_91),
.C(n_94),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_6),
.Y(n_96)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_7),
.B(n_41),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_8),
.B(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_9),
.A2(n_59),
.A3(n_61),
.B1(n_66),
.B2(n_127),
.C1(n_129),
.C2(n_162),
.Y(n_126)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_10),
.B(n_68),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_12),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_12),
.B(n_72),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_14),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_14),
.B(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_15),
.B(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_15),
.Y(n_142)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_17),
.B(n_86),
.C(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_18),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_19),
.A2(n_146),
.B1(n_147),
.B2(n_150),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_19),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_20),
.B(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_145),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_144),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_135),
.B(n_141),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_38),
.B(n_133),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_37),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_32),
.B(n_37),
.Y(n_134)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_36),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_48),
.B(n_132),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_47),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_46),
.Y(n_140)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI31xp67_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_77),
.A3(n_113),
.B(n_122),
.Y(n_49)
);

NOR3xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_65),
.C(n_71),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_51),
.A2(n_123),
.B(n_126),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_53),
.B(n_71),
.C(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_153),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_63),
.Y(n_84)
);

OA21x2_ASAP7_75t_SL g123 ( 
.A1(n_65),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_107),
.C(n_108),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_98),
.B(n_106),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_85),
.B1(n_96),
.B2(n_97),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_158),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_105),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_105),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_152),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_154),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_155),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_156),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_157),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_159),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_160),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_161),
.Y(n_116)
);


endmodule