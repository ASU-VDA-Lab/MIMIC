module real_aes_6159_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g464 ( .A1(n_0), .A2(n_165), .B(n_465), .C(n_468), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_1), .B(n_459), .Y(n_470) );
INVx1_ASAP7_75t_L g428 ( .A(n_2), .Y(n_428) );
INVx1_ASAP7_75t_L g214 ( .A(n_3), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_4), .B(n_153), .Y(n_493) );
XNOR2xp5_ASAP7_75t_SL g763 ( .A(n_5), .B(n_102), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_6), .A2(n_443), .B(n_513), .Y(n_512) );
OAI22xp5_ASAP7_75t_SL g758 ( .A1(n_7), .A2(n_10), .B1(n_423), .B2(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_7), .Y(n_759) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_8), .A2(n_170), .B(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g164 ( .A1(n_9), .A2(n_40), .B1(n_126), .B2(n_138), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g109 ( .A1(n_10), .A2(n_110), .B1(n_111), .B2(n_423), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_10), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_11), .B(n_170), .Y(n_203) );
AND2x6_ASAP7_75t_L g141 ( .A(n_12), .B(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_13), .A2(n_141), .B(n_446), .C(n_535), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_14), .B(n_41), .Y(n_429) );
INVx1_ASAP7_75t_L g122 ( .A(n_15), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_16), .B(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g208 ( .A(n_17), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_18), .B(n_153), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_19), .B(n_168), .Y(n_186) );
AO32x2_ASAP7_75t_L g162 ( .A1(n_20), .A2(n_163), .A3(n_167), .B1(n_169), .B2(n_170), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_21), .A2(n_59), .B1(n_732), .B2(n_733), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_21), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_22), .B(n_126), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_23), .B(n_168), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_24), .A2(n_57), .B1(n_126), .B2(n_138), .Y(n_166) );
AOI22xp33_ASAP7_75t_SL g179 ( .A1(n_25), .A2(n_84), .B1(n_126), .B2(n_130), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_26), .B(n_126), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_27), .A2(n_169), .B(n_446), .C(n_448), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_28), .Y(n_768) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_29), .A2(n_169), .B(n_446), .C(n_525), .Y(n_524) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_30), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_31), .B(n_118), .Y(n_228) );
AOI222xp33_ASAP7_75t_L g106 ( .A1(n_32), .A2(n_107), .B1(n_725), .B2(n_726), .C1(n_735), .C2(n_739), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_33), .A2(n_443), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_34), .B(n_118), .Y(n_160) );
INVx2_ASAP7_75t_L g128 ( .A(n_35), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_36), .A2(n_477), .B(n_478), .C(n_482), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_37), .B(n_126), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_38), .B(n_118), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_39), .B(n_133), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_42), .B(n_442), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_43), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_44), .B(n_153), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_45), .B(n_443), .Y(n_523) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_46), .A2(n_727), .B1(n_728), .B2(n_734), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_46), .Y(n_734) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_47), .A2(n_477), .B(n_482), .C(n_504), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_48), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_48), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_49), .B(n_126), .Y(n_196) );
INVx1_ASAP7_75t_L g466 ( .A(n_50), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_51), .A2(n_92), .B1(n_138), .B2(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g505 ( .A(n_52), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_53), .B(n_126), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_54), .B(n_126), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_55), .B(n_443), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_56), .B(n_201), .Y(n_200) );
AOI22xp33_ASAP7_75t_SL g190 ( .A1(n_58), .A2(n_63), .B1(n_126), .B2(n_130), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_59), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_60), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g125 ( .A(n_61), .B(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_62), .B(n_126), .Y(n_227) );
INVx1_ASAP7_75t_L g142 ( .A(n_64), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_65), .B(n_443), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_66), .B(n_459), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_67), .A2(n_201), .B(n_211), .C(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_68), .B(n_126), .Y(n_215) );
INVx1_ASAP7_75t_L g121 ( .A(n_69), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_70), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_71), .B(n_153), .Y(n_480) );
AO32x2_ASAP7_75t_L g175 ( .A1(n_72), .A2(n_169), .A3(n_170), .B1(n_176), .B2(n_180), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_73), .B(n_154), .Y(n_536) );
INVx1_ASAP7_75t_L g226 ( .A(n_74), .Y(n_226) );
INVx1_ASAP7_75t_L g151 ( .A(n_75), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_76), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_77), .B(n_450), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_78), .A2(n_446), .B(n_482), .C(n_491), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_79), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_79), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_80), .B(n_130), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_81), .Y(n_514) );
INVx1_ASAP7_75t_L g745 ( .A(n_82), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_83), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_85), .B(n_138), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_86), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_87), .B(n_130), .Y(n_157) );
INVx2_ASAP7_75t_L g119 ( .A(n_88), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_89), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_90), .B(n_140), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_91), .B(n_130), .Y(n_197) );
OR2x2_ASAP7_75t_L g426 ( .A(n_93), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g724 ( .A(n_93), .Y(n_724) );
OR2x2_ASAP7_75t_L g749 ( .A(n_93), .B(n_738), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_94), .A2(n_103), .B1(n_130), .B2(n_131), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_95), .B(n_443), .Y(n_475) );
INVx1_ASAP7_75t_L g479 ( .A(n_96), .Y(n_479) );
INVxp67_ASAP7_75t_L g517 ( .A(n_97), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_98), .B(n_130), .Y(n_224) );
INVx1_ASAP7_75t_L g492 ( .A(n_99), .Y(n_492) );
INVx1_ASAP7_75t_L g532 ( .A(n_100), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_101), .B(n_745), .Y(n_744) );
AOI222xp33_ASAP7_75t_L g104 ( .A1(n_102), .A2(n_105), .B1(n_741), .B2(n_750), .C1(n_771), .C2(n_777), .Y(n_104) );
AND2x2_ASAP7_75t_L g507 ( .A(n_102), .B(n_118), .Y(n_507) );
INVxp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22x1_ASAP7_75t_SL g107 ( .A1(n_108), .A2(n_424), .B1(n_430), .B2(n_721), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_109), .A2(n_431), .B1(n_721), .B2(n_740), .Y(n_739) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_110), .A2(n_111), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_345), .Y(n_111) );
NAND5xp2_ASAP7_75t_L g112 ( .A(n_113), .B(n_264), .C(n_279), .D(n_305), .E(n_327), .Y(n_112) );
NOR2xp33_ASAP7_75t_SL g113 ( .A(n_114), .B(n_244), .Y(n_113) );
OAI221xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_181), .B1(n_217), .B2(n_233), .C(n_234), .Y(n_114) );
NOR2xp33_ASAP7_75t_SL g115 ( .A(n_116), .B(n_171), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_116), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_SL g421 ( .A(n_116), .Y(n_421) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_144), .Y(n_116) );
INVx1_ASAP7_75t_L g261 ( .A(n_117), .Y(n_261) );
AND2x2_ASAP7_75t_L g263 ( .A(n_117), .B(n_162), .Y(n_263) );
AND2x2_ASAP7_75t_L g273 ( .A(n_117), .B(n_161), .Y(n_273) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_117), .Y(n_291) );
INVx1_ASAP7_75t_L g301 ( .A(n_117), .Y(n_301) );
OR2x2_ASAP7_75t_L g339 ( .A(n_117), .B(n_238), .Y(n_339) );
INVx2_ASAP7_75t_L g389 ( .A(n_117), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_117), .B(n_237), .Y(n_406) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_143), .Y(n_117) );
OA21x2_ASAP7_75t_L g147 ( .A1(n_118), .A2(n_148), .B(n_160), .Y(n_147) );
INVx2_ASAP7_75t_L g180 ( .A(n_118), .Y(n_180) );
INVx1_ASAP7_75t_L g456 ( .A(n_118), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_118), .A2(n_475), .B(n_476), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_118), .A2(n_502), .B(n_503), .Y(n_501) );
AND2x2_ASAP7_75t_SL g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x2_ASAP7_75t_L g168 ( .A(n_119), .B(n_120), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_135), .B(n_141), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B(n_132), .Y(n_124) );
INVx3_ASAP7_75t_L g150 ( .A(n_126), .Y(n_150) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_126), .Y(n_494) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g138 ( .A(n_127), .Y(n_138) );
BUFx3_ASAP7_75t_L g178 ( .A(n_127), .Y(n_178) );
AND2x6_ASAP7_75t_L g446 ( .A(n_127), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g131 ( .A(n_128), .Y(n_131) );
INVx1_ASAP7_75t_L g202 ( .A(n_128), .Y(n_202) );
INVx2_ASAP7_75t_L g209 ( .A(n_130), .Y(n_209) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
INVx3_ASAP7_75t_L g154 ( .A(n_134), .Y(n_154) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_134), .Y(n_159) );
AND2x2_ASAP7_75t_L g444 ( .A(n_134), .B(n_202), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_134), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B(n_139), .Y(n_135) );
O2A1O1Ixp5_ASAP7_75t_L g225 ( .A1(n_139), .A2(n_213), .B(n_226), .C(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g163 ( .A1(n_140), .A2(n_164), .B1(n_165), .B2(n_166), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g176 ( .A1(n_140), .A2(n_154), .B1(n_177), .B2(n_179), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g188 ( .A1(n_140), .A2(n_165), .B1(n_189), .B2(n_190), .Y(n_188) );
INVx4_ASAP7_75t_L g467 ( .A(n_140), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g148 ( .A1(n_141), .A2(n_149), .B(n_155), .Y(n_148) );
BUFx3_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_141), .A2(n_195), .B(n_198), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_141), .A2(n_207), .B(n_212), .Y(n_206) );
AND2x4_ASAP7_75t_L g443 ( .A(n_141), .B(n_444), .Y(n_443) );
INVx4_ASAP7_75t_SL g469 ( .A(n_141), .Y(n_469) );
NAND2x1p5_ASAP7_75t_L g533 ( .A(n_141), .B(n_444), .Y(n_533) );
NOR2xp67_ASAP7_75t_L g144 ( .A(n_145), .B(n_161), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_146), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_146), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_SL g321 ( .A(n_146), .B(n_261), .Y(n_321) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_147), .Y(n_173) );
INVx2_ASAP7_75t_L g238 ( .A(n_147), .Y(n_238) );
OR2x2_ASAP7_75t_L g300 ( .A(n_147), .B(n_301), .Y(n_300) );
O2A1O1Ixp5_ASAP7_75t_SL g149 ( .A1(n_150), .A2(n_151), .B(n_152), .C(n_153), .Y(n_149) );
INVx2_ASAP7_75t_L g165 ( .A(n_153), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_153), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_153), .A2(n_223), .B(n_224), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_153), .B(n_517), .Y(n_516) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_158), .Y(n_155) );
INVx1_ASAP7_75t_L g211 ( .A(n_158), .Y(n_211) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g450 ( .A(n_159), .Y(n_450) );
AND2x2_ASAP7_75t_L g239 ( .A(n_161), .B(n_175), .Y(n_239) );
AND2x2_ASAP7_75t_L g256 ( .A(n_161), .B(n_236), .Y(n_256) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g174 ( .A(n_162), .B(n_175), .Y(n_174) );
BUFx2_ASAP7_75t_L g259 ( .A(n_162), .Y(n_259) );
AND2x2_ASAP7_75t_L g388 ( .A(n_162), .B(n_389), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_165), .A2(n_199), .B(n_200), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_165), .A2(n_213), .B(n_214), .C(n_215), .Y(n_212) );
INVx2_ASAP7_75t_L g205 ( .A(n_167), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_167), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_168), .Y(n_170) );
NAND3xp33_ASAP7_75t_L g187 ( .A(n_169), .B(n_188), .C(n_191), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_169), .A2(n_222), .B(n_225), .Y(n_221) );
INVx4_ASAP7_75t_L g191 ( .A(n_170), .Y(n_191) );
OA21x2_ASAP7_75t_L g193 ( .A1(n_170), .A2(n_194), .B(n_203), .Y(n_193) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_170), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_170), .A2(n_523), .B(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g233 ( .A(n_171), .Y(n_233) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_174), .Y(n_171) );
AND2x2_ASAP7_75t_L g351 ( .A(n_172), .B(n_239), .Y(n_351) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g352 ( .A(n_173), .B(n_263), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_174), .A2(n_320), .B(n_322), .C(n_324), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_174), .B(n_320), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_174), .A2(n_250), .B1(n_393), .B2(n_394), .C(n_396), .Y(n_392) );
INVx1_ASAP7_75t_L g236 ( .A(n_175), .Y(n_236) );
INVx1_ASAP7_75t_L g272 ( .A(n_175), .Y(n_272) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_175), .Y(n_281) );
INVx2_ASAP7_75t_L g468 ( .A(n_178), .Y(n_468) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_178), .Y(n_481) );
INVx1_ASAP7_75t_L g453 ( .A(n_180), .Y(n_453) );
INVx1_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_192), .Y(n_182) );
AND2x2_ASAP7_75t_L g298 ( .A(n_183), .B(n_243), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_183), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_184), .B(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g390 ( .A(n_184), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g422 ( .A(n_184), .Y(n_422) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx3_ASAP7_75t_L g252 ( .A(n_185), .Y(n_252) );
AND2x2_ASAP7_75t_L g278 ( .A(n_185), .B(n_232), .Y(n_278) );
NOR2x1_ASAP7_75t_L g287 ( .A(n_185), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g294 ( .A(n_185), .B(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
INVx1_ASAP7_75t_L g230 ( .A(n_186), .Y(n_230) );
AO21x1_ASAP7_75t_L g229 ( .A1(n_188), .A2(n_191), .B(n_230), .Y(n_229) );
INVx3_ASAP7_75t_L g459 ( .A(n_191), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_191), .B(n_484), .Y(n_483) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_191), .A2(n_489), .B(n_496), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_191), .B(n_497), .Y(n_496) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_191), .A2(n_531), .B(n_538), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_192), .B(n_334), .Y(n_369) );
INVx1_ASAP7_75t_SL g373 ( .A(n_192), .Y(n_373) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_204), .Y(n_192) );
INVx3_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
AND2x2_ASAP7_75t_L g243 ( .A(n_193), .B(n_220), .Y(n_243) );
AND2x2_ASAP7_75t_L g265 ( .A(n_193), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g310 ( .A(n_193), .B(n_304), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_193), .B(n_242), .Y(n_391) );
INVx2_ASAP7_75t_L g213 ( .A(n_201), .Y(n_213) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g231 ( .A(n_204), .B(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g242 ( .A(n_204), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_204), .B(n_220), .Y(n_267) );
AND2x2_ASAP7_75t_L g303 ( .A(n_204), .B(n_304), .Y(n_303) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_216), .Y(n_204) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_205), .A2(n_221), .B(n_228), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .C(n_211), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_209), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_209), .A2(n_536), .B(n_537), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_211), .A2(n_492), .B(n_493), .C(n_494), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_213), .A2(n_449), .B(n_451), .Y(n_448) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_231), .Y(n_218) );
INVx1_ASAP7_75t_L g283 ( .A(n_219), .Y(n_283) );
AND2x2_ASAP7_75t_L g325 ( .A(n_219), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_219), .B(n_246), .Y(n_331) );
AOI21xp5_ASAP7_75t_SL g405 ( .A1(n_219), .A2(n_237), .B(n_260), .Y(n_405) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_229), .Y(n_219) );
OR2x2_ASAP7_75t_L g248 ( .A(n_220), .B(n_229), .Y(n_248) );
AND2x2_ASAP7_75t_L g295 ( .A(n_220), .B(n_232), .Y(n_295) );
INVx2_ASAP7_75t_L g304 ( .A(n_220), .Y(n_304) );
INVx1_ASAP7_75t_L g410 ( .A(n_220), .Y(n_410) );
AND2x2_ASAP7_75t_L g334 ( .A(n_229), .B(n_304), .Y(n_334) );
INVx1_ASAP7_75t_L g359 ( .A(n_229), .Y(n_359) );
AND2x2_ASAP7_75t_L g268 ( .A(n_231), .B(n_252), .Y(n_268) );
AND2x2_ASAP7_75t_L g280 ( .A(n_231), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_SL g398 ( .A(n_231), .Y(n_398) );
INVx2_ASAP7_75t_L g288 ( .A(n_232), .Y(n_288) );
AND2x2_ASAP7_75t_L g326 ( .A(n_232), .B(n_242), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_232), .B(n_410), .Y(n_409) );
OAI21xp33_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_239), .B(n_240), .Y(n_234) );
AND2x2_ASAP7_75t_L g341 ( .A(n_235), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g395 ( .A(n_235), .Y(n_395) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx1_ASAP7_75t_L g315 ( .A(n_236), .Y(n_315) );
BUFx2_ASAP7_75t_L g414 ( .A(n_236), .Y(n_414) );
BUFx2_ASAP7_75t_L g285 ( .A(n_237), .Y(n_285) );
AND2x2_ASAP7_75t_L g387 ( .A(n_237), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g370 ( .A(n_238), .Y(n_370) );
AND2x4_ASAP7_75t_L g297 ( .A(n_239), .B(n_260), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_239), .B(n_321), .Y(n_333) );
AOI32xp33_ASAP7_75t_L g257 ( .A1(n_240), .A2(n_258), .A3(n_260), .B1(n_262), .B2(n_263), .Y(n_257) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_243), .Y(n_240) );
INVx3_ASAP7_75t_L g246 ( .A(n_241), .Y(n_246) );
OR2x2_ASAP7_75t_L g382 ( .A(n_241), .B(n_338), .Y(n_382) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g251 ( .A(n_242), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g358 ( .A(n_242), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g250 ( .A(n_243), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g262 ( .A(n_243), .B(n_252), .Y(n_262) );
INVx1_ASAP7_75t_L g383 ( .A(n_243), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_243), .B(n_358), .Y(n_416) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_249), .B(n_253), .C(n_257), .Y(n_244) );
OAI322xp33_ASAP7_75t_L g353 ( .A1(n_245), .A2(n_290), .A3(n_354), .B1(n_356), .B2(n_360), .C1(n_361), .C2(n_365), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVxp67_ASAP7_75t_L g318 ( .A(n_246), .Y(n_318) );
INVx1_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g372 ( .A(n_248), .B(n_373), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_248), .B(n_288), .Y(n_419) );
INVxp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g311 ( .A(n_251), .Y(n_311) );
OR2x2_ASAP7_75t_L g397 ( .A(n_252), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_255), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g306 ( .A(n_256), .B(n_285), .Y(n_306) );
AND2x2_ASAP7_75t_L g377 ( .A(n_256), .B(n_290), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_256), .B(n_364), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_258), .A2(n_265), .B1(n_268), .B2(n_269), .C(n_274), .Y(n_264) );
OR2x2_ASAP7_75t_L g275 ( .A(n_258), .B(n_271), .Y(n_275) );
AND2x2_ASAP7_75t_L g363 ( .A(n_258), .B(n_364), .Y(n_363) );
AOI32xp33_ASAP7_75t_L g402 ( .A1(n_258), .A2(n_288), .A3(n_403), .B1(n_404), .B2(n_407), .Y(n_402) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_259), .B(n_295), .C(n_318), .Y(n_336) );
AND2x2_ASAP7_75t_L g362 ( .A(n_259), .B(n_355), .Y(n_362) );
INVxp67_ASAP7_75t_L g342 ( .A(n_260), .Y(n_342) );
BUFx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_263), .B(n_315), .Y(n_371) );
INVx2_ASAP7_75t_L g381 ( .A(n_263), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_263), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g350 ( .A(n_266), .Y(n_350) );
OR2x2_ASAP7_75t_L g276 ( .A(n_267), .B(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_269), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_273), .Y(n_269) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_272), .Y(n_355) );
AND2x2_ASAP7_75t_L g314 ( .A(n_273), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g360 ( .A(n_273), .Y(n_360) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_273), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AOI21xp33_ASAP7_75t_SL g299 ( .A1(n_275), .A2(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g393 ( .A(n_278), .B(n_303), .Y(n_393) );
AOI211xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_282), .B(n_292), .C(n_299), .Y(n_279) );
AND2x2_ASAP7_75t_L g323 ( .A(n_281), .B(n_291), .Y(n_323) );
INVx2_ASAP7_75t_L g338 ( .A(n_281), .Y(n_338) );
OR2x2_ASAP7_75t_L g376 ( .A(n_281), .B(n_339), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_281), .B(n_419), .Y(n_418) );
AOI211xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_284), .B(n_286), .C(n_289), .Y(n_282) );
INVxp67_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_285), .B(n_323), .Y(n_322) );
OAI211xp5_ASAP7_75t_L g404 ( .A1(n_286), .A2(n_381), .B(n_405), .C(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2x1p5_ASAP7_75t_L g302 ( .A(n_287), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g344 ( .A(n_288), .B(n_334), .Y(n_344) );
INVx1_ASAP7_75t_L g349 ( .A(n_288), .Y(n_349) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_293), .B(n_296), .Y(n_292) );
INVxp33_ASAP7_75t_L g400 ( .A(n_294), .Y(n_400) );
AND2x2_ASAP7_75t_L g379 ( .A(n_295), .B(n_358), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_300), .A2(n_362), .B(n_363), .Y(n_361) );
OAI322xp33_ASAP7_75t_L g380 ( .A1(n_302), .A2(n_381), .A3(n_382), .B1(n_383), .B2(n_384), .C1(n_386), .C2(n_390), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B1(n_312), .B2(n_316), .C(n_319), .Y(n_305) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g357 ( .A(n_310), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g401 ( .A(n_314), .Y(n_401) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_317), .B(n_337), .Y(n_403) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g366 ( .A(n_326), .B(n_334), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B1(n_332), .B2(n_334), .C(n_335), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_330), .A2(n_347), .B1(n_351), .B2(n_352), .C(n_353), .Y(n_346) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVxp67_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_334), .B(n_349), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B1(n_340), .B2(n_343), .Y(n_335) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx2_ASAP7_75t_SL g364 ( .A(n_339), .Y(n_364) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND5xp2_ASAP7_75t_L g345 ( .A(n_346), .B(n_367), .C(n_392), .D(n_402), .E(n_412), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_348), .B(n_350), .Y(n_347) );
NOR4xp25_ASAP7_75t_L g420 ( .A(n_349), .B(n_355), .C(n_421), .D(n_422), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_352), .A2(n_413), .B1(n_415), .B2(n_417), .C(n_420), .Y(n_412) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g411 ( .A(n_358), .Y(n_411) );
OAI322xp33_ASAP7_75t_L g368 ( .A1(n_362), .A2(n_369), .A3(n_370), .B1(n_371), .B2(n_372), .C1(n_374), .C2(n_378), .Y(n_368) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_380), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g413 ( .A(n_388), .B(n_414), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B1(n_400), .B2(n_401), .Y(n_396) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g740 ( .A(n_425), .Y(n_740) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g723 ( .A(n_427), .B(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g738 ( .A(n_427), .Y(n_738) );
AND2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_SL g431 ( .A(n_432), .B(n_676), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_611), .Y(n_432) );
NAND4xp25_ASAP7_75t_SL g433 ( .A(n_434), .B(n_556), .C(n_580), .D(n_603), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_498), .B1(n_528), .B2(n_540), .C(n_543), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_471), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_437), .A2(n_457), .B1(n_499), .B2(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_437), .B(n_472), .Y(n_614) );
AND2x2_ASAP7_75t_L g633 ( .A(n_437), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_437), .B(n_617), .Y(n_703) );
AND2x4_ASAP7_75t_L g437 ( .A(n_438), .B(n_457), .Y(n_437) );
AND2x2_ASAP7_75t_L g571 ( .A(n_438), .B(n_472), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_438), .B(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g594 ( .A(n_438), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g599 ( .A(n_438), .B(n_458), .Y(n_599) );
INVx2_ASAP7_75t_L g631 ( .A(n_438), .Y(n_631) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_438), .Y(n_675) );
AND2x2_ASAP7_75t_L g692 ( .A(n_438), .B(n_569), .Y(n_692) );
INVx5_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g610 ( .A(n_439), .B(n_569), .Y(n_610) );
AND2x4_ASAP7_75t_L g624 ( .A(n_439), .B(n_457), .Y(n_624) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_439), .Y(n_628) );
AND2x2_ASAP7_75t_L g648 ( .A(n_439), .B(n_563), .Y(n_648) );
AND2x2_ASAP7_75t_L g698 ( .A(n_439), .B(n_473), .Y(n_698) );
AND2x2_ASAP7_75t_L g708 ( .A(n_439), .B(n_458), .Y(n_708) );
OR2x6_ASAP7_75t_L g439 ( .A(n_440), .B(n_454), .Y(n_439) );
AOI21xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_445), .B(n_453), .Y(n_440) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx5_ASAP7_75t_L g463 ( .A(n_446), .Y(n_463) );
INVx2_ASAP7_75t_L g452 ( .A(n_450), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_452), .A2(n_479), .B(n_480), .C(n_481), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g504 ( .A1(n_452), .A2(n_481), .B(n_505), .C(n_506), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
AND2x2_ASAP7_75t_L g564 ( .A(n_457), .B(n_472), .Y(n_564) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_457), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_457), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g654 ( .A(n_457), .Y(n_654) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g542 ( .A(n_458), .B(n_487), .Y(n_542) );
AND2x2_ASAP7_75t_L g569 ( .A(n_458), .B(n_488), .Y(n_569) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B(n_470), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_463), .B(n_464), .C(n_469), .Y(n_461) );
INVx2_ASAP7_75t_L g477 ( .A(n_463), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_463), .A2(n_469), .B(n_514), .C(n_515), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g482 ( .A(n_469), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_471), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_485), .Y(n_471) );
OR2x2_ASAP7_75t_L g595 ( .A(n_472), .B(n_486), .Y(n_595) );
AND2x2_ASAP7_75t_L g632 ( .A(n_472), .B(n_542), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_472), .B(n_563), .Y(n_643) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_472), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_472), .B(n_599), .Y(n_716) );
INVx5_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g541 ( .A(n_473), .Y(n_541) );
AND2x2_ASAP7_75t_L g550 ( .A(n_473), .B(n_486), .Y(n_550) );
AND2x2_ASAP7_75t_L g666 ( .A(n_473), .B(n_561), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_473), .B(n_599), .Y(n_688) );
OR2x6_ASAP7_75t_L g473 ( .A(n_474), .B(n_483), .Y(n_473) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_486), .Y(n_634) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_487), .Y(n_586) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g563 ( .A(n_488), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_495), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_508), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_499), .B(n_576), .Y(n_695) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_500), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g547 ( .A(n_500), .B(n_548), .Y(n_547) );
INVx5_ASAP7_75t_SL g555 ( .A(n_500), .Y(n_555) );
OR2x2_ASAP7_75t_L g578 ( .A(n_500), .B(n_548), .Y(n_578) );
OR2x2_ASAP7_75t_L g588 ( .A(n_500), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g651 ( .A(n_500), .B(n_510), .Y(n_651) );
AND2x2_ASAP7_75t_SL g689 ( .A(n_500), .B(n_509), .Y(n_689) );
NOR4xp25_ASAP7_75t_L g710 ( .A(n_500), .B(n_631), .C(n_711), .D(n_712), .Y(n_710) );
AND2x2_ASAP7_75t_L g720 ( .A(n_500), .B(n_552), .Y(n_720) );
OR2x6_ASAP7_75t_L g500 ( .A(n_501), .B(n_507), .Y(n_500) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g545 ( .A(n_509), .B(n_541), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_509), .B(n_547), .Y(n_714) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
OR2x2_ASAP7_75t_L g554 ( .A(n_510), .B(n_555), .Y(n_554) );
INVx3_ASAP7_75t_L g561 ( .A(n_510), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_510), .B(n_530), .Y(n_573) );
INVxp67_ASAP7_75t_L g576 ( .A(n_510), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_510), .B(n_548), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_510), .B(n_520), .Y(n_642) );
AND2x2_ASAP7_75t_L g657 ( .A(n_510), .B(n_552), .Y(n_657) );
OR2x2_ASAP7_75t_L g686 ( .A(n_510), .B(n_520), .Y(n_686) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_518), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_519), .B(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_519), .B(n_555), .Y(n_694) );
OR2x2_ASAP7_75t_L g715 ( .A(n_519), .B(n_592), .Y(n_715) );
INVx1_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g529 ( .A(n_520), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g552 ( .A(n_520), .B(n_548), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_520), .B(n_530), .Y(n_567) );
AND2x2_ASAP7_75t_L g637 ( .A(n_520), .B(n_561), .Y(n_637) );
AND2x2_ASAP7_75t_L g671 ( .A(n_520), .B(n_555), .Y(n_671) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_521), .B(n_555), .Y(n_574) );
AND2x2_ASAP7_75t_L g602 ( .A(n_521), .B(n_530), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_528), .B(n_610), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_529), .A2(n_617), .B1(n_653), .B2(n_670), .C(n_672), .Y(n_669) );
INVx5_ASAP7_75t_SL g548 ( .A(n_530), .Y(n_548) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_534), .Y(n_531) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
OAI33xp33_ASAP7_75t_L g568 ( .A1(n_541), .A2(n_569), .A3(n_570), .B1(n_572), .B2(n_575), .B3(n_579), .Y(n_568) );
OR2x2_ASAP7_75t_L g584 ( .A(n_541), .B(n_585), .Y(n_584) );
AOI322xp5_ASAP7_75t_L g693 ( .A1(n_541), .A2(n_610), .A3(n_617), .B1(n_694), .B2(n_695), .C1(n_696), .C2(n_699), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_541), .B(n_569), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_SL g717 ( .A1(n_541), .A2(n_569), .B(n_718), .C(n_720), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_542), .A2(n_557), .B1(n_562), .B2(n_565), .C(n_568), .Y(n_556) );
INVx1_ASAP7_75t_L g649 ( .A(n_542), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_542), .B(n_698), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_546), .B1(n_549), .B2(n_551), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g626 ( .A(n_547), .B(n_561), .Y(n_626) );
AND2x2_ASAP7_75t_L g684 ( .A(n_547), .B(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g592 ( .A(n_548), .B(n_555), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_548), .B(n_561), .Y(n_620) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_550), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_550), .B(n_628), .Y(n_682) );
OAI321xp33_ASAP7_75t_L g701 ( .A1(n_550), .A2(n_623), .A3(n_702), .B1(n_703), .B2(n_704), .C(n_705), .Y(n_701) );
INVx1_ASAP7_75t_L g668 ( .A(n_551), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_552), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g607 ( .A(n_552), .B(n_555), .Y(n_607) );
AOI321xp33_ASAP7_75t_L g665 ( .A1(n_552), .A2(n_569), .A3(n_666), .B1(n_667), .B2(n_668), .C(n_669), .Y(n_665) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g582 ( .A(n_554), .B(n_567), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_555), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_555), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_555), .B(n_641), .Y(n_678) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x4_ASAP7_75t_L g601 ( .A(n_559), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g566 ( .A(n_560), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g674 ( .A(n_561), .Y(n_674) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_564), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g597 ( .A(n_569), .Y(n_597) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_571), .B(n_606), .Y(n_655) );
OR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
OR2x2_ASAP7_75t_L g619 ( .A(n_574), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g664 ( .A(n_574), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_575), .A2(n_622), .B1(n_625), .B2(n_627), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g719 ( .A(n_578), .B(n_642), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_583), .B1(n_587), .B2(n_593), .C(n_596), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx2_ASAP7_75t_L g617 ( .A(n_586), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx1_ASAP7_75t_SL g663 ( .A(n_589), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_591), .B(n_641), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_591), .A2(n_659), .B(n_661), .Y(n_658) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g704 ( .A(n_592), .B(n_686), .Y(n_704) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_SL g606 ( .A(n_595), .Y(n_606) );
AOI21xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_600), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g650 ( .A(n_602), .B(n_651), .Y(n_650) );
INVxp67_ASAP7_75t_L g712 ( .A(n_602), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_607), .B(n_608), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_606), .B(n_624), .Y(n_660) );
INVxp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g681 ( .A(n_610), .Y(n_681) );
NAND5xp2_ASAP7_75t_L g611 ( .A(n_612), .B(n_629), .C(n_638), .D(n_658), .E(n_665), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B(n_618), .C(n_621), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g653 ( .A(n_617), .Y(n_653) );
CKINVDCx16_ASAP7_75t_R g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_625), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g667 ( .A(n_627), .Y(n_667) );
OAI21xp5_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_633), .B(n_635), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_630), .A2(n_684), .B1(n_687), .B2(n_689), .C(n_690), .Y(n_683) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
AOI321xp33_ASAP7_75t_L g638 ( .A1(n_631), .A2(n_639), .A3(n_643), .B1(n_644), .B2(n_650), .C(n_652), .Y(n_638) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g709 ( .A(n_643), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_645), .B(n_649), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g661 ( .A(n_646), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NOR2xp67_ASAP7_75t_SL g673 ( .A(n_647), .B(n_654), .Y(n_673) );
AOI321xp33_ASAP7_75t_SL g705 ( .A1(n_650), .A2(n_706), .A3(n_707), .B1(n_708), .B2(n_709), .C(n_710), .Y(n_705) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B(n_655), .C(n_656), .Y(n_652) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_663), .B(n_671), .Y(n_700) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .C(n_675), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_701), .C(n_713), .Y(n_676) );
OAI211xp5_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_679), .B(n_683), .C(n_693), .Y(n_677) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_681), .B(n_682), .Y(n_680) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_682), .A2(n_714), .B1(n_715), .B2(n_716), .C(n_717), .Y(n_713) );
INVx1_ASAP7_75t_L g702 ( .A(n_684), .Y(n_702) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g706 ( .A(n_704), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
CKINVDCx14_ASAP7_75t_R g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_724), .B(n_738), .Y(n_737) );
CKINVDCx14_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
NAND2xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .Y(n_742) );
NOR2xp33_ASAP7_75t_SL g743 ( .A(n_744), .B(n_746), .Y(n_743) );
INVx1_ASAP7_75t_SL g776 ( .A(n_744), .Y(n_776) );
INVx1_ASAP7_75t_L g775 ( .A(n_746), .Y(n_775) );
OA21x2_ASAP7_75t_L g778 ( .A1(n_746), .A2(n_766), .B(n_776), .Y(n_778) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
BUFx2_ASAP7_75t_L g766 ( .A(n_749), .Y(n_766) );
INVx2_ASAP7_75t_L g770 ( .A(n_749), .Y(n_770) );
INVxp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_765), .B(n_767), .Y(n_751) );
OAI22xp33_ASAP7_75t_SL g752 ( .A1(n_753), .A2(n_754), .B1(n_760), .B2(n_761), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
BUFx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
CKINVDCx6p67_ASAP7_75t_R g772 ( .A(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
endmodule