module real_aes_7477_n_207 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_174, n_156, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_183, n_205, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_3, n_41, n_140, n_153, n_75, n_178, n_19, n_71, n_180, n_40, n_49, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_81, n_133, n_48, n_204, n_37, n_117, n_97, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_207);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_97;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_207;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_216;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_455;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_498;
wire n_481;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_639;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_208;
wire n_215;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
AOI22xp5_ASAP7_75t_SL g399 ( .A1(n_0), .A2(n_179), .B1(n_371), .B2(n_400), .Y(n_399) );
AOI222xp33_ASAP7_75t_L g288 ( .A1(n_1), .A2(n_60), .B1(n_191), .B2(n_289), .C1(n_292), .C2(n_296), .Y(n_288) );
INVx1_ASAP7_75t_L g356 ( .A(n_2), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_3), .A2(n_85), .B1(n_284), .B2(n_408), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_4), .A2(n_15), .B1(n_463), .B2(n_464), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_5), .B(n_275), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_6), .A2(n_39), .B1(n_281), .B2(n_435), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g601 ( .A1(n_7), .A2(n_13), .B1(n_411), .B2(n_479), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_8), .A2(n_174), .B1(n_310), .B2(n_639), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_9), .A2(n_134), .B1(n_346), .B2(n_347), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_10), .A2(n_118), .B1(n_444), .B2(n_568), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_11), .A2(n_93), .B1(n_310), .B2(n_443), .Y(n_532) );
AOI222xp33_ASAP7_75t_L g507 ( .A1(n_12), .A2(n_95), .B1(n_165), .B2(n_408), .C1(n_508), .C2(n_509), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_14), .A2(n_112), .B1(n_505), .B2(n_575), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_16), .Y(n_405) );
AOI222xp33_ASAP7_75t_L g478 ( .A1(n_17), .A2(n_61), .B1(n_111), .B2(n_422), .C1(n_479), .C2(n_480), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_18), .B(n_575), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_19), .Y(n_390) );
AO22x2_ASAP7_75t_L g229 ( .A1(n_20), .A2(n_64), .B1(n_230), .B2(n_231), .Y(n_229) );
INVx1_ASAP7_75t_L g625 ( .A(n_20), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_21), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_22), .A2(n_151), .B1(n_497), .B2(n_498), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g370 ( .A1(n_23), .A2(n_205), .B1(n_244), .B2(n_371), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_24), .A2(n_160), .B1(n_292), .B2(n_411), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_25), .A2(n_206), .B1(n_369), .B2(n_568), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_26), .A2(n_190), .B1(n_361), .B2(n_563), .Y(n_562) );
AOI222xp33_ASAP7_75t_L g649 ( .A1(n_27), .A2(n_149), .B1(n_188), .B2(n_289), .C1(n_296), .C2(n_509), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_28), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_29), .A2(n_186), .B1(n_244), .B2(n_249), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_30), .B(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_31), .Y(n_436) );
INVx1_ASAP7_75t_L g556 ( .A(n_32), .Y(n_556) );
AO22x2_ASAP7_75t_L g233 ( .A1(n_33), .A2(n_67), .B1(n_230), .B2(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g626 ( .A(n_33), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_34), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_35), .A2(n_197), .B1(n_340), .B2(n_344), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_36), .A2(n_129), .B1(n_360), .B2(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_37), .A2(n_59), .B1(n_470), .B2(n_471), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_38), .A2(n_97), .B1(n_312), .B2(n_314), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_40), .A2(n_48), .B1(n_244), .B2(n_565), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_41), .Y(n_542) );
AOI22xp5_ASAP7_75t_SL g395 ( .A1(n_42), .A2(n_125), .B1(n_396), .B2(n_397), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_43), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_44), .A2(n_168), .B1(n_223), .B2(n_240), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_45), .A2(n_120), .B1(n_347), .B2(n_411), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_46), .A2(n_148), .B1(n_263), .B2(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_47), .Y(n_376) );
XNOR2x2_ASAP7_75t_L g219 ( .A(n_49), .B(n_220), .Y(n_219) );
AOI22xp5_ASAP7_75t_SL g393 ( .A1(n_50), .A2(n_110), .B1(n_361), .B2(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_51), .A2(n_167), .B1(n_341), .B2(n_344), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_52), .A2(n_629), .B1(n_630), .B2(n_650), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_52), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g334 ( .A1(n_53), .A2(n_130), .B1(n_335), .B2(n_337), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_54), .Y(n_424) );
AOI211xp5_ASAP7_75t_L g421 ( .A1(n_55), .A2(n_422), .B(n_423), .C(n_432), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_56), .A2(n_182), .B1(n_306), .B2(n_308), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_57), .A2(n_170), .B1(n_475), .B2(n_476), .Y(n_474) );
AOI22xp5_ASAP7_75t_SL g359 ( .A1(n_58), .A2(n_117), .B1(n_360), .B2(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g569 ( .A(n_62), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_63), .A2(n_119), .B1(n_369), .B2(n_498), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_65), .A2(n_108), .B1(n_337), .B2(n_479), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_66), .A2(n_200), .B1(n_396), .B2(n_642), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_68), .A2(n_156), .B1(n_245), .B2(n_315), .Y(n_609) );
INVx1_ASAP7_75t_L g215 ( .A(n_69), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_70), .A2(n_100), .B1(n_255), .B2(n_257), .Y(n_254) );
INVx1_ASAP7_75t_L g590 ( .A(n_71), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_72), .A2(n_194), .B1(n_534), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_73), .A2(n_106), .B1(n_443), .B2(n_444), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_74), .A2(n_155), .B1(n_319), .B2(n_568), .Y(n_606) );
AOI22xp5_ASAP7_75t_SL g366 ( .A1(n_75), .A2(n_181), .B1(n_367), .B2(n_369), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_76), .A2(n_143), .B1(n_296), .B2(n_347), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_77), .Y(n_317) );
INVx1_ASAP7_75t_L g211 ( .A(n_78), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_79), .A2(n_157), .B1(n_443), .B2(n_444), .Y(n_442) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_80), .A2(n_132), .B1(n_494), .B2(n_497), .Y(n_608) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_81), .A2(n_208), .B(n_216), .C(n_627), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_82), .A2(n_144), .B1(n_263), .B2(n_266), .Y(n_262) );
INVxp67_ASAP7_75t_L g659 ( .A(n_83), .Y(n_659) );
XOR2x2_ASAP7_75t_L g661 ( .A(n_83), .B(n_631), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_84), .B(n_340), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_86), .A2(n_185), .B1(n_500), .B2(n_501), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_87), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_88), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_89), .A2(n_166), .B1(n_292), .B2(n_411), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_90), .A2(n_135), .B1(n_241), .B2(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_91), .B(n_505), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_92), .A2(n_139), .B1(n_498), .B2(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_94), .B(n_343), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_96), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_98), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g579 ( .A(n_99), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_101), .A2(n_177), .B1(n_315), .B2(n_494), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_102), .A2(n_183), .B1(n_279), .B2(n_347), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_103), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_104), .A2(n_142), .B1(n_285), .B2(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_105), .A2(n_162), .B1(n_346), .B2(n_430), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_107), .A2(n_201), .B1(n_314), .B2(n_534), .Y(n_533) );
AOI22xp5_ASAP7_75t_SL g514 ( .A1(n_109), .A2(n_515), .B1(n_544), .B2(n_545), .Y(n_514) );
INVx1_ASAP7_75t_L g545 ( .A(n_109), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g320 ( .A(n_113), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_114), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_115), .B(n_275), .Y(n_428) );
AND2x2_ASAP7_75t_L g214 ( .A(n_116), .B(n_215), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_121), .A2(n_176), .B1(n_285), .B2(n_346), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_122), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_123), .A2(n_159), .B1(n_279), .B2(n_284), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_124), .Y(n_518) );
AND2x6_ASAP7_75t_L g210 ( .A(n_126), .B(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_126), .Y(n_619) );
AO22x2_ASAP7_75t_L g237 ( .A1(n_127), .A2(n_175), .B1(n_230), .B2(n_234), .Y(n_237) );
CKINVDCx16_ASAP7_75t_R g419 ( .A(n_128), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_131), .A2(n_189), .B1(n_319), .B2(n_363), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_133), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_136), .Y(n_503) );
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_137), .A2(n_192), .B1(n_319), .B2(n_360), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_138), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_140), .A2(n_154), .B1(n_322), .B2(n_494), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_141), .Y(n_610) );
AO22x2_ASAP7_75t_L g239 ( .A1(n_145), .A2(n_187), .B1(n_230), .B2(n_231), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_146), .A2(n_199), .B1(n_408), .B2(n_581), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_147), .Y(n_540) );
INVx1_ASAP7_75t_L g456 ( .A(n_150), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_152), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_153), .A2(n_163), .B1(n_314), .B2(n_467), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_158), .A2(n_203), .B1(n_559), .B2(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_161), .B(n_505), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_164), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_169), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_171), .Y(n_450) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_172), .A2(n_180), .B1(n_500), .B2(n_565), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_173), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_175), .B(n_624), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_178), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_184), .A2(n_301), .B1(n_302), .B2(n_348), .Y(n_300) );
INVx1_ASAP7_75t_L g348 ( .A(n_184), .Y(n_348) );
INVx1_ASAP7_75t_L g622 ( .A(n_187), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_193), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_195), .A2(n_198), .B1(n_634), .B2(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g230 ( .A(n_196), .Y(n_230) );
INVx1_ASAP7_75t_L g232 ( .A(n_196), .Y(n_232) );
OA22x2_ASAP7_75t_L g458 ( .A1(n_202), .A2(n_459), .B1(n_460), .B2(n_481), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_202), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_204), .Y(n_598) );
INVx1_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_212), .Y(n_209) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_211), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g657 ( .A1(n_212), .A2(n_617), .B(n_658), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_213), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI221xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_487), .B1(n_612), .B2(n_613), .C(n_614), .Y(n_216) );
INVx1_ASAP7_75t_L g612 ( .A(n_217), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_351), .B1(n_485), .B2(n_486), .Y(n_217) );
INVx1_ASAP7_75t_L g485 ( .A(n_218), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_299), .B1(n_349), .B2(n_350), .Y(n_218) );
INVx1_ASAP7_75t_L g350 ( .A(n_219), .Y(n_350) );
NAND4xp75_ASAP7_75t_L g220 ( .A(n_221), .B(n_253), .C(n_269), .D(n_288), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_243), .Y(n_221) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx5_ASAP7_75t_SL g319 ( .A(n_224), .Y(n_319) );
INVx4_ASAP7_75t_L g539 ( .A(n_224), .Y(n_539) );
INVx2_ASAP7_75t_SL g585 ( .A(n_224), .Y(n_585) );
INVx11_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx11_ASAP7_75t_L g368 ( .A(n_225), .Y(n_368) );
AND2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_235), .Y(n_225) );
AND2x4_ASAP7_75t_L g277 ( .A(n_226), .B(n_248), .Y(n_277) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g383 ( .A(n_227), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_233), .Y(n_227) );
AND2x2_ASAP7_75t_L g242 ( .A(n_228), .B(n_233), .Y(n_242) );
AND2x2_ASAP7_75t_L g246 ( .A(n_228), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g283 ( .A(n_229), .B(n_237), .Y(n_283) );
AND2x2_ASAP7_75t_L g287 ( .A(n_229), .B(n_233), .Y(n_287) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g234 ( .A(n_232), .Y(n_234) );
INVx2_ASAP7_75t_L g247 ( .A(n_233), .Y(n_247) );
INVx1_ASAP7_75t_L g268 ( .A(n_233), .Y(n_268) );
AND2x4_ASAP7_75t_L g241 ( .A(n_235), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g256 ( .A(n_235), .B(n_246), .Y(n_256) );
AND2x6_ASAP7_75t_L g291 ( .A(n_235), .B(n_287), .Y(n_291) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
AND2x2_ASAP7_75t_L g248 ( .A(n_236), .B(n_239), .Y(n_248) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_237), .B(n_239), .Y(n_252) );
AND2x2_ASAP7_75t_L g260 ( .A(n_237), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g261 ( .A(n_239), .Y(n_261) );
INVx1_ASAP7_75t_L g295 ( .A(n_239), .Y(n_295) );
INVx3_ASAP7_75t_L g643 ( .A(n_240), .Y(n_643) );
BUFx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
BUFx3_ASAP7_75t_L g322 ( .A(n_241), .Y(n_322) );
BUFx3_ASAP7_75t_L g397 ( .A(n_241), .Y(n_397) );
INVx6_ASAP7_75t_L g451 ( .A(n_241), .Y(n_451) );
AND2x2_ASAP7_75t_L g265 ( .A(n_242), .B(n_260), .Y(n_265) );
NAND2x1p5_ASAP7_75t_L g273 ( .A(n_242), .B(n_248), .Y(n_273) );
AND2x6_ASAP7_75t_L g341 ( .A(n_242), .B(n_248), .Y(n_341) );
INVx4_ASAP7_75t_L g307 ( .A(n_244), .Y(n_307) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
BUFx3_ASAP7_75t_L g402 ( .A(n_245), .Y(n_402) );
BUFx3_ASAP7_75t_L g500 ( .A(n_245), .Y(n_500) );
BUFx3_ASAP7_75t_L g639 ( .A(n_245), .Y(n_639) );
AND2x4_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
AND2x4_ASAP7_75t_L g250 ( .A(n_246), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g259 ( .A(n_246), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_246), .B(n_260), .Y(n_330) );
AND2x2_ASAP7_75t_L g294 ( .A(n_247), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g372 ( .A(n_247), .Y(n_372) );
INVx1_ASAP7_75t_L g384 ( .A(n_248), .Y(n_384) );
BUFx2_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
BUFx3_ASAP7_75t_L g310 ( .A(n_250), .Y(n_310) );
BUFx3_ASAP7_75t_L g369 ( .A(n_250), .Y(n_369) );
BUFx3_ASAP7_75t_L g400 ( .A(n_250), .Y(n_400) );
BUFx2_ASAP7_75t_L g444 ( .A(n_250), .Y(n_444) );
BUFx3_ASAP7_75t_L g501 ( .A(n_250), .Y(n_501) );
AND2x2_ASAP7_75t_L g371 ( .A(n_251), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x6_ASAP7_75t_L g267 ( .A(n_252), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_262), .Y(n_253) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_255), .Y(n_455) );
BUFx3_ASAP7_75t_L g470 ( .A(n_255), .Y(n_470) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
BUFx2_ASAP7_75t_SL g326 ( .A(n_256), .Y(n_326) );
INVx2_ASAP7_75t_L g364 ( .A(n_256), .Y(n_364) );
BUFx2_ASAP7_75t_SL g396 ( .A(n_256), .Y(n_396) );
BUFx4f_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
BUFx3_ASAP7_75t_L g360 ( .A(n_259), .Y(n_360) );
BUFx3_ASAP7_75t_L g498 ( .A(n_259), .Y(n_498) );
BUFx3_ASAP7_75t_L g637 ( .A(n_259), .Y(n_637) );
INVx1_ASAP7_75t_L g286 ( .A(n_261), .Y(n_286) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx4_ASAP7_75t_L g313 ( .A(n_264), .Y(n_313) );
INVx3_ASAP7_75t_L g361 ( .A(n_264), .Y(n_361) );
INVx5_ASAP7_75t_L g494 ( .A(n_264), .Y(n_494) );
INVx8_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx6_ASAP7_75t_SL g315 ( .A(n_267), .Y(n_315) );
INVx1_ASAP7_75t_SL g446 ( .A(n_267), .Y(n_446) );
INVx1_ASAP7_75t_SL g565 ( .A(n_267), .Y(n_565) );
INVx1_ASAP7_75t_L g282 ( .A(n_268), .Y(n_282) );
OA211x2_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_271), .B(n_274), .C(n_278), .Y(n_269) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g375 ( .A(n_272), .Y(n_375) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx3_ASAP7_75t_L g427 ( .A(n_273), .Y(n_427) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx5_ASAP7_75t_L g344 ( .A(n_276), .Y(n_344) );
INVx2_ASAP7_75t_L g505 ( .A(n_276), .Y(n_505) );
INVx4_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx2_ASAP7_75t_L g346 ( .A(n_281), .Y(n_346) );
BUFx3_ASAP7_75t_L g411 ( .A(n_281), .Y(n_411) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x4_ASAP7_75t_L g293 ( .A(n_283), .B(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g297 ( .A(n_283), .B(n_298), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g379 ( .A(n_283), .B(n_372), .Y(n_379) );
BUFx2_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_285), .Y(n_347) );
BUFx2_ASAP7_75t_SL g560 ( .A(n_285), .Y(n_560) );
BUFx3_ASAP7_75t_L g581 ( .A(n_285), .Y(n_581) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g528 ( .A(n_286), .Y(n_528) );
INVx1_ASAP7_75t_L g527 ( .A(n_287), .Y(n_527) );
INVx4_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI21xp5_ASAP7_75t_SL g332 ( .A1(n_290), .A2(n_333), .B(n_334), .Y(n_332) );
OAI22xp5_ASAP7_75t_SL g387 ( .A1(n_290), .A2(n_388), .B1(n_389), .B2(n_390), .Y(n_387) );
OAI21xp5_ASAP7_75t_SL g520 ( .A1(n_290), .A2(n_521), .B(n_522), .Y(n_520) );
INVx4_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g406 ( .A(n_291), .Y(n_406) );
BUFx3_ASAP7_75t_L g422 ( .A(n_291), .Y(n_422) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_291), .Y(n_508) );
INVx2_ASAP7_75t_L g557 ( .A(n_291), .Y(n_557) );
INVx4_ASAP7_75t_L g336 ( .A(n_292), .Y(n_336) );
INVx2_ASAP7_75t_L g389 ( .A(n_292), .Y(n_389) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_293), .Y(n_435) );
BUFx4f_ASAP7_75t_SL g479 ( .A(n_293), .Y(n_479) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_293), .Y(n_509) );
INVx1_ASAP7_75t_L g298 ( .A(n_295), .Y(n_298) );
BUFx4f_ASAP7_75t_L g337 ( .A(n_296), .Y(n_337) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx12f_ASAP7_75t_L g408 ( .A(n_297), .Y(n_408) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_297), .Y(n_559) );
INVx1_ASAP7_75t_L g349 ( .A(n_299), .Y(n_349) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_SL g302 ( .A(n_303), .B(n_331), .Y(n_302) );
NOR3xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_316), .C(n_323), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_311), .Y(n_304) );
INVx4_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx3_ASAP7_75t_L g443 ( .A(n_307), .Y(n_443) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx2_ASAP7_75t_L g467 ( .A(n_313), .Y(n_467) );
INVx2_ASAP7_75t_L g535 ( .A(n_313), .Y(n_535) );
BUFx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx2_ASAP7_75t_L g645 ( .A(n_315), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_320), .B2(n_321), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B1(n_327), .B2(n_328), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_325), .A2(n_328), .B1(n_542), .B2(n_543), .Y(n_541) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_328), .A2(n_453), .B1(n_454), .B2(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_332), .B(n_338), .Y(n_331) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND3xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_342), .C(n_345), .Y(n_338) );
BUFx4f_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx2_ASAP7_75t_L g476 ( .A(n_341), .Y(n_476) );
BUFx2_ASAP7_75t_L g575 ( .A(n_341), .Y(n_575) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_344), .Y(n_475) );
INVx1_ASAP7_75t_SL g431 ( .A(n_347), .Y(n_431) );
INVx1_ASAP7_75t_L g486 ( .A(n_351), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_415), .B1(n_483), .B2(n_484), .Y(n_351) );
INVx1_ASAP7_75t_L g483 ( .A(n_352), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_391), .B2(n_414), .Y(n_352) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
XNOR2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
NAND3x1_ASAP7_75t_SL g357 ( .A(n_358), .B(n_365), .C(n_373), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_362), .Y(n_358) );
INVx1_ASAP7_75t_L g465 ( .A(n_360), .Y(n_465) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g568 ( .A(n_364), .Y(n_568) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_370), .Y(n_365) );
INVx4_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g394 ( .A(n_368), .Y(n_394) );
INVx2_ASAP7_75t_SL g471 ( .A(n_368), .Y(n_471) );
INVx4_ASAP7_75t_L g634 ( .A(n_368), .Y(n_634) );
NOR3xp33_ASAP7_75t_L g373 ( .A(n_374), .B(n_381), .C(n_387), .Y(n_373) );
OAI22xp5_ASAP7_75t_SL g374 ( .A1(n_375), .A2(n_376), .B1(n_377), .B2(n_380), .Y(n_374) );
OAI22xp5_ASAP7_75t_SL g523 ( .A1(n_377), .A2(n_524), .B1(n_525), .B2(n_529), .Y(n_523) );
INVx3_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx4_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI21xp5_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_385), .B(n_386), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp5_ASAP7_75t_SL g517 ( .A1(n_383), .A2(n_427), .B1(n_518), .B2(n_519), .Y(n_517) );
INVx2_ASAP7_75t_L g414 ( .A(n_391), .Y(n_414) );
XOR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_413), .Y(n_391) );
NAND4xp75_ASAP7_75t_SL g392 ( .A(n_393), .B(n_395), .C(n_398), .D(n_403), .Y(n_392) );
INVx1_ASAP7_75t_L g449 ( .A(n_394), .Y(n_449) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_409), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B(n_407), .Y(n_404) );
INVx2_ASAP7_75t_L g439 ( .A(n_408), .Y(n_439) );
BUFx4f_ASAP7_75t_SL g480 ( .A(n_408), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
INVx1_ASAP7_75t_L g484 ( .A(n_415), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_457), .B1(n_458), .B2(n_482), .Y(n_415) );
INVx1_ASAP7_75t_SL g482 ( .A(n_416), .Y(n_482) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
XNOR2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_440), .Y(n_420) );
OAI211xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B(n_428), .C(n_429), .Y(n_423) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OA211x2_ASAP7_75t_L g502 ( .A1(n_427), .A2(n_503), .B(n_504), .C(n_506), .Y(n_502) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_436), .B2(n_437), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_447), .C(n_452), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_445), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B1(n_450), .B2(n_451), .Y(n_447) );
INVx2_ASAP7_75t_L g463 ( .A(n_451), .Y(n_463) );
INVx3_ASAP7_75t_L g497 ( .A(n_451), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_451), .A2(n_537), .B1(n_538), .B2(n_540), .Y(n_536) );
INVx2_ASAP7_75t_L g563 ( .A(n_451), .Y(n_563) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g481 ( .A(n_460), .Y(n_481) );
NAND4xp75_ASAP7_75t_L g460 ( .A(n_461), .B(n_468), .C(n_473), .D(n_478), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_466), .Y(n_461) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_472), .Y(n_468) );
AND2x2_ASAP7_75t_SL g473 ( .A(n_474), .B(n_477), .Y(n_473) );
INVx1_ASAP7_75t_L g613 ( .A(n_487), .Y(n_613) );
AOI22xp5_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_593), .B1(n_594), .B2(n_611), .Y(n_487) );
INVx1_ASAP7_75t_L g611 ( .A(n_488), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_511), .B1(n_591), .B2(n_592), .Y(n_488) );
INVx2_ASAP7_75t_SL g591 ( .A(n_489), .Y(n_591) );
XOR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_510), .Y(n_489) );
NAND4xp75_ASAP7_75t_L g490 ( .A(n_491), .B(n_495), .C(n_502), .D(n_507), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_499), .Y(n_495) );
INVx1_ASAP7_75t_L g592 ( .A(n_511), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B1(n_546), .B2(n_547), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g544 ( .A(n_515), .Y(n_544) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_530), .Y(n_515) );
NOR3xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_520), .C(n_523), .Y(n_516) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x6_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
NOR3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .C(n_541), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
XOR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_570), .Y(n_547) );
XOR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_569), .Y(n_548) );
NAND4xp75_ASAP7_75t_SL g549 ( .A(n_550), .B(n_561), .C(n_566), .D(n_567), .Y(n_549) );
NOR2xp67_ASAP7_75t_SL g550 ( .A(n_551), .B(n_555), .Y(n_550) );
NAND3xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .C(n_554), .Y(n_551) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B(n_558), .Y(n_555) );
OAI21xp5_ASAP7_75t_SL g578 ( .A1(n_557), .A2(n_579), .B(n_580), .Y(n_578) );
OAI21xp5_ASAP7_75t_L g597 ( .A1(n_557), .A2(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
XOR2x2_ASAP7_75t_SL g570 ( .A(n_571), .B(n_590), .Y(n_570) );
NAND2x1p5_ASAP7_75t_L g571 ( .A(n_572), .B(n_582), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_578), .Y(n_572) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .C(n_577), .Y(n_573) );
NOR2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_587), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx3_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
XOR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_610), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_596), .B(n_603), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_600), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
NOR2x1_ASAP7_75t_L g615 ( .A(n_616), .B(n_620), .Y(n_615) );
OR2x2_ASAP7_75t_SL g664 ( .A(n_616), .B(n_621), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_618), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_618), .B(n_655), .Y(n_658) );
CKINVDCx16_ASAP7_75t_R g655 ( .A(n_619), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
OAI322xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_651), .A3(n_652), .B1(n_656), .B2(n_659), .C1(n_660), .C2(n_662), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_630), .Y(n_629) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND4xp75_ASAP7_75t_L g631 ( .A(n_632), .B(n_640), .C(n_646), .D(n_649), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_638), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_644), .Y(n_640) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_SL g646 ( .A(n_647), .B(n_648), .Y(n_646) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
CKINVDCx16_ASAP7_75t_R g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_663), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_664), .Y(n_663) );
endmodule