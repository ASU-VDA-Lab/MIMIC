module fake_jpeg_27193_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_48),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_39),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_39),
.B1(n_31),
.B2(n_29),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_62),
.B1(n_37),
.B2(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_42),
.Y(n_68)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

CKINVDCx11_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_31),
.B(n_29),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_33),
.B1(n_30),
.B2(n_28),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_31),
.B1(n_29),
.B2(n_16),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_75),
.B1(n_76),
.B2(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_24),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_91),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_25),
.B1(n_27),
.B2(n_24),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_56),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_77),
.C(n_36),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_18),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_37),
.B1(n_16),
.B2(n_21),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_37),
.B1(n_16),
.B2(n_21),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_42),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_37),
.B1(n_40),
.B2(n_36),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_63),
.B1(n_51),
.B2(n_47),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_18),
.B1(n_33),
.B2(n_30),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_40),
.B1(n_36),
.B2(n_34),
.Y(n_86)
);

AO22x1_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_45),
.B1(n_51),
.B2(n_49),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_17),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_92),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_40),
.Y(n_90)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_103),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_93),
.B1(n_78),
.B2(n_92),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_124),
.Y(n_141)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_77),
.B1(n_73),
.B2(n_84),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_52),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_118),
.Y(n_126)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_63),
.B1(n_50),
.B2(n_45),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_122),
.B1(n_91),
.B2(n_57),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_52),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_121),
.B(n_86),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_71),
.A2(n_63),
.B1(n_57),
.B2(n_49),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_72),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_129),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_69),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_69),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_131),
.A2(n_136),
.B1(n_145),
.B2(n_109),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_142),
.B1(n_146),
.B2(n_152),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_103),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_112),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_77),
.B1(n_86),
.B2(n_79),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_137),
.B(n_99),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_150),
.Y(n_182)
);

BUFx12f_ASAP7_75t_SL g139 ( 
.A(n_120),
.Y(n_139)
);

OR2x2_ASAP7_75t_SL g178 ( 
.A(n_139),
.B(n_145),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_140),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_86),
.B1(n_85),
.B2(n_81),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_81),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_123),
.Y(n_183)
);

AO22x2_ASAP7_75t_SL g145 ( 
.A1(n_99),
.A2(n_82),
.B1(n_52),
.B2(n_85),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_118),
.A2(n_40),
.B1(n_36),
.B2(n_34),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_34),
.B(n_17),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_148),
.B(n_154),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_107),
.A2(n_0),
.B(n_1),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_94),
.Y(n_150)
);

AO22x1_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_155),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_32),
.B1(n_23),
.B2(n_17),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_32),
.B(n_23),
.Y(n_154)
);

AO22x1_ASAP7_75t_SL g155 ( 
.A1(n_114),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_106),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_187),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_158),
.B(n_160),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_109),
.C(n_104),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_166),
.C(n_189),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_113),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_161),
.B(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_164),
.A2(n_172),
.B1(n_13),
.B2(n_12),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_104),
.C(n_116),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_116),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_100),
.Y(n_170)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_175),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_125),
.A2(n_115),
.B1(n_110),
.B2(n_108),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_177),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_188),
.B(n_154),
.Y(n_204)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_181),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_141),
.B(n_100),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_147),
.Y(n_197)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_149),
.B1(n_102),
.B2(n_101),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_129),
.B(n_123),
.Y(n_187)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_145),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_127),
.B(n_101),
.C(n_102),
.Y(n_189)
);

AO22x1_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_145),
.B1(n_131),
.B2(n_136),
.Y(n_190)
);

AO22x1_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_178),
.B1(n_188),
.B2(n_176),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_169),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_199),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_185),
.A2(n_141),
.B1(n_155),
.B2(n_142),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_203),
.B1(n_210),
.B2(n_217),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_207),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_152),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_202),
.C(n_205),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_146),
.C(n_133),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_185),
.A2(n_155),
.B1(n_151),
.B2(n_148),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_158),
.B(n_156),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_151),
.C(n_149),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_151),
.C(n_155),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_15),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_211),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_173),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_14),
.C(n_13),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_176),
.B1(n_187),
.B2(n_182),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_157),
.B(n_12),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_215),
.B(n_180),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_173),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_206),
.Y(n_219)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_226),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_223),
.B(n_235),
.Y(n_243)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_175),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_224),
.B(n_217),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_163),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_238),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_212),
.A2(n_174),
.B1(n_177),
.B2(n_163),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_230),
.A2(n_232),
.B1(n_236),
.B2(n_237),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_169),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_233),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_196),
.A2(n_172),
.B1(n_174),
.B2(n_160),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_190),
.B(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_182),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_240),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_203),
.A2(n_180),
.B1(n_184),
.B2(n_186),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_207),
.A2(n_179),
.B1(n_5),
.B2(n_6),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_242),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_199),
.A2(n_179),
.B(n_5),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_192),
.C(n_209),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_244),
.B(n_245),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_192),
.C(n_198),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_224),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_254),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_202),
.C(n_201),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_257),
.C(n_233),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_201),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_215),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_259),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_208),
.C(n_218),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_225),
.C(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_261),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_211),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_249),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_210),
.C(n_190),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_270),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_268),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_233),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_232),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_269),
.B(n_272),
.Y(n_280)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_221),
.B1(n_219),
.B2(n_242),
.Y(n_271)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_246),
.A2(n_221),
.B1(n_226),
.B2(n_237),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_274),
.A2(n_266),
.B1(n_273),
.B2(n_276),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_250),
.C(n_254),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_277),
.C(n_266),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_241),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_243),
.A2(n_223),
.B1(n_11),
.B2(n_10),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_281),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_255),
.C(n_262),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_269),
.B1(n_274),
.B2(n_223),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_286),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_264),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_249),
.C(n_251),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_288),
.Y(n_300)
);

NAND3xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_11),
.C(n_10),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_277),
.A2(n_11),
.B(n_10),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_290),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_3),
.B(n_5),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_7),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_6),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_299),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_281),
.B(n_6),
.Y(n_295)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_295),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_303),
.C(n_291),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_283),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_283),
.A2(n_8),
.B1(n_9),
.B2(n_285),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_280),
.A2(n_8),
.B(n_9),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_304),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_289),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_311),
.C(n_279),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_SL g309 ( 
.A(n_300),
.B(n_289),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_310),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_287),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_293),
.B1(n_294),
.B2(n_297),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_292),
.C(n_302),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_315),
.A2(n_308),
.B(n_307),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_316),
.C(n_312),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_316),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_317),
.B(n_305),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_8),
.Y(n_322)
);


endmodule