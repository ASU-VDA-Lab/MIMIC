module fake_ariane_1514_n_837 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_837);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_837;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_677;
wire n_614;
wire n_604;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_804;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

BUFx3_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_79),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_52),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_132),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_63),
.Y(n_173)
);

BUFx2_ASAP7_75t_SL g174 ( 
.A(n_95),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_54),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_36),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_8),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_38),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_17),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_53),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_9),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_12),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_70),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_2),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_50),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_98),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_L g191 ( 
.A(n_33),
.B(n_31),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_78),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_24),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_58),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_127),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_57),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_82),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_16),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_46),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_65),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_156),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_138),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_14),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_34),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_112),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_74),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_106),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_137),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_28),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_80),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_83),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_93),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_88),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_47),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_102),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_149),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_20),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_30),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_115),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_89),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_69),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_96),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_62),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_141),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_73),
.B(n_6),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_61),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_113),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_9),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_23),
.Y(n_235)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

AND2x6_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_15),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_178),
.B(n_0),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_176),
.A2(n_207),
.B1(n_188),
.B2(n_200),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_179),
.A2(n_0),
.B(n_1),
.Y(n_247)
);

BUFx8_ASAP7_75t_SL g248 ( 
.A(n_206),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_177),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_186),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_181),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_189),
.B(n_1),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

OAI22x1_ASAP7_75t_R g260 ( 
.A1(n_234),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_205),
.Y(n_261)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_171),
.Y(n_262)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_192),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_193),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_201),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_231),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_199),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_210),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_214),
.Y(n_273)
);

OAI21x1_ASAP7_75t_L g274 ( 
.A1(n_222),
.A2(n_94),
.B(n_167),
.Y(n_274)
);

BUFx8_ASAP7_75t_SL g275 ( 
.A(n_170),
.Y(n_275)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_174),
.Y(n_276)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_185),
.Y(n_277)
);

OA21x2_ASAP7_75t_L g278 ( 
.A1(n_230),
.A2(n_5),
.B(n_6),
.Y(n_278)
);

OA21x2_ASAP7_75t_L g279 ( 
.A1(n_216),
.A2(n_7),
.B(n_8),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_199),
.B(n_7),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_185),
.B(n_10),
.Y(n_281)
);

BUFx12f_ASAP7_75t_L g282 ( 
.A(n_172),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_185),
.B(n_10),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_211),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_275),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_175),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_282),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_257),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_242),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_251),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_243),
.Y(n_292)
);

NOR2x1p5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_180),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_241),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_248),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_239),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_246),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_242),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_236),
.B(n_184),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_236),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_272),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_R g308 ( 
.A(n_236),
.B(n_194),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_256),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_256),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_238),
.B(n_11),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_196),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_280),
.B(n_235),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_265),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_259),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_268),
.B(n_197),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_R g320 ( 
.A(n_254),
.B(n_233),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_276),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_276),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_259),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_255),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_260),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_260),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_261),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_261),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_270),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_267),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_245),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_271),
.B(n_202),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_284),
.B(n_203),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_254),
.B(n_204),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_267),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_307),
.Y(n_336)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_283),
.C(n_258),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_312),
.B(n_266),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_266),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_320),
.B(n_240),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_315),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_290),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_286),
.B(n_332),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_261),
.Y(n_347)
);

INVx8_ASAP7_75t_L g348 ( 
.A(n_297),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_313),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_292),
.B(n_269),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_300),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_299),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_244),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_269),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_309),
.B(n_245),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_303),
.B(n_244),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_262),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_317),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_288),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_306),
.B(n_262),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_308),
.B(n_250),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_302),
.B(n_262),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_330),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_310),
.B(n_250),
.Y(n_365)
);

OR2x6_ASAP7_75t_L g366 ( 
.A(n_316),
.B(n_279),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_303),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_291),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_291),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_302),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_305),
.B(n_277),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_293),
.B(n_277),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_291),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_304),
.B(n_277),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_327),
.B(n_263),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_324),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_263),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_324),
.Y(n_380)
);

INVx8_ASAP7_75t_L g381 ( 
.A(n_287),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_323),
.B(n_263),
.Y(n_382)
);

AO22x1_ASAP7_75t_L g383 ( 
.A1(n_289),
.A2(n_237),
.B1(n_281),
.B2(n_226),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_304),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_319),
.B(n_249),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_311),
.B(n_249),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_331),
.B(n_213),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_319),
.B(n_237),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_329),
.A2(n_279),
.B1(n_278),
.B2(n_247),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_331),
.B(n_237),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_333),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_329),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_294),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_294),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_285),
.B(n_215),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_296),
.Y(n_396)
);

AOI221xp5_ASAP7_75t_L g397 ( 
.A1(n_325),
.A2(n_224),
.B1(n_218),
.B2(n_229),
.C(n_228),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_325),
.B(n_217),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_326),
.B(n_247),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_326),
.B(n_278),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_288),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_346),
.B(n_219),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_336),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_351),
.B(n_221),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_339),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_355),
.B(n_223),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_401),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_353),
.B(n_225),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_350),
.B(n_227),
.Y(n_410)
);

NAND3xp33_ASAP7_75t_SL g411 ( 
.A(n_397),
.B(n_13),
.C(n_14),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

BUFx12f_ASAP7_75t_L g413 ( 
.A(n_396),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_348),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_354),
.B(n_185),
.Y(n_415)
);

AND2x6_ASAP7_75t_SL g416 ( 
.A(n_395),
.B(n_191),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_347),
.B(n_185),
.Y(n_417)
);

BUFx4f_ASAP7_75t_L g418 ( 
.A(n_348),
.Y(n_418)
);

INVx5_ASAP7_75t_L g419 ( 
.A(n_366),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_357),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_341),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_337),
.B(n_274),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_337),
.B(n_18),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_348),
.Y(n_425)
);

AOI211xp5_ASAP7_75t_L g426 ( 
.A1(n_360),
.A2(n_168),
.B(n_21),
.C(n_22),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_343),
.B(n_19),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

INVx5_ASAP7_75t_L g429 ( 
.A(n_366),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_371),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_399),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_29),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_357),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_381),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_369),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_338),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_165),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_338),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_356),
.B(n_32),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_386),
.B(n_163),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_373),
.B(n_35),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_373),
.B(n_37),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_344),
.Y(n_443)
);

NOR2x1p5_ASAP7_75t_L g444 ( 
.A(n_396),
.B(n_39),
.Y(n_444)
);

NOR3x1_ASAP7_75t_L g445 ( 
.A(n_398),
.B(n_40),
.C(n_41),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_359),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_381),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_381),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_389),
.A2(n_42),
.B(n_43),
.Y(n_449)
);

INVx5_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_370),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_396),
.B(n_44),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_393),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_400),
.Y(n_454)
);

AO22x1_ASAP7_75t_L g455 ( 
.A1(n_391),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_L g456 ( 
.A(n_382),
.B(n_358),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_364),
.B(n_160),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_367),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_379),
.B(n_159),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_374),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_378),
.B(n_380),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_375),
.B(n_59),
.Y(n_462)
);

BUFx8_ASAP7_75t_L g463 ( 
.A(n_392),
.Y(n_463)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_361),
.B(n_158),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_383),
.A2(n_60),
.B1(n_64),
.B2(n_66),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_394),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_387),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_467)
);

NOR2x1p5_ASAP7_75t_L g468 ( 
.A(n_377),
.B(n_72),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_365),
.B(n_157),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_384),
.B(n_75),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_362),
.Y(n_471)
);

NOR2x1_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_363),
.Y(n_472)
);

BUFx12f_ASAP7_75t_L g473 ( 
.A(n_413),
.Y(n_473)
);

O2A1O1Ixp5_ASAP7_75t_L g474 ( 
.A1(n_410),
.A2(n_422),
.B(n_415),
.C(n_427),
.Y(n_474)
);

INVx3_ASAP7_75t_SL g475 ( 
.A(n_434),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_368),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_408),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_453),
.Y(n_478)
);

NAND3xp33_ASAP7_75t_SL g479 ( 
.A(n_406),
.B(n_372),
.C(n_385),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_418),
.B(n_372),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_436),
.B(n_438),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_466),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_405),
.B(n_352),
.Y(n_483)
);

NAND3xp33_ASAP7_75t_L g484 ( 
.A(n_402),
.B(n_376),
.C(n_349),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_407),
.A2(n_390),
.B(n_388),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_448),
.B(n_376),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_404),
.B(n_345),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_342),
.Y(n_488)
);

O2A1O1Ixp5_ASAP7_75t_L g489 ( 
.A1(n_440),
.A2(n_76),
.B(n_81),
.C(n_84),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_420),
.A2(n_85),
.B(n_86),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_419),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_403),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_411),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_439),
.B(n_92),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_449),
.B(n_419),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_443),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_439),
.B(n_97),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_414),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_419),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_433),
.B(n_99),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_446),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_461),
.A2(n_100),
.B(n_101),
.Y(n_502)
);

NAND3xp33_ASAP7_75t_L g503 ( 
.A(n_423),
.B(n_103),
.C(n_104),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_424),
.B(n_105),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_463),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_R g506 ( 
.A(n_425),
.B(n_107),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_430),
.B(n_108),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_456),
.B(n_109),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_412),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_421),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_452),
.B(n_110),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_429),
.B(n_111),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_429),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_R g514 ( 
.A(n_424),
.B(n_114),
.Y(n_514)
);

O2A1O1Ixp33_ASAP7_75t_L g515 ( 
.A1(n_409),
.A2(n_116),
.B(n_117),
.C(n_118),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_429),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_417),
.A2(n_123),
.B(n_125),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_450),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_424),
.Y(n_519)
);

BUFx12f_ASAP7_75t_L g520 ( 
.A(n_416),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_428),
.B(n_130),
.Y(n_521)
);

XOR2x2_ASAP7_75t_SL g522 ( 
.A(n_431),
.B(n_131),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_451),
.B(n_133),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_435),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_428),
.B(n_134),
.Y(n_525)
);

O2A1O1Ixp33_ASAP7_75t_L g526 ( 
.A1(n_441),
.A2(n_135),
.B(n_136),
.C(n_140),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_428),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_450),
.B(n_435),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_450),
.Y(n_529)
);

O2A1O1Ixp33_ASAP7_75t_L g530 ( 
.A1(n_442),
.A2(n_142),
.B(n_143),
.C(n_144),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_491),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_477),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_495),
.A2(n_437),
.B1(n_432),
.B2(n_460),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_492),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_491),
.Y(n_535)
);

OA21x2_ASAP7_75t_L g536 ( 
.A1(n_490),
.A2(n_470),
.B(n_462),
.Y(n_536)
);

AO21x2_ASAP7_75t_L g537 ( 
.A1(n_490),
.A2(n_459),
.B(n_457),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_496),
.Y(n_538)
);

BUFx12f_ASAP7_75t_L g539 ( 
.A(n_473),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_499),
.B(n_444),
.Y(n_540)
);

AO21x2_ASAP7_75t_L g541 ( 
.A1(n_484),
.A2(n_465),
.B(n_464),
.Y(n_541)
);

AO21x2_ASAP7_75t_L g542 ( 
.A1(n_485),
.A2(n_458),
.B(n_467),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_510),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_509),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_501),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_483),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_481),
.B(n_445),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_519),
.B(n_460),
.Y(n_548)
);

BUFx2_ASAP7_75t_SL g549 ( 
.A(n_491),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_529),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_476),
.Y(n_551)
);

BUFx4f_ASAP7_75t_L g552 ( 
.A(n_529),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_478),
.B(n_460),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_529),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_482),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_488),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_527),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_479),
.A2(n_469),
.B(n_468),
.Y(n_558)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_474),
.A2(n_455),
.B(n_426),
.Y(n_559)
);

OAI21x1_ASAP7_75t_L g560 ( 
.A1(n_500),
.A2(n_517),
.B(n_489),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_511),
.B(n_435),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_524),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_487),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_499),
.Y(n_564)
);

BUFx6f_ASAP7_75t_SL g565 ( 
.A(n_475),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_504),
.Y(n_566)
);

OR2x6_ASAP7_75t_L g567 ( 
.A(n_528),
.B(n_145),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_521),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_498),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_525),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_494),
.Y(n_571)
);

INVx6_ASAP7_75t_L g572 ( 
.A(n_520),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_503),
.Y(n_573)
);

OAI21x1_ASAP7_75t_SL g574 ( 
.A1(n_497),
.A2(n_146),
.B(n_147),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_505),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_513),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_513),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_514),
.Y(n_578)
);

AO21x2_ASAP7_75t_L g579 ( 
.A1(n_508),
.A2(n_150),
.B(n_153),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_539),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_532),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_534),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_560),
.A2(n_502),
.B(n_526),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_538),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_545),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_545),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_544),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_544),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_543),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_560),
.A2(n_530),
.B(n_515),
.Y(n_590)
);

NAND2x1p5_ASAP7_75t_L g591 ( 
.A(n_554),
.B(n_507),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_552),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_547),
.A2(n_495),
.B1(n_493),
.B2(n_512),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_543),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_546),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_550),
.Y(n_596)
);

OA21x2_ASAP7_75t_L g597 ( 
.A1(n_559),
.A2(n_523),
.B(n_518),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_547),
.A2(n_563),
.B1(n_556),
.B2(n_537),
.Y(n_598)
);

INVx3_ASAP7_75t_SL g599 ( 
.A(n_572),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_555),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_551),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_551),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_562),
.Y(n_603)
);

OAI21x1_ASAP7_75t_L g604 ( 
.A1(n_559),
.A2(n_516),
.B(n_472),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_562),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_552),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_550),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_546),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_533),
.A2(n_522),
.B1(n_486),
.B2(n_480),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_563),
.B(n_512),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_548),
.B(n_506),
.Y(n_611)
);

AOI21x1_ASAP7_75t_L g612 ( 
.A1(n_536),
.A2(n_154),
.B(n_155),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_548),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_573),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_573),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_536),
.A2(n_570),
.B(n_568),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_557),
.Y(n_617)
);

BUFx4f_ASAP7_75t_L g618 ( 
.A(n_550),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_539),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_569),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_572),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_566),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_550),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_550),
.Y(n_624)
);

AO21x2_ASAP7_75t_L g625 ( 
.A1(n_537),
.A2(n_542),
.B(n_541),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_R g626 ( 
.A(n_580),
.B(n_565),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_614),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_581),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_581),
.B(n_575),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_585),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_583),
.A2(n_574),
.B(n_536),
.Y(n_631)
);

NOR3xp33_ASAP7_75t_SL g632 ( 
.A(n_580),
.B(n_553),
.C(n_565),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_R g633 ( 
.A(n_619),
.B(n_565),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_586),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_582),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_613),
.B(n_569),
.Y(n_636)
);

BUFx5_ASAP7_75t_L g637 ( 
.A(n_595),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_584),
.Y(n_638)
);

CKINVDCx16_ASAP7_75t_R g639 ( 
.A(n_619),
.Y(n_639)
);

NOR2x1p5_ASAP7_75t_L g640 ( 
.A(n_611),
.B(n_531),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_599),
.Y(n_641)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_620),
.Y(n_642)
);

NAND2xp33_ASAP7_75t_R g643 ( 
.A(n_610),
.B(n_540),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_618),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_592),
.B(n_578),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_592),
.B(n_554),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_600),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_617),
.B(n_576),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_606),
.B(n_578),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_R g650 ( 
.A(n_610),
.B(n_540),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_621),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_593),
.A2(n_540),
.B(n_561),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_621),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_599),
.B(n_577),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_618),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_601),
.B(n_531),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_602),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_608),
.B(n_549),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_588),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_595),
.B(n_549),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_587),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_614),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_587),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_606),
.B(n_554),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_598),
.B(n_531),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_589),
.A2(n_537),
.B1(n_561),
.B2(n_558),
.Y(n_666)
);

XNOR2xp5_ASAP7_75t_L g667 ( 
.A(n_609),
.B(n_572),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_618),
.Y(n_668)
);

AOI222xp33_ASAP7_75t_L g669 ( 
.A1(n_615),
.A2(n_572),
.B1(n_566),
.B2(n_570),
.C1(n_568),
.C2(n_571),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_596),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_596),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_615),
.B(n_535),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_623),
.Y(n_673)
);

OR2x6_ASAP7_75t_L g674 ( 
.A(n_591),
.B(n_567),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_596),
.B(n_554),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_SL g676 ( 
.A1(n_597),
.A2(n_558),
.B1(n_541),
.B2(n_571),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_624),
.B(n_535),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_657),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_637),
.B(n_625),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_647),
.B(n_622),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_628),
.B(n_622),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_673),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_646),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_635),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_642),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_638),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_637),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_637),
.B(n_625),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_654),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_637),
.B(n_625),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_659),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_627),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_630),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_634),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_637),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_663),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_636),
.B(n_607),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_629),
.B(n_607),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_627),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_661),
.B(n_616),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_662),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_662),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_672),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_648),
.B(n_591),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_656),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_658),
.B(n_607),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_665),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_674),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_674),
.B(n_616),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_666),
.B(n_591),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_660),
.B(n_603),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_677),
.B(n_597),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_670),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_671),
.B(n_597),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_669),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_640),
.B(n_605),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_631),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_676),
.B(n_605),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_675),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_678),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_685),
.B(n_641),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_682),
.B(n_705),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_689),
.B(n_639),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_684),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_689),
.B(n_667),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_686),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_691),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_687),
.Y(n_728)
);

NAND3x1_ASAP7_75t_L g729 ( 
.A(n_698),
.B(n_633),
.C(n_626),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_712),
.B(n_675),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_692),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_L g732 ( 
.A(n_713),
.B(n_632),
.C(n_652),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_682),
.B(n_653),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_696),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_709),
.B(n_646),
.Y(n_735)
);

NAND3xp33_ASAP7_75t_L g736 ( 
.A(n_680),
.B(n_649),
.C(n_645),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_712),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_705),
.B(n_651),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_681),
.B(n_645),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_687),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_709),
.B(n_664),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_692),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_699),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_697),
.B(n_655),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_695),
.A2(n_558),
.B(n_542),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_719),
.B(n_649),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_699),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_719),
.B(n_644),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_693),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_737),
.B(n_679),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_734),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_731),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_722),
.B(n_703),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_720),
.Y(n_754)
);

NAND2x1_ASAP7_75t_L g755 ( 
.A(n_728),
.B(n_695),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_723),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_730),
.B(n_737),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_730),
.B(n_679),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_724),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_735),
.B(n_707),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_726),
.B(n_707),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_731),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_728),
.B(n_688),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_727),
.Y(n_764)
);

BUFx2_ASAP7_75t_SL g765 ( 
.A(n_729),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_721),
.B(n_703),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_735),
.B(n_709),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_744),
.B(n_690),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_765),
.A2(n_732),
.B1(n_729),
.B2(n_736),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_767),
.A2(n_745),
.B(n_725),
.C(n_715),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_757),
.B(n_741),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_751),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_766),
.B(n_738),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_754),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_768),
.B(n_739),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_752),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_750),
.B(n_728),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_750),
.B(n_740),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_759),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_760),
.A2(n_650),
.B1(n_643),
.B2(n_688),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_761),
.B(n_758),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_758),
.B(n_735),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_779),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_L g784 ( 
.A1(n_769),
.A2(n_704),
.B1(n_756),
.B2(n_733),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_770),
.A2(n_780),
.B1(n_773),
.B2(n_767),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_779),
.A2(n_764),
.B(n_763),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_772),
.A2(n_763),
.B(n_755),
.Y(n_787)
);

OAI31xp33_ASAP7_75t_L g788 ( 
.A1(n_774),
.A2(n_753),
.A3(n_749),
.B(n_767),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_781),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_789),
.B(n_775),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_788),
.B(n_782),
.Y(n_791)
);

NAND3xp33_ASAP7_75t_SL g792 ( 
.A(n_785),
.B(n_756),
.C(n_778),
.Y(n_792)
);

AOI211xp5_ASAP7_75t_L g793 ( 
.A1(n_784),
.A2(n_777),
.B(n_706),
.C(n_771),
.Y(n_793)
);

XOR2x2_ASAP7_75t_L g794 ( 
.A(n_786),
.B(n_741),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_784),
.B(n_740),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_790),
.B(n_787),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_793),
.B(n_783),
.Y(n_797)
);

AOI211xp5_ASAP7_75t_L g798 ( 
.A1(n_792),
.A2(n_714),
.B(n_741),
.C(n_746),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_791),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_797),
.A2(n_795),
.B(n_794),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_799),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_796),
.A2(n_776),
.B(n_716),
.Y(n_802)
);

OAI221xp5_ASAP7_75t_SL g803 ( 
.A1(n_800),
.A2(n_798),
.B1(n_704),
.B2(n_567),
.C(n_714),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_801),
.A2(n_710),
.B(n_718),
.C(n_690),
.Y(n_804)
);

O2A1O1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_802),
.A2(n_574),
.B(n_567),
.C(n_579),
.Y(n_805)
);

AOI222xp33_ASAP7_75t_L g806 ( 
.A1(n_801),
.A2(n_718),
.B1(n_694),
.B2(n_752),
.C1(n_762),
.C2(n_701),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_803),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_805),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_806),
.Y(n_809)
);

OAI221xp5_ASAP7_75t_L g810 ( 
.A1(n_804),
.A2(n_710),
.B1(n_567),
.B2(n_762),
.C(n_552),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_806),
.A2(n_748),
.B1(n_708),
.B2(n_579),
.Y(n_811)
);

NAND3x1_ASAP7_75t_L g812 ( 
.A(n_808),
.B(n_740),
.C(n_644),
.Y(n_812)
);

NAND4xp75_ASAP7_75t_L g813 ( 
.A(n_807),
.B(n_554),
.C(n_700),
.D(n_702),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_809),
.B(n_668),
.Y(n_814)
);

AOI221xp5_ASAP7_75t_L g815 ( 
.A1(n_811),
.A2(n_579),
.B1(n_542),
.B2(n_571),
.C(n_541),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_810),
.A2(n_717),
.B(n_664),
.Y(n_816)
);

AOI221xp5_ASAP7_75t_L g817 ( 
.A1(n_808),
.A2(n_571),
.B1(n_717),
.B2(n_742),
.C(n_743),
.Y(n_817)
);

NAND4xp25_ASAP7_75t_L g818 ( 
.A(n_808),
.B(n_535),
.C(n_564),
.D(n_708),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_814),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_818),
.Y(n_820)
);

OAI22x1_ASAP7_75t_L g821 ( 
.A1(n_812),
.A2(n_708),
.B1(n_564),
.B2(n_612),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_813),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_816),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_819),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_820),
.A2(n_817),
.B1(n_815),
.B2(n_711),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_822),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_821),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_827),
.A2(n_823),
.B1(n_825),
.B2(n_826),
.Y(n_828)
);

AOI31xp33_ASAP7_75t_L g829 ( 
.A1(n_824),
.A2(n_711),
.A3(n_612),
.B(n_564),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_827),
.A2(n_571),
.B1(n_747),
.B2(n_743),
.Y(n_830)
);

NOR2x1_ASAP7_75t_L g831 ( 
.A(n_824),
.B(n_683),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_831),
.Y(n_832)
);

OA22x2_ASAP7_75t_L g833 ( 
.A1(n_832),
.A2(n_828),
.B1(n_829),
.B2(n_830),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_833),
.A2(n_604),
.B(n_590),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_834),
.A2(n_594),
.B1(n_604),
.B2(n_747),
.Y(n_835)
);

OR2x6_ASAP7_75t_L g836 ( 
.A(n_835),
.B(n_683),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_836),
.A2(n_590),
.B1(n_583),
.B2(n_742),
.Y(n_837)
);


endmodule