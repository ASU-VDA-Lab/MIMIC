module fake_jpeg_9275_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVxp67_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_5),
.B(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_40),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_23),
.B1(n_15),
.B2(n_21),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_13),
.B1(n_29),
.B2(n_35),
.Y(n_54)
);

XNOR2x1_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_18),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_47),
.C(n_13),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_27),
.B1(n_22),
.B2(n_20),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_50),
.B1(n_35),
.B2(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_33),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_24),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_36),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_22),
.B1(n_20),
.B2(n_17),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_58),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_36),
.B1(n_34),
.B2(n_30),
.Y(n_80)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_64),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_61),
.B(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_29),
.B1(n_1),
.B2(n_4),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_63),
.B(n_37),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_61),
.B1(n_56),
.B2(n_62),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_36),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_49),
.B1(n_39),
.B2(n_43),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_79),
.B1(n_82),
.B2(n_65),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_49),
.B1(n_43),
.B2(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_83),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_60),
.A2(n_34),
.B1(n_30),
.B2(n_36),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

AO21x1_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_92),
.B(n_94),
.Y(n_108)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_90),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_67),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_80),
.B1(n_73),
.B2(n_76),
.Y(n_103)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_93),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_59),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_97),
.C(n_73),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_78),
.B1(n_83),
.B2(n_79),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_78),
.B1(n_84),
.B2(n_70),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_97),
.C(n_85),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_34),
.B1(n_30),
.B2(n_36),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_10),
.B1(n_6),
.B2(n_8),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_0),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_112),
.C(n_115),
.Y(n_122)
);

OAI21x1_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_94),
.B(n_92),
.Y(n_110)
);

AOI321xp33_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_113),
.A3(n_98),
.B1(n_105),
.B2(n_106),
.C(n_99),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_88),
.C(n_86),
.Y(n_112)
);

OA21x2_ASAP7_75t_SL g113 ( 
.A1(n_108),
.A2(n_102),
.B(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_114),
.B(n_98),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_88),
.Y(n_115)
);

XOR2x1_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_88),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_107),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_121),
.B(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_120),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_6),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_123),
.B(n_122),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_109),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.C1(n_0),
.C2(n_16),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_125),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_122),
.C(n_11),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_128),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_16),
.C(n_28),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_SL g132 ( 
.A(n_129),
.B(n_130),
.C(n_28),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_28),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_28),
.B1(n_131),
.B2(n_57),
.Y(n_134)
);


endmodule