module fake_jpeg_3580_n_425 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_425);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_425;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_6),
.B(n_11),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_54),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_13),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_58),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_56),
.B(n_61),
.Y(n_117)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_57),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_13),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_60),
.Y(n_167)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g119 ( 
.A(n_62),
.Y(n_119)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_64),
.Y(n_172)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_67),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_66),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_26),
.B(n_14),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_68),
.B(n_72),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_23),
.B(n_14),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_75),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_14),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_23),
.B(n_13),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_77),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_32),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_32),
.B(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_81),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_80),
.A2(n_33),
.B1(n_27),
.B2(n_46),
.Y(n_143)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_83),
.B(n_90),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_39),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_86),
.B(n_92),
.Y(n_151)
);

BUFx4f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_48),
.B(n_3),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_91),
.B(n_98),
.Y(n_182)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_93),
.Y(n_179)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_48),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_95),
.B(n_96),
.Y(n_154)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_38),
.B(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_7),
.Y(n_114)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_17),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_19),
.B(n_4),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_109),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_19),
.B(n_5),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_19),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_46),
.B1(n_36),
.B2(n_24),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

BUFx4f_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_114),
.B(n_135),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_43),
.B1(n_34),
.B2(n_53),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_116),
.A2(n_121),
.B1(n_133),
.B2(n_142),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_110),
.A2(n_43),
.B1(n_34),
.B2(n_39),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_71),
.B(n_51),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_124),
.B(n_139),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_105),
.A2(n_43),
.B1(n_34),
.B2(n_45),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_67),
.B(n_51),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_75),
.B(n_40),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_101),
.A2(n_34),
.B1(n_40),
.B2(n_45),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_143),
.A2(n_148),
.B1(n_150),
.B2(n_171),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_66),
.A2(n_25),
.B1(n_49),
.B2(n_37),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g211 ( 
.A1(n_146),
.A2(n_147),
.B1(n_153),
.B2(n_159),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_66),
.A2(n_25),
.B1(n_49),
.B2(n_37),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_85),
.A2(n_28),
.B1(n_36),
.B2(n_33),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_72),
.B(n_28),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_157),
.B(n_158),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_24),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_85),
.A2(n_27),
.B1(n_50),
.B2(n_44),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_99),
.A2(n_50),
.B1(n_8),
.B2(n_9),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_163),
.B1(n_89),
.B2(n_93),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_69),
.A2(n_7),
.B1(n_9),
.B2(n_112),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_54),
.B(n_90),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_170),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_111),
.B(n_63),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_169),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_87),
.B(n_111),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_59),
.B(n_94),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_79),
.B(n_106),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_177),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_74),
.B(n_103),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_132),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_70),
.B(n_73),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g181 ( 
.A(n_103),
.B(n_99),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_155),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_84),
.B1(n_88),
.B2(n_104),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_184),
.A2(n_198),
.B1(n_207),
.B2(n_231),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_119),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_185),
.B(n_192),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_156),
.A2(n_62),
.B(n_102),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_186),
.B(n_203),
.C(n_228),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_187),
.A2(n_206),
.B1(n_200),
.B2(n_205),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_123),
.A2(n_100),
.B1(n_137),
.B2(n_134),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_119),
.A2(n_153),
.B(n_159),
.C(n_155),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_189),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_125),
.B(n_126),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_191),
.B(n_213),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_193),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_154),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_206),
.Y(n_245)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_195),
.Y(n_242)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_115),
.B1(n_167),
.B2(n_164),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_200),
.B(n_216),
.Y(n_261)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_202),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_126),
.B(n_125),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_205),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_115),
.A2(n_172),
.B1(n_163),
.B2(n_149),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_165),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_214),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_117),
.B(n_182),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_131),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_131),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_232),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_151),
.A2(n_113),
.B1(n_134),
.B2(n_129),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_218),
.Y(n_244)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_132),
.Y(n_219)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_219),
.Y(n_277)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_131),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_138),
.B(n_180),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_221),
.B(n_224),
.Y(n_247)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_136),
.B(n_140),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_240),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_146),
.A2(n_147),
.B(n_116),
.C(n_160),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_225),
.A2(n_227),
.B1(n_234),
.B2(n_200),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_226),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_121),
.A2(n_142),
.B1(n_133),
.B2(n_128),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_118),
.B(n_120),
.Y(n_228)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_145),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_145),
.A2(n_150),
.B1(n_171),
.B2(n_120),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_130),
.B(n_122),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_161),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_SL g267 ( 
.A(n_233),
.B(n_236),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_173),
.A2(n_161),
.B1(n_152),
.B2(n_141),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_152),
.B(n_141),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_238),
.Y(n_257)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_144),
.A2(n_168),
.B1(n_169),
.B2(n_148),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_237),
.A2(n_216),
.B1(n_183),
.B2(n_223),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_144),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_119),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_185),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_125),
.B(n_126),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_119),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_241),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_255),
.A2(n_272),
.B1(n_211),
.B2(n_199),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_264),
.A2(n_274),
.B1(n_189),
.B2(n_234),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_190),
.B(n_228),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_266),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_190),
.B(n_208),
.Y(n_266)
);

OAI32xp33_ASAP7_75t_L g269 ( 
.A1(n_191),
.A2(n_240),
.A3(n_208),
.B1(n_229),
.B2(n_204),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_211),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_212),
.B(n_213),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_279),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_237),
.A2(n_225),
.B1(n_224),
.B2(n_203),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_241),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_273),
.B(n_278),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_226),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_192),
.B(n_219),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_195),
.B(n_217),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_284),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_186),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_287),
.B(n_293),
.Y(n_325)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_288),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_211),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_301),
.C(n_276),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_243),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_296),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_292),
.B(n_309),
.Y(n_335)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_236),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_299),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_243),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_297),
.A2(n_300),
.B1(n_316),
.B2(n_251),
.Y(n_324)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_302),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_259),
.B(n_233),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_272),
.A2(n_199),
.B1(n_211),
.B2(n_231),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_199),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_244),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_193),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_304),
.Y(n_327)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_242),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_264),
.A2(n_199),
.B1(n_209),
.B2(n_196),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_305),
.A2(n_263),
.B1(n_273),
.B2(n_254),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_249),
.B(n_197),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_306),
.B(n_308),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_281),
.B(n_201),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_249),
.B(n_220),
.Y(n_309)
);

A2O1A1O1Ixp25_ASAP7_75t_L g310 ( 
.A1(n_281),
.A2(n_202),
.B(n_222),
.C(n_230),
.D(n_261),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_310),
.A2(n_262),
.B(n_278),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_247),
.B(n_269),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_313),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_312),
.Y(n_339)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_276),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_315),
.Y(n_330)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_283),
.A2(n_255),
.B1(n_261),
.B2(n_247),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_252),
.B(n_248),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_317),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_261),
.A2(n_283),
.B(n_246),
.C(n_245),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_263),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_275),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_332),
.C(n_298),
.Y(n_345)
);

MAJx2_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_275),
.C(n_246),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g344 ( 
.A(n_322),
.B(n_297),
.CI(n_289),
.CON(n_344),
.SN(n_344)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_324),
.A2(n_331),
.B1(n_343),
.B2(n_313),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_300),
.A2(n_251),
.B1(n_242),
.B2(n_254),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_326),
.A2(n_305),
.B1(n_303),
.B2(n_296),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_286),
.B(n_250),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_334),
.A2(n_337),
.B(n_338),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_318),
.A2(n_292),
.B(n_316),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_291),
.Y(n_340)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_340),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_288),
.A2(n_253),
.B(n_270),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_341),
.A2(n_307),
.B(n_310),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_301),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_287),
.A2(n_256),
.B1(n_268),
.B2(n_270),
.Y(n_343)
);

AOI321xp33_ASAP7_75t_L g376 ( 
.A1(n_344),
.A2(n_319),
.A3(n_322),
.B1(n_336),
.B2(n_332),
.C(n_295),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_351),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_330),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_347),
.B(n_348),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_330),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_333),
.Y(n_349)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_342),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_320),
.B(n_286),
.C(n_294),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_338),
.A2(n_293),
.B(n_290),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_352),
.A2(n_354),
.B(n_359),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_353),
.A2(n_355),
.B1(n_357),
.B2(n_361),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_335),
.A2(n_325),
.B(n_329),
.Y(n_354)
);

BUFx24_ASAP7_75t_SL g356 ( 
.A(n_323),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_356),
.B(n_323),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_324),
.A2(n_343),
.B1(n_337),
.B2(n_325),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_358),
.A2(n_319),
.B(n_339),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_325),
.A2(n_285),
.B(n_312),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_334),
.A2(n_285),
.B1(n_302),
.B2(n_306),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_362),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_299),
.Y(n_363)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_363),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_357),
.A2(n_329),
.B1(n_335),
.B2(n_326),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_368),
.A2(n_374),
.B1(n_353),
.B2(n_349),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_355),
.A2(n_328),
.B1(n_339),
.B2(n_321),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_369),
.A2(n_348),
.B1(n_347),
.B2(n_361),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_360),
.A2(n_336),
.B(n_341),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_379),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_359),
.C(n_351),
.Y(n_387)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_376),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_352),
.A2(n_321),
.B1(n_327),
.B2(n_322),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_377),
.B(n_340),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_363),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_375),
.B(n_350),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_382),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_379),
.A2(n_370),
.B1(n_372),
.B2(n_378),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_381),
.A2(n_388),
.B1(n_391),
.B2(n_374),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_345),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_383),
.B(n_390),
.C(n_367),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_378),
.B(n_346),
.Y(n_385)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_385),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_366),
.C(n_364),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_367),
.B(n_346),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_389),
.A2(n_354),
.B(n_366),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_358),
.C(n_360),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_394),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_383),
.C(n_387),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_386),
.C(n_384),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_381),
.A2(n_373),
.B1(n_368),
.B2(n_369),
.Y(n_394)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_395),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_396),
.A2(n_365),
.B(n_327),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_400),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_390),
.B(n_364),
.C(n_354),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_402),
.B(n_408),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_398),
.A2(n_391),
.B(n_365),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_403),
.B(n_406),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_392),
.A2(n_388),
.B(n_386),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_404),
.B(n_262),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_397),
.A2(n_344),
.B1(n_376),
.B2(n_331),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_393),
.Y(n_411)
);

NAND3xp33_ASAP7_75t_L g418 ( 
.A(n_411),
.B(n_413),
.C(n_304),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_407),
.A2(n_344),
.B1(n_315),
.B2(n_314),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_412),
.B(n_402),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_403),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g417 ( 
.A1(n_414),
.A2(n_260),
.B(n_282),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_415),
.B(n_417),
.Y(n_420)
);

O2A1O1Ixp33_ASAP7_75t_L g416 ( 
.A1(n_410),
.A2(n_408),
.B(n_401),
.C(n_253),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_416),
.B(n_409),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_413),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_419),
.B(n_421),
.Y(n_423)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_420),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_422),
.B(n_420),
.C(n_268),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_423),
.Y(n_425)
);


endmodule