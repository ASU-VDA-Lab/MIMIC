module fake_jpeg_29642_n_239 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_239);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_239;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_48),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_0),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_22),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_68),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_21),
.B(n_27),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_27),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_25),
.B1(n_29),
.B2(n_19),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_37),
.A2(n_33),
.B1(n_24),
.B2(n_26),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_25),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_76),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_84),
.Y(n_131)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_80),
.A2(n_85),
.B1(n_89),
.B2(n_102),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_96),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_46),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_43),
.B1(n_41),
.B2(n_44),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_43),
.B1(n_41),
.B2(n_29),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_41),
.B1(n_33),
.B2(n_26),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_100),
.B1(n_101),
.B2(n_51),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_50),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_21),
.B1(n_26),
.B2(n_24),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_65),
.A2(n_26),
.B1(n_24),
.B2(n_33),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_64),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_24),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_105),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_58),
.A2(n_32),
.B1(n_31),
.B2(n_3),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_49),
.A2(n_32),
.B1(n_31),
.B2(n_6),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_64),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_51),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_49),
.A2(n_32),
.B1(n_31),
.B2(n_6),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_62),
.B1(n_4),
.B2(n_7),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_128),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_59),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_113),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_122),
.B1(n_107),
.B2(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_59),
.Y(n_113)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_78),
.A2(n_55),
.A3(n_58),
.B1(n_62),
.B2(n_16),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_103),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_92),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_101),
.B1(n_94),
.B2(n_95),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_16),
.C(n_15),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_84),
.A2(n_4),
.B(n_8),
.C(n_9),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_8),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_131),
.B(n_84),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_88),
.C(n_96),
.Y(n_177)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_143),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_104),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_122),
.B1(n_124),
.B2(n_120),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_147),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_89),
.B1(n_80),
.B2(n_97),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_152),
.B1(n_154),
.B2(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_99),
.B1(n_98),
.B2(n_91),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_98),
.B1(n_106),
.B2(n_104),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_155),
.B(n_81),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_117),
.B(n_125),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_157),
.A2(n_175),
.B(n_9),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_162),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_129),
.B(n_108),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_163),
.B(n_166),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_172),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_139),
.B(n_121),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_113),
.B(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_171),
.B1(n_169),
.B2(n_168),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_140),
.B(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_135),
.B(n_131),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_173),
.A2(n_114),
.B1(n_130),
.B2(n_87),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_128),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_176),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_136),
.C(n_156),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_161),
.B1(n_145),
.B2(n_169),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_182),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_183),
.C(n_186),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_142),
.A3(n_153),
.B1(n_141),
.B2(n_147),
.C1(n_155),
.C2(n_82),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_167),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_153),
.B1(n_114),
.B2(n_130),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_166),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_187),
.B1(n_158),
.B2(n_176),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_79),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_9),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_193),
.C(n_157),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_168),
.B1(n_165),
.B2(n_167),
.Y(n_192)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_14),
.C(n_12),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_163),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_204),
.Y(n_208)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_198),
.B(n_203),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_199),
.A2(n_202),
.B1(n_192),
.B2(n_181),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_191),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_185),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_159),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_162),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_207),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_170),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_184),
.B1(n_201),
.B2(n_207),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_211),
.A2(n_216),
.B1(n_200),
.B2(n_206),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_217),
.Y(n_220)
);

FAx1_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_194),
.CI(n_185),
.CON(n_213),
.SN(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_215),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_204),
.C(n_188),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_197),
.C(n_12),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_189),
.B1(n_178),
.B2(n_182),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_193),
.B(n_12),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_209),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_218),
.B(n_222),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_224),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_11),
.C(n_13),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_220),
.C(n_213),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_13),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_208),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_225),
.B(n_229),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_219),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_223),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_227),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_232),
.C(n_233),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_228),
.C(n_210),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_235),
.B(n_213),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_210),
.C(n_234),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_208),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_217),
.Y(n_239)
);


endmodule