module fake_netlist_1_8161_n_653 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_653);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_653;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_73;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_195;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_522;
wire n_264;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g72 ( .A(n_13), .Y(n_72) );
CKINVDCx16_ASAP7_75t_R g73 ( .A(n_11), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_58), .Y(n_74) );
INVxp33_ASAP7_75t_L g75 ( .A(n_70), .Y(n_75) );
INVx2_ASAP7_75t_L g76 ( .A(n_71), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_30), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_17), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_37), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_66), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_67), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_32), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_56), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_68), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_29), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_47), .Y(n_86) );
OR2x2_ASAP7_75t_L g87 ( .A(n_57), .B(n_14), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_12), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_22), .Y(n_89) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_63), .Y(n_90) );
INVx1_ASAP7_75t_SL g91 ( .A(n_26), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_5), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_50), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_55), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_18), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_69), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_49), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_54), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_13), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_31), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_5), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_64), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_28), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_11), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_3), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_39), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_41), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_46), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_21), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_59), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_52), .Y(n_111) );
INVxp33_ASAP7_75t_SL g112 ( .A(n_23), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_27), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_18), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_36), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_21), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_0), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_9), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_42), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_19), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_74), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_120), .B(n_0), .Y(n_122) );
AND2x6_ASAP7_75t_L g123 ( .A(n_74), .B(n_34), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_76), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_76), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_94), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_119), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_73), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_94), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_120), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_77), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_79), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_100), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_116), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_93), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_100), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_79), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_105), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_80), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_108), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_80), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_81), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_112), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_81), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_108), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_82), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_82), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_84), .Y(n_150) );
NOR2xp33_ASAP7_75t_R g151 ( .A(n_83), .B(n_35), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g152 ( .A1(n_72), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_98), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_90), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_85), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_96), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_75), .B(n_1), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_96), .Y(n_159) );
AND2x6_ASAP7_75t_L g160 ( .A(n_97), .B(n_38), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_72), .B(n_2), .Y(n_161) );
NAND2xp33_ASAP7_75t_L g162 ( .A(n_87), .B(n_40), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_97), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_87), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_121), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_158), .Y(n_167) );
CKINVDCx16_ASAP7_75t_R g168 ( .A(n_164), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_131), .B(n_114), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
INVx1_ASAP7_75t_SL g171 ( .A(n_135), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_131), .B(n_118), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_158), .B(n_118), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_137), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_137), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_137), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_132), .B(n_117), .Y(n_178) );
INVxp67_ASAP7_75t_SL g179 ( .A(n_122), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_123), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_121), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_121), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_154), .B(n_102), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_136), .B(n_102), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_132), .B(n_117), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_121), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_121), .Y(n_188) );
AO22x2_ASAP7_75t_L g189 ( .A1(n_152), .A2(n_115), .B1(n_113), .B2(n_103), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_130), .Y(n_190) );
OR2x2_ASAP7_75t_L g191 ( .A(n_122), .B(n_92), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_130), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_123), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_130), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_130), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_158), .B(n_115), .Y(n_196) );
BUFx2_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_140), .B(n_101), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_144), .B(n_113), .Y(n_199) );
INVxp67_ASAP7_75t_L g200 ( .A(n_128), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_130), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_133), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_133), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_140), .B(n_101), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_123), .A2(n_99), .B1(n_88), .B2(n_109), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_124), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_123), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_124), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_124), .Y(n_209) );
BUFx4f_ASAP7_75t_L g210 ( .A(n_123), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_125), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_133), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_142), .B(n_99), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_123), .Y(n_215) );
AO22x2_ASAP7_75t_L g216 ( .A1(n_152), .A2(n_103), .B1(n_110), .B2(n_106), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_127), .B(n_110), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_125), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_133), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_123), .Y(n_220) );
NAND2x1p5_ASAP7_75t_L g221 ( .A(n_138), .B(n_107), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_138), .Y(n_222) );
INVx5_ASAP7_75t_L g223 ( .A(n_123), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_142), .B(n_95), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_143), .B(n_107), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_143), .B(n_95), .Y(n_226) );
NOR2xp33_ASAP7_75t_R g227 ( .A(n_168), .B(n_164), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_166), .Y(n_228) );
AOI211xp5_ASAP7_75t_L g229 ( .A1(n_184), .A2(n_162), .B(n_161), .C(n_78), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_179), .B(n_145), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_166), .Y(n_231) );
OR2x2_ASAP7_75t_SL g232 ( .A(n_191), .B(n_139), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_197), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_181), .Y(n_234) );
INVx4_ASAP7_75t_L g235 ( .A(n_166), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_222), .Y(n_236) );
NAND2xp33_ASAP7_75t_SL g237 ( .A(n_167), .B(n_151), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_222), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_221), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_196), .B(n_145), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_167), .B(n_148), .Y(n_241) );
AO22x1_ASAP7_75t_L g242 ( .A1(n_171), .A2(n_160), .B1(n_123), .B2(n_104), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_222), .Y(n_243) );
CKINVDCx6p67_ASAP7_75t_R g244 ( .A(n_197), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_178), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_178), .A2(n_148), .B1(n_157), .B2(n_160), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_178), .Y(n_247) );
NOR2xp33_ASAP7_75t_R g248 ( .A(n_210), .B(n_139), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_186), .Y(n_249) );
NOR3xp33_ASAP7_75t_SL g250 ( .A(n_185), .B(n_161), .C(n_88), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_200), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_186), .Y(n_252) );
NOR2xp33_ASAP7_75t_R g253 ( .A(n_210), .B(n_162), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_174), .B(n_157), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_173), .B(n_138), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_181), .B(n_138), .Y(n_256) );
INVx4_ASAP7_75t_L g257 ( .A(n_221), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_220), .Y(n_258) );
AND3x1_ASAP7_75t_SL g259 ( .A(n_189), .B(n_89), .C(n_109), .Y(n_259) );
OR2x6_ASAP7_75t_L g260 ( .A(n_189), .B(n_216), .Y(n_260) );
OAI22xp5_ASAP7_75t_SL g261 ( .A1(n_169), .A2(n_89), .B1(n_106), .B2(n_86), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_181), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_174), .B(n_138), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_181), .Y(n_264) );
NOR2xp67_ASAP7_75t_L g265 ( .A(n_191), .B(n_150), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_173), .B(n_150), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_173), .B(n_155), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_220), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_186), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_204), .B(n_150), .Y(n_270) );
INVx4_ASAP7_75t_L g271 ( .A(n_221), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_204), .Y(n_272) );
NAND2x1p5_ASAP7_75t_L g273 ( .A(n_204), .B(n_156), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_224), .B(n_150), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_206), .Y(n_275) );
NOR3xp33_ASAP7_75t_SL g276 ( .A(n_199), .B(n_160), .C(n_6), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_224), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_224), .B(n_150), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_198), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_198), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_214), .Y(n_281) );
NOR3xp33_ASAP7_75t_SL g282 ( .A(n_217), .B(n_160), .C(n_6), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_214), .B(n_155), .Y(n_283) );
CKINVDCx8_ASAP7_75t_R g284 ( .A(n_181), .Y(n_284) );
NOR3xp33_ASAP7_75t_SL g285 ( .A(n_225), .B(n_160), .C(n_7), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_226), .B(n_156), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_206), .Y(n_287) );
NOR3xp33_ASAP7_75t_SL g288 ( .A(n_189), .B(n_160), .C(n_7), .Y(n_288) );
INVx4_ASAP7_75t_L g289 ( .A(n_223), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_226), .Y(n_290) );
NAND2x1p5_ASAP7_75t_L g291 ( .A(n_210), .B(n_156), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_208), .B(n_156), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_208), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_293), .Y(n_294) );
NOR2xp67_ASAP7_75t_L g295 ( .A(n_257), .B(n_223), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_257), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_260), .A2(n_189), .B1(n_216), .B2(n_205), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_244), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_239), .Y(n_299) );
OR2x6_ASAP7_75t_SL g300 ( .A(n_233), .B(n_216), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_293), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_271), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_271), .B(n_223), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_239), .B(n_193), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_235), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_275), .Y(n_306) );
OR2x6_ASAP7_75t_L g307 ( .A(n_260), .B(n_216), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_265), .B(n_182), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_234), .Y(n_309) );
OAI22xp33_ASAP7_75t_L g310 ( .A1(n_260), .A2(n_193), .B1(n_215), .B2(n_207), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_256), .A2(n_223), .B(n_193), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_273), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_279), .B(n_223), .Y(n_313) );
NAND2x1_ASAP7_75t_L g314 ( .A(n_289), .B(n_160), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_240), .B(n_182), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_280), .B(n_209), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_273), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_292), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_287), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_234), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_231), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_255), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_256), .A2(n_223), .B(n_193), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_258), .B(n_193), .Y(n_324) );
OA21x2_ASAP7_75t_L g325 ( .A1(n_276), .A2(n_282), .B(n_288), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_236), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_286), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_245), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_281), .A2(n_267), .B1(n_255), .B2(n_261), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_290), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_230), .A2(n_207), .B(n_215), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_240), .B(n_183), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_281), .B(n_209), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_267), .B(n_212), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_259), .A2(n_219), .B1(n_183), .B2(n_187), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_284), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_234), .Y(n_337) );
BUFx10_ASAP7_75t_L g338 ( .A(n_247), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_266), .A2(n_207), .B(n_215), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_227), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_254), .B(n_212), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_249), .Y(n_342) );
AO21x1_ASAP7_75t_L g343 ( .A1(n_229), .A2(n_163), .B(n_147), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_243), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_234), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_270), .A2(n_207), .B(n_215), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_307), .A2(n_251), .B1(n_248), .B2(n_277), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_306), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_307), .A2(n_248), .B1(n_252), .B2(n_269), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_307), .A2(n_259), .B1(n_250), .B2(n_272), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_307), .A2(n_237), .B1(n_235), .B2(n_246), .Y(n_351) );
OR2x6_ASAP7_75t_L g352 ( .A(n_307), .B(n_291), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_341), .B(n_263), .Y(n_353) );
INVx8_ASAP7_75t_L g354 ( .A(n_302), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_316), .Y(n_355) );
INVx4_ASAP7_75t_L g356 ( .A(n_299), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_316), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_297), .A2(n_246), .B1(n_243), .B2(n_241), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_330), .A2(n_228), .B1(n_238), .B2(n_253), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_299), .B(n_250), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_331), .A2(n_274), .B(n_278), .Y(n_361) );
OAI22xp33_ASAP7_75t_L g362 ( .A1(n_300), .A2(n_283), .B1(n_232), .B2(n_291), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_294), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_333), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_302), .Y(n_365) );
INVx4_ASAP7_75t_L g366 ( .A(n_299), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_294), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_306), .Y(n_368) );
BUFx2_ASAP7_75t_R g369 ( .A(n_300), .Y(n_369) );
CKINVDCx11_ASAP7_75t_R g370 ( .A(n_298), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_320), .A2(n_155), .B(n_156), .Y(n_371) );
INVx4_ASAP7_75t_L g372 ( .A(n_302), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_301), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_333), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g375 ( .A1(n_330), .A2(n_207), .B1(n_215), .B2(n_288), .Y(n_375) );
OR2x6_ASAP7_75t_L g376 ( .A(n_317), .B(n_242), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_317), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_318), .B(n_187), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_301), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_348), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_356), .B(n_302), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_362), .B(n_329), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g383 ( .A1(n_350), .A2(n_340), .B1(n_335), .B2(n_327), .C(n_322), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g384 ( .A1(n_360), .A2(n_325), .B1(n_336), .B2(n_296), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_348), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_356), .B(n_302), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_363), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_363), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_360), .A2(n_335), .B1(n_343), .B2(n_325), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_367), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_353), .B(n_341), .Y(n_391) );
OAI221xp5_ASAP7_75t_L g392 ( .A1(n_347), .A2(n_327), .B1(n_322), .B2(n_282), .C(n_276), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_355), .A2(n_318), .B1(n_343), .B2(n_328), .C(n_342), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_377), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_360), .A2(n_325), .B1(n_336), .B2(n_296), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_353), .B(n_312), .Y(n_396) );
AOI21x1_ASAP7_75t_L g397 ( .A1(n_361), .A2(n_314), .B(n_325), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_354), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_357), .B(n_312), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_352), .A2(n_328), .B1(n_342), .B2(n_296), .Y(n_400) );
AO31x2_ASAP7_75t_L g401 ( .A1(n_368), .A2(n_163), .A3(n_159), .B(n_149), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_352), .A2(n_310), .B1(n_315), .B2(n_332), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_354), .Y(n_403) );
OAI211xp5_ASAP7_75t_L g404 ( .A1(n_359), .A2(n_253), .B(n_285), .C(n_149), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_352), .A2(n_296), .B1(n_336), .B2(n_319), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_356), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_352), .A2(n_314), .B1(n_305), .B2(n_308), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_354), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_387), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_403), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_380), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_403), .Y(n_412) );
OAI211xp5_ASAP7_75t_SL g413 ( .A1(n_394), .A2(n_370), .B(n_349), .C(n_111), .Y(n_413) );
OAI33xp33_ASAP7_75t_L g414 ( .A1(n_387), .A2(n_375), .A3(n_159), .B1(n_163), .B2(n_149), .B3(n_147), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_381), .B(n_366), .Y(n_415) );
NOR3xp33_ASAP7_75t_SL g416 ( .A(n_383), .B(n_369), .C(n_374), .Y(n_416) );
AO21x2_ASAP7_75t_L g417 ( .A1(n_389), .A2(n_285), .B(n_371), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_388), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_388), .Y(n_419) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_382), .A2(n_366), .B1(n_354), .B2(n_367), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_389), .A2(n_366), .B1(n_376), .B2(n_373), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_391), .A2(n_364), .B1(n_351), .B2(n_358), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_399), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_402), .A2(n_379), .B1(n_373), .B2(n_376), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_399), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_403), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_390), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_390), .Y(n_428) );
OAI22xp33_ASAP7_75t_L g429 ( .A1(n_396), .A2(n_376), .B1(n_379), .B2(n_378), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_391), .A2(n_376), .B1(n_370), .B2(n_160), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_380), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_398), .B(n_378), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_403), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_406), .B(n_368), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_385), .Y(n_435) );
NAND4xp25_ASAP7_75t_L g436 ( .A(n_384), .B(n_159), .C(n_147), .D(n_155), .Y(n_436) );
NOR2xp33_ASAP7_75t_SL g437 ( .A(n_398), .B(n_372), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_385), .Y(n_438) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_381), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_381), .B(n_372), .Y(n_440) );
OR2x6_ASAP7_75t_L g441 ( .A(n_381), .B(n_372), .Y(n_441) );
OAI31xp33_ASAP7_75t_L g442 ( .A1(n_392), .A2(n_334), .A3(n_155), .B(n_305), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_409), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_423), .B(n_393), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_411), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_410), .B(n_395), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_410), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_418), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_418), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_425), .B(n_386), .Y(n_450) );
OAI33xp33_ASAP7_75t_L g451 ( .A1(n_413), .A2(n_125), .A3(n_126), .B1(n_129), .B2(n_134), .B3(n_141), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_419), .Y(n_452) );
OAI31xp33_ASAP7_75t_L g453 ( .A1(n_429), .A2(n_404), .A3(n_405), .B(n_407), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_434), .B(n_401), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_433), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_411), .Y(n_456) );
OAI31xp33_ASAP7_75t_L g457 ( .A1(n_436), .A2(n_386), .A3(n_400), .B(n_408), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_438), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_437), .B(n_386), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_427), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_431), .B(n_386), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_432), .B(n_408), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_434), .B(n_401), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_431), .B(n_401), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_428), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_438), .B(n_401), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_435), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_439), .B(n_401), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_441), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_415), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_422), .A2(n_126), .B1(n_129), .B2(n_134), .C(n_141), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_439), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_439), .Y(n_473) );
NAND3xp33_ASAP7_75t_L g474 ( .A(n_420), .B(n_146), .C(n_129), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_439), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_439), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_415), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_440), .B(n_365), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_416), .B(n_126), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_441), .B(n_365), .Y(n_480) );
OAI221xp5_ASAP7_75t_SL g481 ( .A1(n_442), .A2(n_134), .B1(n_141), .B2(n_146), .C(n_91), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_433), .B(n_146), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_441), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_441), .B(n_424), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_412), .B(n_365), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_421), .B(n_218), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_412), .Y(n_487) );
OAI33xp33_ASAP7_75t_L g488 ( .A1(n_430), .A2(n_177), .A3(n_176), .B1(n_175), .B2(n_172), .B3(n_170), .Y(n_488) );
INVx1_ASAP7_75t_SL g489 ( .A(n_447), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_445), .Y(n_490) );
AND4x1_ASAP7_75t_L g491 ( .A(n_457), .B(n_414), .C(n_8), .D(n_9), .Y(n_491) );
NAND2xp33_ASAP7_75t_SL g492 ( .A(n_469), .B(n_426), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_460), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_454), .B(n_426), .Y(n_494) );
NOR3xp33_ASAP7_75t_L g495 ( .A(n_479), .B(n_426), .C(n_397), .Y(n_495) );
AOI22x1_ASAP7_75t_L g496 ( .A1(n_469), .A2(n_218), .B1(n_8), .B2(n_10), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_465), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_443), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_448), .B(n_417), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_463), .B(n_4), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_470), .Y(n_501) );
NOR3xp33_ASAP7_75t_L g502 ( .A(n_451), .B(n_397), .C(n_165), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_449), .B(n_452), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_445), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_483), .B(n_417), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_456), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_463), .B(n_4), .Y(n_507) );
NOR3xp33_ASAP7_75t_SL g508 ( .A(n_446), .B(n_304), .C(n_12), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_478), .B(n_10), .Y(n_509) );
NOR4xp25_ASAP7_75t_SL g510 ( .A(n_481), .B(n_417), .C(n_15), .D(n_16), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_478), .B(n_14), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_467), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_470), .B(n_15), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_444), .B(n_16), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_450), .B(n_17), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_461), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_483), .B(n_19), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_477), .B(n_20), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_461), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_458), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_464), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_468), .B(n_24), .Y(n_522) );
NOR4xp25_ASAP7_75t_SL g523 ( .A(n_459), .B(n_22), .C(n_175), .D(n_177), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_464), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_462), .B(n_25), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_458), .Y(n_526) );
OAI33xp33_ASAP7_75t_L g527 ( .A1(n_484), .A2(n_165), .A3(n_170), .B1(n_172), .B2(n_176), .B3(n_180), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_466), .B(n_319), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_477), .B(n_371), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_468), .Y(n_530) );
BUFx2_ASAP7_75t_L g531 ( .A(n_455), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_472), .B(n_33), .Y(n_532) );
OR2x6_ASAP7_75t_L g533 ( .A(n_484), .B(n_303), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_473), .B(n_43), .Y(n_534) );
BUFx2_ASAP7_75t_L g535 ( .A(n_487), .Y(n_535) );
AOI21xp33_ASAP7_75t_L g536 ( .A1(n_514), .A2(n_480), .B(n_482), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_493), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_497), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_512), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_498), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_489), .B(n_487), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_530), .B(n_475), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_521), .B(n_476), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_516), .B(n_475), .Y(n_544) );
OAI21xp33_ASAP7_75t_L g545 ( .A1(n_508), .A2(n_476), .B(n_485), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_527), .A2(n_453), .B(n_488), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_519), .B(n_486), .Y(n_547) );
NOR4xp25_ASAP7_75t_L g548 ( .A(n_500), .B(n_474), .C(n_486), .D(n_471), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_504), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_504), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_508), .A2(n_295), .B(n_180), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_524), .B(n_321), .Y(n_552) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_515), .A2(n_151), .B1(n_344), .B2(n_203), .C(n_201), .Y(n_553) );
NAND2x1_ASAP7_75t_L g554 ( .A(n_531), .B(n_303), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_501), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_496), .A2(n_295), .B(n_303), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_525), .A2(n_344), .B1(n_326), .B2(n_305), .Y(n_557) );
AOI21xp5_ASAP7_75t_SL g558 ( .A1(n_517), .A2(n_303), .B(n_313), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_533), .A2(n_326), .B1(n_313), .B2(n_338), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_535), .B(n_44), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_495), .B(n_346), .C(n_339), .Y(n_561) );
AOI33xp33_ASAP7_75t_L g562 ( .A1(n_509), .A2(n_195), .A3(n_188), .B1(n_219), .B2(n_213), .B3(n_211), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_501), .B(n_45), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_507), .A2(n_313), .B1(n_337), .B2(n_320), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_525), .A2(n_338), .B1(n_313), .B2(n_324), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_533), .A2(n_345), .B1(n_337), .B2(n_320), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g567 ( .A1(n_491), .A2(n_195), .B1(n_213), .B2(n_211), .C(n_203), .Y(n_567) );
OAI21xp33_ASAP7_75t_L g568 ( .A1(n_499), .A2(n_345), .B(n_337), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_506), .Y(n_569) );
XOR2x2_ASAP7_75t_L g570 ( .A(n_511), .B(n_48), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_533), .A2(n_345), .B1(n_202), .B2(n_201), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_503), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_494), .B(n_51), .Y(n_573) );
OAI221xp5_ASAP7_75t_SL g574 ( .A1(n_513), .A2(n_323), .B1(n_311), .B2(n_202), .C(n_190), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_528), .B(n_53), .Y(n_575) );
NOR2xp33_ASAP7_75t_SL g576 ( .A(n_527), .B(n_338), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_526), .Y(n_577) );
OAI21xp5_ASAP7_75t_L g578 ( .A1(n_518), .A2(n_190), .B(n_188), .Y(n_578) );
AOI311xp33_ASAP7_75t_L g579 ( .A1(n_495), .A2(n_192), .A3(n_194), .B(n_62), .C(n_65), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_537), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_555), .B(n_492), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_541), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_572), .B(n_505), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_544), .B(n_505), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_538), .B(n_490), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_569), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_549), .Y(n_587) );
CKINVDCx16_ASAP7_75t_R g588 ( .A(n_560), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_539), .Y(n_589) );
INVxp33_ASAP7_75t_L g590 ( .A(n_554), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_540), .Y(n_591) );
NOR2x1_ASAP7_75t_L g592 ( .A(n_558), .B(n_522), .Y(n_592) );
NOR4xp25_ASAP7_75t_SL g593 ( .A(n_545), .B(n_510), .C(n_523), .D(n_522), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g594 ( .A(n_536), .B(n_502), .C(n_534), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_550), .B(n_520), .Y(n_595) );
OAI21xp5_ASAP7_75t_SL g596 ( .A1(n_563), .A2(n_534), .B(n_529), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_543), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_543), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_577), .B(n_532), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_570), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_L g601 ( .A1(n_548), .A2(n_546), .B(n_567), .C(n_574), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_542), .B(n_60), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_547), .B(n_61), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_552), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_576), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_573), .B(n_309), .Y(n_606) );
OAI21xp5_ASAP7_75t_SL g607 ( .A1(n_557), .A2(n_309), .B(n_338), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_597), .B(n_568), .Y(n_608) );
OAI21xp33_ASAP7_75t_L g609 ( .A1(n_583), .A2(n_562), .B(n_575), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_598), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_586), .Y(n_611) );
XNOR2xp5_ASAP7_75t_L g612 ( .A(n_600), .B(n_564), .Y(n_612) );
XOR2x2_ASAP7_75t_L g613 ( .A(n_582), .B(n_571), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_580), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_589), .B(n_578), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_596), .A2(n_566), .B1(n_565), .B2(n_553), .Y(n_616) );
A2O1A1Ixp33_ASAP7_75t_SL g617 ( .A1(n_593), .A2(n_551), .B(n_556), .C(n_559), .Y(n_617) );
AOI211xp5_ASAP7_75t_L g618 ( .A1(n_590), .A2(n_566), .B(n_561), .C(n_579), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_604), .B(n_309), .Y(n_619) );
INVxp67_ASAP7_75t_L g620 ( .A(n_591), .Y(n_620) );
AOI222xp33_ASAP7_75t_L g621 ( .A1(n_594), .A2(n_262), .B1(n_264), .B2(n_268), .C1(n_309), .C2(n_581), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_585), .Y(n_622) );
OAI211xp5_ASAP7_75t_L g623 ( .A1(n_605), .A2(n_262), .B(n_264), .C(n_607), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_584), .B(n_262), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_614), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_611), .B(n_595), .Y(n_626) );
NOR2xp33_ASAP7_75t_R g627 ( .A(n_612), .B(n_588), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_613), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_622), .Y(n_629) );
AOI221x1_ASAP7_75t_SL g630 ( .A1(n_618), .A2(n_603), .B1(n_602), .B2(n_587), .C(n_599), .Y(n_630) );
OAI211xp5_ASAP7_75t_L g631 ( .A1(n_617), .A2(n_599), .B(n_606), .C(n_616), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_621), .B(n_623), .Y(n_632) );
BUFx2_ASAP7_75t_L g633 ( .A(n_620), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_624), .B(n_608), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_608), .B(n_609), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_619), .A2(n_588), .B1(n_592), .B2(n_590), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_611), .A2(n_588), .B1(n_590), .B2(n_592), .Y(n_637) );
OAI322xp33_ASAP7_75t_L g638 ( .A1(n_611), .A2(n_612), .A3(n_615), .B1(n_620), .B2(n_600), .C1(n_589), .C2(n_601), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_610), .Y(n_639) );
AND2x4_ASAP7_75t_L g640 ( .A(n_633), .B(n_634), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_630), .B(n_635), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_625), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_639), .Y(n_643) );
INVx4_ASAP7_75t_L g644 ( .A(n_628), .Y(n_644) );
NOR2xp67_ASAP7_75t_L g645 ( .A(n_644), .B(n_637), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_641), .A2(n_628), .B1(n_636), .B2(n_631), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_643), .Y(n_647) );
OAI222xp33_ASAP7_75t_L g648 ( .A1(n_646), .A2(n_641), .B1(n_644), .B2(n_636), .C1(n_632), .C2(n_640), .Y(n_648) );
NAND2xp33_ASAP7_75t_R g649 ( .A(n_645), .B(n_627), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_649), .Y(n_650) );
BUFx2_ASAP7_75t_L g651 ( .A(n_648), .Y(n_651) );
AOI322xp5_ASAP7_75t_L g652 ( .A1(n_651), .A2(n_647), .A3(n_640), .B1(n_629), .B2(n_638), .C1(n_642), .C2(n_626), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_652), .A2(n_651), .B(n_650), .Y(n_653) );
endmodule