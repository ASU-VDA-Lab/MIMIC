module fake_jpeg_27574_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_17),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_31),
.Y(n_49)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_20),
.B1(n_22),
.B2(n_32),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_43),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_63),
.B1(n_40),
.B2(n_24),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_32),
.B1(n_24),
.B2(n_22),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_59),
.C(n_66),
.Y(n_73)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_22),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_60),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_20),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_21),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_21),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_43),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_72),
.B(n_77),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_24),
.B1(n_16),
.B2(n_26),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_86),
.B1(n_89),
.B2(n_40),
.Y(n_102)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_80),
.B(n_82),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_59),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_50),
.A2(n_18),
.B1(n_19),
.B2(n_30),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_82),
.B1(n_80),
.B2(n_56),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_90),
.A2(n_97),
.B1(n_105),
.B2(n_64),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_111),
.Y(n_118)
);

AOI32xp33_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_58),
.A3(n_49),
.B1(n_36),
.B2(n_59),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_99),
.B(n_41),
.Y(n_129)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_100),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_46),
.B1(n_52),
.B2(n_48),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_49),
.B(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_59),
.B1(n_44),
.B2(n_48),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_110),
.B1(n_69),
.B2(n_79),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_57),
.B1(n_51),
.B2(n_19),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_74),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_104),
.Y(n_125)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_44),
.B1(n_60),
.B2(n_64),
.Y(n_105)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_28),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_78),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_75),
.B1(n_71),
.B2(n_44),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_75),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_27),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_25),
.C(n_30),
.Y(n_117)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_116),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_97),
.B1(n_109),
.B2(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_91),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_45),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_119),
.A2(n_129),
.B(n_134),
.Y(n_157)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_102),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_131),
.B1(n_99),
.B2(n_100),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_27),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_132),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_68),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_83),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_103),
.A2(n_18),
.B1(n_28),
.B2(n_26),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_90),
.B(n_25),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_136),
.B(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_23),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_154),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_140),
.A2(n_153),
.B(n_160),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_144),
.B1(n_147),
.B2(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_143),
.B(n_146),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_94),
.B1(n_107),
.B2(n_104),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_125),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_68),
.B1(n_57),
.B2(n_106),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_159),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_41),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_150),
.B(n_151),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_43),
.Y(n_151)
);

AOI32xp33_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_47),
.A3(n_29),
.B1(n_45),
.B2(n_83),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_123),
.B(n_23),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_119),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_121),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_134),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_158),
.A2(n_122),
.B1(n_118),
.B2(n_136),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_165),
.A2(n_168),
.B1(n_170),
.B2(n_173),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_171),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_115),
.B1(n_119),
.B2(n_114),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_151),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_187),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_132),
.B1(n_133),
.B2(n_124),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_135),
.B1(n_120),
.B2(n_137),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_183),
.B1(n_152),
.B2(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_117),
.B(n_0),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_155),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_184),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_143),
.C(n_160),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_161),
.C(n_163),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_47),
.B1(n_29),
.B2(n_45),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_141),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_47),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_148),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_203),
.Y(n_214)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_162),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_198),
.C(n_176),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_163),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_196),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_205),
.B1(n_206),
.B2(n_189),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_205),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_175),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_202),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_170),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_29),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_207),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_3),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_190),
.C(n_198),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_211),
.C(n_218),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_168),
.C(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_213),
.B(n_177),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_177),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_172),
.C(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_220),
.Y(n_231)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_185),
.C(n_186),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_224),
.C(n_207),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_185),
.C(n_174),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_216),
.A2(n_171),
.B(n_194),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_227),
.A2(n_208),
.B(n_214),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_222),
.Y(n_230)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_237),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_221),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_194),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_217),
.C(n_4),
.Y(n_247)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_218),
.CI(n_223),
.CON(n_238),
.SN(n_238)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_243),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_228),
.B(n_234),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_217),
.B1(n_4),
.B2(n_5),
.Y(n_243)
);

OA21x2_ASAP7_75t_SL g244 ( 
.A1(n_236),
.A2(n_229),
.B(n_231),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_238),
.B(n_245),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_247),
.B(n_3),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_249),
.B(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_228),
.C(n_4),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_251),
.B(n_252),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_5),
.B(n_7),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_255),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_240),
.B(n_7),
.Y(n_254)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_242),
.B1(n_238),
.B2(n_240),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_257),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_251),
.A2(n_242),
.B1(n_247),
.B2(n_243),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_245),
.C(n_249),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_262),
.B(n_264),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g263 ( 
.A1(n_258),
.A2(n_8),
.B(n_10),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_263),
.A2(n_11),
.B(n_12),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_8),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_11),
.C(n_12),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_261),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.C(n_264),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_271),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_259),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_265),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_13),
.B(n_14),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_14),
.B(n_15),
.Y(n_274)
);


endmodule