module fake_netlist_6_3793_n_1731 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1731);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1731;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1605;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_952;
wire n_725;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_69),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_173),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_186),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_57),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_179),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_78),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_165),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_21),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_21),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_54),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_133),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_22),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_127),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_14),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_83),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_6),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_3),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_71),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_161),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_131),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_14),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_97),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_74),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_84),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_142),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_115),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_56),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_26),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_130),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_35),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_36),
.Y(n_224)
);

BUFx8_ASAP7_75t_SL g225 ( 
.A(n_45),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_13),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_41),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_121),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_62),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_114),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_119),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_135),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_160),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_151),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_87),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_17),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_91),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_41),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_20),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_107),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_95),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_31),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_19),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_73),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_18),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_27),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_159),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_52),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_152),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_100),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_143),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_92),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_146),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_144),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_169),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_70),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_117),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_128),
.Y(n_258)
);

BUFx8_ASAP7_75t_SL g259 ( 
.A(n_118),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_43),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_11),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_180),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_40),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_79),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_167),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_5),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_58),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_26),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_182),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_75),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_164),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_132),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_112),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_62),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_99),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_66),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_1),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_57),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_19),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_58),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_23),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_108),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_1),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_86),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_177),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_16),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_153),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_120),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_17),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_18),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_65),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_10),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_38),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_181),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_7),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_157),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_4),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_27),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_166),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_126),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_39),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_101),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_6),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_82),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_52),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_34),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_183),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_96),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_12),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_3),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_93),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_185),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_102),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_134),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_28),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_36),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_104),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_72),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_67),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_170),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_156),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_47),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_88),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_109),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_85),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_24),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_184),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_24),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_106),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_5),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_4),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_89),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_64),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_38),
.Y(n_335)
);

BUFx8_ASAP7_75t_SL g336 ( 
.A(n_22),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_34),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_35),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_158),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_55),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_23),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_154),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_150),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_140),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_129),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_123),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_149),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_0),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_39),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_155),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_116),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_30),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_94),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_12),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_59),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_122),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_76),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_54),
.Y(n_358)
);

BUFx10_ASAP7_75t_L g359 ( 
.A(n_49),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_66),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_110),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_47),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_63),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_25),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_43),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_67),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_98),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_28),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_49),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_8),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_37),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_174),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_147),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_81),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_15),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_2),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_32),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_105),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_145),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_50),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_46),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_225),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_371),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_336),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_307),
.B(n_0),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_371),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_196),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_237),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_270),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_196),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_195),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_339),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_371),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_259),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_288),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_371),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_371),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_209),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_238),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_268),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_242),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_220),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_245),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_231),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_246),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_343),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_248),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_282),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_217),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_268),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_264),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_267),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_282),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_244),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_274),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_247),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_287),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_195),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_214),
.B(n_2),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_316),
.B(n_7),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_214),
.B(n_8),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_220),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_331),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_253),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_254),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_354),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_354),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_202),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_268),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_284),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_281),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_255),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_291),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_375),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_257),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_262),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_375),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_202),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_197),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_223),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_284),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_239),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_265),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_243),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_293),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_261),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_295),
.B(n_9),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_204),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_294),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_284),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_263),
.Y(n_452)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_341),
.B(n_10),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_269),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_359),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_266),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_275),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_224),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_277),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_296),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_359),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_278),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_306),
.Y(n_463)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_226),
.B(n_11),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_271),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_272),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_310),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_224),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_317),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_298),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_359),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_298),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_276),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_274),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_292),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_381),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_199),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_302),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_383),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_410),
.B(n_309),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_388),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_392),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_383),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_388),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_386),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_386),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_R g487 ( 
.A(n_400),
.B(n_187),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_389),
.B(n_190),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_226),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

AND2x2_ASAP7_75t_R g491 ( 
.A(n_477),
.B(n_311),
.Y(n_491)
);

OA21x2_ASAP7_75t_L g492 ( 
.A1(n_394),
.A2(n_398),
.B(n_397),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_410),
.B(n_309),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_388),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_431),
.B(n_199),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_395),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_422),
.A2(n_207),
.B(n_203),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_397),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_415),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_423),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_423),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_407),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_390),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_417),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_410),
.B(n_303),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_407),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_399),
.B(n_318),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_425),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_407),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_458),
.Y(n_513)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_382),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_407),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_407),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_416),
.B(n_303),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_426),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_433),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_475),
.Y(n_521)
);

OA21x2_ASAP7_75t_L g522 ( 
.A1(n_403),
.A2(n_470),
.B(n_468),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_436),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_416),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_448),
.A2(n_207),
.B(n_203),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_476),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_476),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_478),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_387),
.B(n_304),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_470),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_472),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_420),
.B(n_187),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_437),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_478),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_391),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_385),
.B(n_304),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_393),
.B(n_229),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_444),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_456),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_465),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_402),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_409),
.B(n_241),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_440),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_441),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_466),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_445),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_419),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_473),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_447),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_452),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_454),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_457),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_459),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_508),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_508),
.B(n_405),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_532),
.B(n_402),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_532),
.B(n_404),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_518),
.B(n_404),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_SL g560 ( 
.A(n_496),
.B(n_260),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_492),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_508),
.B(n_406),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_507),
.B(n_401),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_510),
.B(n_408),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_507),
.B(n_411),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_484),
.Y(n_566)
);

INVx3_ASAP7_75t_R g567 ( 
.A(n_541),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_535),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_481),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_518),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_481),
.Y(n_571)
);

INVx11_ASAP7_75t_L g572 ( 
.A(n_514),
.Y(n_572)
);

BUFx4f_ASAP7_75t_L g573 ( 
.A(n_541),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_484),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_489),
.B(n_408),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_482),
.B(n_439),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_524),
.B(n_414),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_524),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_543),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_489),
.B(n_412),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_492),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_543),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_482),
.B(n_430),
.Y(n_583)
);

OAI22xp33_ASAP7_75t_L g584 ( 
.A1(n_536),
.A2(n_363),
.B1(n_299),
.B2(n_206),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_524),
.Y(n_585)
);

OAI22xp33_ASAP7_75t_L g586 ( 
.A1(n_536),
.A2(n_206),
.B1(n_208),
.B2(n_204),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_L g587 ( 
.A(n_529),
.B(n_412),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_524),
.B(n_413),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_529),
.B(n_542),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_522),
.A2(n_464),
.B1(n_250),
.B2(n_258),
.Y(n_590)
);

AND2x2_ASAP7_75t_SL g591 ( 
.A(n_480),
.B(n_241),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_544),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_544),
.B(n_413),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_546),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_544),
.B(n_432),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_488),
.A2(n_327),
.B1(n_355),
.B2(n_290),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_484),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_544),
.B(n_250),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_547),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_548),
.B(n_439),
.Y(n_600)
);

INVxp33_ASAP7_75t_L g601 ( 
.A(n_548),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_481),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_536),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_544),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_480),
.B(n_432),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_536),
.B(n_442),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_488),
.Y(n_607)
);

NAND3xp33_ASAP7_75t_L g608 ( 
.A(n_487),
.B(n_446),
.C(n_434),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_484),
.Y(n_609)
);

INVx4_ASAP7_75t_SL g610 ( 
.A(n_490),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_547),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_542),
.B(n_418),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_536),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_550),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_550),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_554),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_536),
.A2(n_377),
.B1(n_208),
.B2(n_213),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_493),
.B(n_481),
.Y(n_618)
);

BUFx4f_ASAP7_75t_L g619 ( 
.A(n_544),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_493),
.B(n_429),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_554),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_553),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_553),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_490),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_553),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_553),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_492),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_553),
.B(n_434),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_492),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_553),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_517),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_490),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_542),
.B(n_258),
.Y(n_633)
);

INVx4_ASAP7_75t_SL g634 ( 
.A(n_490),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_485),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_494),
.B(n_446),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_479),
.B(n_450),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_522),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_494),
.B(n_450),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_517),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_551),
.B(n_460),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_494),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_521),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_479),
.B(n_460),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_522),
.A2(n_286),
.B1(n_335),
.B2(n_334),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_530),
.B(n_286),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_521),
.Y(n_647)
);

NAND3xp33_ASAP7_75t_L g648 ( 
.A(n_526),
.B(n_467),
.C(n_463),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_526),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_485),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_L g651 ( 
.A(n_527),
.B(n_463),
.Y(n_651)
);

AND2x6_ASAP7_75t_L g652 ( 
.A(n_528),
.B(n_343),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_490),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_494),
.B(n_467),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_522),
.A2(n_337),
.B1(n_332),
.B2(n_348),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_551),
.A2(n_396),
.B1(n_469),
.B2(n_455),
.Y(n_656)
);

AND2x6_ASAP7_75t_L g657 ( 
.A(n_528),
.B(n_343),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_551),
.B(n_469),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_552),
.B(n_451),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_495),
.Y(n_660)
);

OAI21xp33_ASAP7_75t_SL g661 ( 
.A1(n_499),
.A2(n_453),
.B(n_421),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_534),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_485),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_530),
.B(n_343),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_516),
.Y(n_665)
);

INVx5_ASAP7_75t_L g666 ( 
.A(n_490),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_483),
.B(n_449),
.Y(n_667)
);

AND2x6_ASAP7_75t_L g668 ( 
.A(n_534),
.B(n_353),
.Y(n_668)
);

BUFx4f_ASAP7_75t_L g669 ( 
.A(n_530),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_516),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_516),
.Y(n_671)
);

INVx4_ASAP7_75t_SL g672 ( 
.A(n_504),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_495),
.Y(n_673)
);

NOR3xp33_ASAP7_75t_L g674 ( 
.A(n_552),
.B(n_461),
.C(n_471),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_537),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_486),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_486),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_483),
.Y(n_678)
);

AO22x2_ASAP7_75t_L g679 ( 
.A1(n_491),
.A2(n_352),
.B1(n_358),
.B2(n_362),
.Y(n_679)
);

NOR2x1p5_ASAP7_75t_L g680 ( 
.A(n_501),
.B(n_382),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_504),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_504),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_509),
.Y(n_683)
);

INVx6_ASAP7_75t_L g684 ( 
.A(n_509),
.Y(n_684)
);

AND2x6_ASAP7_75t_L g685 ( 
.A(n_498),
.B(n_353),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_537),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_498),
.B(n_424),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_500),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_509),
.B(n_289),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_570),
.Y(n_690)
);

OR2x2_ASAP7_75t_SL g691 ( 
.A(n_608),
.B(n_564),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_590),
.B(n_531),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_590),
.A2(n_201),
.B1(n_351),
.B2(n_218),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_570),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_580),
.B(n_506),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_557),
.B(n_531),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_557),
.B(n_384),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_555),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_558),
.B(n_531),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_555),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_561),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_591),
.B(n_353),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_559),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_578),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_591),
.B(n_530),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_596),
.B(n_519),
.C(n_511),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_579),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_638),
.B(n_662),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_L g709 ( 
.A(n_651),
.B(n_575),
.C(n_648),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_582),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_629),
.Y(n_711)
);

NOR2xp67_ASAP7_75t_L g712 ( 
.A(n_585),
.B(n_520),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_576),
.Y(n_713)
);

OR2x6_ASAP7_75t_L g714 ( 
.A(n_563),
.B(n_427),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_605),
.B(n_384),
.Y(n_715)
);

AND2x2_ASAP7_75t_SL g716 ( 
.A(n_645),
.B(n_655),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_593),
.A2(n_308),
.B1(n_301),
.B2(n_300),
.Y(n_717)
);

AOI221xp5_ASAP7_75t_L g718 ( 
.A1(n_584),
.A2(n_279),
.B1(n_227),
.B2(n_219),
.C(n_213),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_600),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_561),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_629),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_620),
.B(n_523),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_638),
.A2(n_499),
.B1(n_525),
.B2(n_346),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_662),
.B(n_353),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_593),
.B(n_499),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_655),
.A2(n_525),
.B(n_370),
.C(n_364),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_589),
.B(n_525),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_581),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_581),
.B(n_221),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_595),
.B(n_228),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_627),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_583),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_562),
.B(n_533),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_659),
.Y(n_734)
);

INVx8_ASAP7_75t_L g735 ( 
.A(n_659),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_594),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_601),
.B(n_538),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_599),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_631),
.A2(n_249),
.B1(n_315),
.B2(n_313),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_572),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_595),
.B(n_230),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_628),
.B(n_232),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_628),
.B(n_240),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_649),
.B(n_618),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_611),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_614),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_641),
.A2(n_325),
.B1(n_319),
.B2(n_321),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_L g748 ( 
.A(n_603),
.B(n_251),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_615),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_616),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_661),
.B(n_256),
.Y(n_751)
);

AND2x6_ASAP7_75t_SL g752 ( 
.A(n_583),
.B(n_368),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_601),
.B(n_539),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_640),
.B(n_273),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_556),
.B(n_545),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_643),
.A2(n_633),
.B(n_587),
.C(n_667),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_658),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_577),
.B(n_283),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_647),
.B(n_285),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_621),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_635),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_643),
.Y(n_762)
);

OAI22xp33_ASAP7_75t_L g763 ( 
.A1(n_603),
.A2(n_305),
.B1(n_312),
.B2(n_324),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_577),
.B(n_326),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_667),
.A2(n_435),
.B(n_438),
.C(n_428),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_613),
.A2(n_328),
.B1(n_322),
.B2(n_330),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_568),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_612),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_650),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_636),
.B(n_374),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_678),
.B(n_500),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_588),
.B(n_540),
.Y(n_772)
);

OR2x2_ASAP7_75t_SL g773 ( 
.A(n_560),
.B(n_491),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_665),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_573),
.B(n_549),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_573),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_637),
.B(n_505),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_644),
.B(n_497),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_665),
.Y(n_779)
);

NOR2x1_ASAP7_75t_R g780 ( 
.A(n_607),
.B(n_188),
.Y(n_780)
);

OAI22xp33_ASAP7_75t_L g781 ( 
.A1(n_659),
.A2(n_219),
.B1(n_227),
.B2(n_236),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_612),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_639),
.B(n_188),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_583),
.B(n_462),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_633),
.A2(n_486),
.B1(n_297),
.B2(n_222),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_654),
.B(n_189),
.Y(n_786)
);

NAND2xp33_ASAP7_75t_L g787 ( 
.A(n_652),
.B(n_189),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_688),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_656),
.B(n_606),
.Y(n_789)
);

NAND3xp33_ASAP7_75t_L g790 ( 
.A(n_674),
.B(n_560),
.C(n_687),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_606),
.B(n_191),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_660),
.B(n_502),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_586),
.B(n_191),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_675),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_606),
.B(n_192),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_687),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_622),
.A2(n_345),
.B1(n_222),
.B2(n_252),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_663),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_673),
.B(n_502),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_683),
.B(n_503),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_586),
.B(n_192),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_623),
.A2(n_345),
.B1(n_222),
.B2(n_252),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_686),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_617),
.B(n_193),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_683),
.B(n_503),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_670),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_617),
.B(n_193),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_670),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_663),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_674),
.B(n_194),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_689),
.B(n_513),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_679),
.A2(n_194),
.B1(n_198),
.B2(n_333),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_676),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_569),
.B(n_68),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_571),
.B(n_198),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_619),
.A2(n_669),
.B(n_626),
.Y(n_816)
);

BUFx6f_ASAP7_75t_SL g817 ( 
.A(n_563),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_676),
.Y(n_818)
);

OAI221xp5_ASAP7_75t_L g819 ( 
.A1(n_646),
.A2(n_323),
.B1(n_329),
.B2(n_320),
.C(n_380),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_602),
.B(n_200),
.Y(n_820)
);

BUFx12f_ASAP7_75t_L g821 ( 
.A(n_680),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_642),
.B(n_200),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_679),
.A2(n_205),
.B1(n_210),
.B2(n_211),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_677),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_677),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_609),
.B(n_624),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_774),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_716),
.B(n_625),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_744),
.B(n_624),
.Y(n_829)
);

AOI21x1_ASAP7_75t_L g830 ( 
.A1(n_729),
.A2(n_630),
.B(n_671),
.Y(n_830)
);

BUFx12f_ASAP7_75t_L g831 ( 
.A(n_740),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_757),
.B(n_565),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_692),
.A2(n_592),
.B(n_604),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_693),
.A2(n_584),
.B(n_598),
.C(n_646),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_756),
.A2(n_664),
.B(n_356),
.C(n_350),
.Y(n_835)
);

CKINVDCx11_ASAP7_75t_R g836 ( 
.A(n_821),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_716),
.B(n_566),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_727),
.A2(n_664),
.B(n_653),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_709),
.A2(n_679),
.B1(n_565),
.B2(n_684),
.Y(n_839)
);

INVx11_ASAP7_75t_L g840 ( 
.A(n_821),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_774),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_703),
.B(n_567),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_765),
.A2(n_565),
.B(n_682),
.C(n_681),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_727),
.A2(n_682),
.B(n_681),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_768),
.B(n_610),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_761),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_729),
.A2(n_811),
.B(n_711),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_762),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_690),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_796),
.B(n_696),
.Y(n_850)
);

O2A1O1Ixp5_ASAP7_75t_L g851 ( 
.A1(n_751),
.A2(n_685),
.B(n_652),
.C(n_668),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_SL g852 ( 
.A1(n_702),
.A2(n_199),
.B(n_372),
.C(n_314),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_721),
.A2(n_357),
.B1(n_210),
.B2(n_211),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_711),
.A2(n_632),
.B(n_597),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_711),
.A2(n_632),
.B(n_597),
.Y(n_855)
);

AOI21xp33_ASAP7_75t_L g856 ( 
.A1(n_697),
.A2(n_279),
.B(n_236),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_774),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_694),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_699),
.B(n_610),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_792),
.A2(n_666),
.B(n_574),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_794),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_799),
.A2(n_666),
.B(n_574),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_702),
.A2(n_349),
.B1(n_280),
.B2(n_369),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_713),
.B(n_280),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_708),
.A2(n_205),
.B1(n_212),
.B2(n_215),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_800),
.A2(n_666),
.B(n_574),
.Y(n_866)
);

AO21x1_ASAP7_75t_L g867 ( 
.A1(n_751),
.A2(n_372),
.B(n_314),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_701),
.B(n_720),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_793),
.A2(n_372),
.B(n_297),
.C(n_314),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_805),
.A2(n_666),
.B(n_574),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_701),
.B(n_634),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_776),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_720),
.B(n_672),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_816),
.A2(n_708),
.B(n_705),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_728),
.B(n_672),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_728),
.B(n_216),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_755),
.A2(n_361),
.B1(n_233),
.B2(n_234),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_700),
.B(n_233),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_R g879 ( 
.A(n_778),
.B(n_234),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_826),
.A2(n_512),
.B(n_515),
.Y(n_880)
);

BUFx4f_ASAP7_75t_L g881 ( 
.A(n_735),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_700),
.B(n_731),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_731),
.B(n_235),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_784),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_691),
.A2(n_235),
.B1(n_333),
.B2(n_342),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_774),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_L g887 ( 
.A(n_804),
.B(n_379),
.C(n_378),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_700),
.B(n_342),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_790),
.A2(n_379),
.B(n_378),
.C(n_373),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_786),
.B(n_344),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_719),
.B(n_338),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_SL g892 ( 
.A1(n_726),
.A2(n_297),
.B(n_15),
.C(n_16),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_730),
.A2(n_367),
.B1(n_344),
.B2(n_347),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_769),
.Y(n_894)
);

BUFx8_ASAP7_75t_SL g895 ( 
.A(n_817),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_782),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_698),
.A2(n_367),
.B1(n_373),
.B2(n_357),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_742),
.A2(n_350),
.B1(n_356),
.B2(n_340),
.Y(n_898)
);

NOR2x1_ASAP7_75t_L g899 ( 
.A(n_712),
.B(n_340),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_743),
.A2(n_349),
.B(n_360),
.C(n_365),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_768),
.B(n_103),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_775),
.Y(n_902)
);

OR2x6_ASAP7_75t_L g903 ( 
.A(n_735),
.B(n_732),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_770),
.A2(n_657),
.B1(n_652),
.B2(n_380),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_695),
.B(n_360),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_806),
.A2(n_657),
.B(n_377),
.Y(n_906)
);

AND2x6_ASAP7_75t_SL g907 ( 
.A(n_737),
.B(n_376),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_806),
.A2(n_376),
.B(n_369),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_779),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_707),
.B(n_366),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_SL g911 ( 
.A(n_753),
.B(n_366),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_710),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_798),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_726),
.A2(n_175),
.B(n_171),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_779),
.B(n_163),
.Y(n_915)
);

NOR2x1p5_ASAP7_75t_SL g916 ( 
.A(n_798),
.B(n_162),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_736),
.B(n_13),
.Y(n_917)
);

OAI321xp33_ASAP7_75t_L g918 ( 
.A1(n_718),
.A2(n_25),
.A3(n_29),
.B1(n_30),
.B2(n_31),
.C(n_32),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_738),
.B(n_29),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_770),
.A2(n_139),
.B1(n_138),
.B2(n_137),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_745),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_733),
.B(n_33),
.Y(n_922)
);

AOI21x1_ASAP7_75t_L g923 ( 
.A1(n_741),
.A2(n_136),
.B(n_124),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_746),
.B(n_33),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_723),
.A2(n_113),
.B(n_111),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_734),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_704),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_777),
.B(n_37),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_749),
.B(n_42),
.Y(n_929)
);

O2A1O1Ixp5_ASAP7_75t_L g930 ( 
.A1(n_724),
.A2(n_42),
.B(n_44),
.C(n_45),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_715),
.B(n_44),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_758),
.A2(n_90),
.B(n_80),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_764),
.A2(n_77),
.B(n_48),
.Y(n_933)
);

AOI22x1_ASAP7_75t_L g934 ( 
.A1(n_767),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_814),
.B(n_51),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_724),
.A2(n_51),
.B(n_53),
.Y(n_936)
);

CKINVDCx10_ASAP7_75t_R g937 ( 
.A(n_817),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_793),
.A2(n_801),
.B(n_807),
.C(n_748),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_772),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_939)
);

BUFx12f_ASAP7_75t_L g940 ( 
.A(n_752),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_814),
.B(n_59),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_771),
.A2(n_825),
.B(n_824),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_809),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_750),
.A2(n_65),
.B1(n_61),
.B2(n_63),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_760),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_714),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_788),
.B(n_60),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_801),
.B(n_64),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_809),
.A2(n_60),
.B(n_61),
.Y(n_949)
);

CKINVDCx10_ASAP7_75t_R g950 ( 
.A(n_714),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_813),
.A2(n_818),
.B(n_783),
.Y(n_951)
);

NAND2x1p5_ASAP7_75t_L g952 ( 
.A(n_814),
.B(n_808),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_735),
.B(n_714),
.Y(n_953)
);

AOI21x1_ASAP7_75t_L g954 ( 
.A1(n_818),
.A2(n_754),
.B(n_759),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_SL g955 ( 
.A1(n_807),
.A2(n_763),
.B(n_810),
.C(n_783),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_808),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_704),
.Y(n_957)
);

CKINVDCx6p67_ASAP7_75t_R g958 ( 
.A(n_803),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_717),
.B(n_747),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_722),
.B(n_781),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_815),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_748),
.A2(n_820),
.B(n_822),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_810),
.B(n_789),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_735),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_812),
.B(n_823),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_766),
.B(n_795),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_787),
.A2(n_791),
.B(n_819),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_706),
.B(n_797),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_739),
.B(n_785),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_847),
.A2(n_787),
.B(n_802),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_850),
.B(n_780),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_837),
.A2(n_773),
.B(n_828),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_841),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_955),
.A2(n_938),
.B(n_922),
.C(n_948),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_837),
.A2(n_828),
.B(n_874),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_861),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_905),
.B(n_884),
.Y(n_977)
);

OA21x2_ASAP7_75t_L g978 ( 
.A1(n_914),
.A2(n_925),
.B(n_844),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_963),
.A2(n_922),
.B1(n_965),
.B2(n_966),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_958),
.Y(n_980)
);

AO21x1_ASAP7_75t_L g981 ( 
.A1(n_928),
.A2(n_948),
.B(n_966),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_931),
.B(n_961),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_965),
.A2(n_918),
.B(n_960),
.C(n_834),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_921),
.B(n_945),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_882),
.A2(n_835),
.B(n_962),
.Y(n_985)
);

AND2x2_ASAP7_75t_SL g986 ( 
.A(n_959),
.B(n_863),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_890),
.B(n_952),
.Y(n_987)
);

NAND2x1_ASAP7_75t_L g988 ( 
.A(n_857),
.B(n_841),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_952),
.B(n_829),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_856),
.B(n_960),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_868),
.A2(n_941),
.B(n_935),
.Y(n_991)
);

NAND2x1p5_ASAP7_75t_L g992 ( 
.A(n_964),
.B(n_857),
.Y(n_992)
);

AO21x1_ASAP7_75t_L g993 ( 
.A1(n_843),
.A2(n_941),
.B(n_935),
.Y(n_993)
);

OA21x2_ASAP7_75t_L g994 ( 
.A1(n_838),
.A2(n_942),
.B(n_954),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_896),
.B(n_863),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_896),
.B(n_849),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_854),
.A2(n_855),
.B(n_880),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_831),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_968),
.A2(n_911),
.B1(n_839),
.B2(n_888),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_858),
.B(n_876),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_SL g1001 ( 
.A(n_872),
.B(n_964),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_841),
.Y(n_1002)
);

AOI21x1_ASAP7_75t_L g1003 ( 
.A1(n_878),
.A2(n_888),
.B(n_860),
.Y(n_1003)
);

OAI22x1_ASAP7_75t_L g1004 ( 
.A1(n_939),
.A2(n_934),
.B1(n_927),
.B2(n_926),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_SL g1005 ( 
.A1(n_923),
.A2(n_933),
.B(n_932),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_841),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_L g1007 ( 
.A(n_877),
.B(n_887),
.C(n_864),
.Y(n_1007)
);

AO31x2_ASAP7_75t_L g1008 ( 
.A1(n_867),
.A2(n_889),
.A3(n_900),
.B(n_949),
.Y(n_1008)
);

AND2x2_ASAP7_75t_SL g1009 ( 
.A(n_881),
.B(n_915),
.Y(n_1009)
);

OR2x6_ASAP7_75t_L g1010 ( 
.A(n_953),
.B(n_903),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_871),
.A2(n_875),
.B(n_873),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_862),
.A2(n_870),
.B(n_866),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_955),
.A2(n_878),
.B(n_969),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_883),
.A2(n_846),
.B(n_894),
.Y(n_1014)
);

OAI21xp33_ASAP7_75t_L g1015 ( 
.A1(n_879),
.A2(n_864),
.B(n_891),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_881),
.Y(n_1016)
);

AOI21xp33_ASAP7_75t_L g1017 ( 
.A1(n_869),
.A2(n_891),
.B(n_910),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_848),
.B(n_927),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_836),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_930),
.A2(n_936),
.B(n_924),
.C(n_917),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_956),
.B(n_947),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_902),
.B(n_957),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_886),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_957),
.B(n_832),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_913),
.A2(n_943),
.B(n_929),
.Y(n_1025)
);

NOR2x1_ASAP7_75t_SL g1026 ( 
.A(n_886),
.B(n_909),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_851),
.A2(n_906),
.B(n_919),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_901),
.A2(n_909),
.B1(n_886),
.B2(n_827),
.Y(n_1028)
);

INVx3_ASAP7_75t_SL g1029 ( 
.A(n_953),
.Y(n_1029)
);

INVx6_ASAP7_75t_L g1030 ( 
.A(n_886),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_845),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_946),
.Y(n_1032)
);

AO31x2_ASAP7_75t_L g1033 ( 
.A1(n_944),
.A2(n_885),
.A3(n_898),
.B(n_893),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_930),
.A2(n_920),
.B(n_908),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_853),
.A2(n_865),
.B(n_897),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_899),
.A2(n_916),
.B(n_904),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_909),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_879),
.B(n_842),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_909),
.B(n_845),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_892),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_892),
.A2(n_852),
.B(n_842),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_903),
.A2(n_953),
.B(n_840),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_903),
.B(n_907),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_940),
.B(n_950),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_895),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_937),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_912),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_837),
.A2(n_828),
.B(n_874),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_861),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_837),
.A2(n_828),
.B(n_874),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_912),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_850),
.B(n_744),
.Y(n_1052)
);

AOI21x1_ASAP7_75t_SL g1053 ( 
.A1(n_859),
.A2(n_959),
.B(n_725),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_830),
.A2(n_951),
.B(n_833),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_841),
.Y(n_1055)
);

OR2x6_ASAP7_75t_L g1056 ( 
.A(n_953),
.B(n_735),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_850),
.B(n_744),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_850),
.B(n_744),
.Y(n_1058)
);

O2A1O1Ixp5_ASAP7_75t_L g1059 ( 
.A1(n_922),
.A2(n_741),
.B(n_925),
.C(n_751),
.Y(n_1059)
);

AND3x4_ASAP7_75t_L g1060 ( 
.A(n_946),
.B(n_706),
.C(n_674),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_830),
.A2(n_951),
.B(n_833),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_905),
.B(n_580),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_948),
.A2(n_716),
.B(n_938),
.C(n_922),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_850),
.B(n_744),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_850),
.B(n_744),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_841),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_948),
.A2(n_716),
.B(n_938),
.C(n_922),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_905),
.B(n_580),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_850),
.B(n_744),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_912),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_964),
.B(n_957),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_830),
.A2(n_951),
.B(n_833),
.Y(n_1072)
);

AOI221x1_ASAP7_75t_L g1073 ( 
.A1(n_922),
.A2(n_963),
.B1(n_928),
.B2(n_967),
.C(n_914),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_964),
.B(n_957),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_830),
.A2(n_951),
.B(n_833),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_850),
.B(n_744),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_912),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_830),
.A2(n_951),
.B(n_833),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_905),
.B(n_580),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_837),
.A2(n_828),
.B(n_874),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_850),
.B(n_744),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_959),
.B(n_716),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_963),
.B(n_777),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_837),
.A2(n_828),
.B(n_874),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_850),
.B(n_744),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_830),
.A2(n_951),
.B(n_833),
.Y(n_1086)
);

OAI22x1_ASAP7_75t_L g1087 ( 
.A1(n_928),
.A2(n_965),
.B1(n_963),
.B2(n_804),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_850),
.B(n_744),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_964),
.B(n_957),
.Y(n_1089)
);

NOR2x1_ASAP7_75t_L g1090 ( 
.A(n_861),
.B(n_709),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_948),
.A2(n_716),
.B(n_938),
.C(n_922),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_850),
.B(n_744),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_837),
.A2(n_828),
.B(n_874),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_1016),
.B(n_1010),
.Y(n_1094)
);

BUFx12f_ASAP7_75t_L g1095 ( 
.A(n_1019),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_1016),
.B(n_1010),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_1018),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_979),
.A2(n_983),
.B1(n_1058),
.B2(n_1064),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1083),
.B(n_1062),
.Y(n_1099)
);

BUFx4_ASAP7_75t_SL g1100 ( 
.A(n_976),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_1083),
.B(n_990),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_998),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1051),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1065),
.B(n_1069),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1010),
.B(n_1056),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1068),
.B(n_1079),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_990),
.B(n_1015),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1076),
.B(n_1081),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_SL g1109 ( 
.A1(n_986),
.A2(n_1007),
.B1(n_1035),
.B2(n_1001),
.Y(n_1109)
);

BUFx8_ASAP7_75t_SL g1110 ( 
.A(n_1046),
.Y(n_1110)
);

BUFx2_ASAP7_75t_R g1111 ( 
.A(n_1049),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1056),
.B(n_1042),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1085),
.B(n_1088),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1070),
.Y(n_1114)
);

BUFx8_ASAP7_75t_L g1115 ( 
.A(n_980),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_1002),
.Y(n_1116)
);

O2A1O1Ixp5_ASAP7_75t_SL g1117 ( 
.A1(n_1017),
.A2(n_1040),
.B(n_1082),
.C(n_985),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_SL g1118 ( 
.A(n_983),
.B(n_986),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_1073),
.B(n_974),
.C(n_1067),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_971),
.B(n_1092),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1002),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1056),
.B(n_1031),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1071),
.Y(n_1123)
);

BUFx4f_ASAP7_75t_SL g1124 ( 
.A(n_1029),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1071),
.B(n_1074),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1074),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1063),
.A2(n_1067),
.B1(n_1091),
.B2(n_999),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_SL g1128 ( 
.A(n_1045),
.B(n_1044),
.Y(n_1128)
);

AOI21xp33_ASAP7_75t_L g1129 ( 
.A1(n_1087),
.A2(n_974),
.B(n_981),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1077),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_977),
.B(n_1038),
.Y(n_1131)
);

INVx6_ASAP7_75t_L g1132 ( 
.A(n_1089),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1063),
.A2(n_1091),
.B(n_1059),
.C(n_1013),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_1032),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_995),
.B(n_1082),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1089),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_1024),
.B(n_1022),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1013),
.A2(n_991),
.B(n_970),
.C(n_972),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_982),
.A2(n_1020),
.B(n_1000),
.C(n_1041),
.Y(n_1139)
);

NAND2xp33_ASAP7_75t_L g1140 ( 
.A(n_987),
.B(n_984),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1090),
.Y(n_1141)
);

BUFx8_ASAP7_75t_L g1142 ( 
.A(n_1002),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1039),
.B(n_996),
.Y(n_1143)
);

OR2x2_ASAP7_75t_L g1144 ( 
.A(n_1021),
.B(n_1043),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_1029),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_991),
.B(n_989),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_973),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_L g1148 ( 
.A(n_1020),
.B(n_1041),
.C(n_978),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_993),
.B(n_1093),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_975),
.B(n_1048),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1060),
.A2(n_1004),
.B1(n_1084),
.B2(n_1080),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1037),
.B(n_1066),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1009),
.A2(n_1060),
.B1(n_1028),
.B2(n_1050),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1030),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1037),
.B(n_1066),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_1033),
.B(n_1008),
.Y(n_1156)
);

BUFx12f_ASAP7_75t_L g1157 ( 
.A(n_1030),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_973),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1009),
.A2(n_1034),
.B1(n_1014),
.B2(n_1027),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1006),
.B(n_1023),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1025),
.B(n_1033),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1006),
.Y(n_1162)
);

OR2x6_ASAP7_75t_L g1163 ( 
.A(n_992),
.B(n_988),
.Y(n_1163)
);

BUFx4f_ASAP7_75t_L g1164 ( 
.A(n_992),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1003),
.B(n_1055),
.Y(n_1165)
);

INVx1_ASAP7_75t_SL g1166 ( 
.A(n_1030),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1005),
.A2(n_1044),
.B(n_1055),
.C(n_994),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1026),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_994),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_L g1170 ( 
.A(n_1033),
.B(n_1053),
.C(n_1008),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1008),
.B(n_1036),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1011),
.Y(n_1172)
);

BUFx4_ASAP7_75t_SL g1173 ( 
.A(n_1053),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_997),
.B(n_1061),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1012),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_1054),
.Y(n_1176)
);

AOI21xp33_ASAP7_75t_SL g1177 ( 
.A1(n_1072),
.A2(n_1075),
.B(n_1078),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1086),
.A2(n_990),
.B1(n_1083),
.B2(n_777),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1073),
.A2(n_1067),
.B(n_1063),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1052),
.B(n_1057),
.Y(n_1180)
);

NOR2xp67_ASAP7_75t_L g1181 ( 
.A(n_971),
.B(n_740),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1016),
.B(n_1010),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_1018),
.B(n_803),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1083),
.B(n_1062),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1018),
.B(n_803),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_976),
.Y(n_1186)
);

NAND2xp33_ASAP7_75t_L g1187 ( 
.A(n_979),
.B(n_983),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1016),
.B(n_1010),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1083),
.B(n_1062),
.Y(n_1189)
);

OAI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_979),
.A2(n_1083),
.B1(n_990),
.B2(n_911),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1047),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1018),
.B(n_803),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1016),
.B(n_1010),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1047),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1016),
.B(n_1010),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1083),
.B(n_1062),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_979),
.A2(n_983),
.B1(n_716),
.B2(n_1052),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1083),
.B(n_1085),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1052),
.B(n_1057),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_SL g1200 ( 
.A1(n_990),
.A2(n_922),
.B(n_697),
.C(n_928),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1047),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1083),
.B(n_1062),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_979),
.B(n_573),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1019),
.Y(n_1204)
);

NOR2x1_ASAP7_75t_L g1205 ( 
.A(n_976),
.B(n_861),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1018),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_976),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1071),
.Y(n_1208)
);

INVx6_ASAP7_75t_L g1209 ( 
.A(n_976),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1052),
.B(n_1057),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_976),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1083),
.B(n_1085),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_976),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1083),
.B(n_1085),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1016),
.B(n_1010),
.Y(n_1215)
);

INVx4_ASAP7_75t_L g1216 ( 
.A(n_1002),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1016),
.B(n_1010),
.Y(n_1217)
);

OAI321xp33_ASAP7_75t_L g1218 ( 
.A1(n_979),
.A2(n_990),
.A3(n_1083),
.B1(n_922),
.B2(n_948),
.C(n_983),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1201),
.Y(n_1219)
);

NAND2x1p5_ASAP7_75t_L g1220 ( 
.A(n_1164),
.B(n_1105),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1103),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1114),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1190),
.A2(n_1187),
.B1(n_1109),
.B2(n_1107),
.Y(n_1223)
);

CKINVDCx11_ASAP7_75t_R g1224 ( 
.A(n_1095),
.Y(n_1224)
);

INVx6_ASAP7_75t_L g1225 ( 
.A(n_1142),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1097),
.Y(n_1226)
);

NAND2x1p5_ASAP7_75t_L g1227 ( 
.A(n_1164),
.B(n_1105),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1191),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1194),
.Y(n_1229)
);

BUFx12f_ASAP7_75t_L g1230 ( 
.A(n_1102),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1100),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1118),
.A2(n_1127),
.B1(n_1203),
.B2(n_1120),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_1183),
.Y(n_1233)
);

INVx6_ASAP7_75t_L g1234 ( 
.A(n_1142),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1198),
.B(n_1212),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1169),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1204),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_SL g1238 ( 
.A1(n_1118),
.A2(n_1127),
.B1(n_1153),
.B2(n_1197),
.Y(n_1238)
);

OAI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1214),
.A2(n_1218),
.B1(n_1113),
.B2(n_1178),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1104),
.B(n_1108),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_SL g1241 ( 
.A(n_1111),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1169),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1143),
.Y(n_1243)
);

INVx4_ASAP7_75t_L g1244 ( 
.A(n_1157),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1185),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_1192),
.Y(n_1246)
);

NAND2x1_ASAP7_75t_L g1247 ( 
.A(n_1112),
.B(n_1172),
.Y(n_1247)
);

OAI21xp33_ASAP7_75t_L g1248 ( 
.A1(n_1108),
.A2(n_1210),
.B(n_1199),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1143),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1121),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1153),
.A2(n_1197),
.B1(n_1098),
.B2(n_1141),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1206),
.Y(n_1252)
);

BUFx10_ASAP7_75t_L g1253 ( 
.A(n_1209),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1147),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1158),
.Y(n_1255)
);

AO21x1_ASAP7_75t_L g1256 ( 
.A1(n_1129),
.A2(n_1098),
.B(n_1179),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1180),
.A2(n_1210),
.B1(n_1199),
.B2(n_1151),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_SL g1258 ( 
.A1(n_1167),
.A2(n_1139),
.B(n_1135),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1162),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1099),
.A2(n_1189),
.B1(n_1196),
.B2(n_1202),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1218),
.A2(n_1200),
.B(n_1180),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1146),
.Y(n_1262)
);

CKINVDCx6p67_ASAP7_75t_R g1263 ( 
.A(n_1211),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1184),
.B(n_1179),
.Y(n_1264)
);

AO21x1_ASAP7_75t_L g1265 ( 
.A1(n_1129),
.A2(n_1149),
.B(n_1161),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1144),
.A2(n_1131),
.B1(n_1137),
.B2(n_1119),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1156),
.B(n_1137),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1106),
.B(n_1140),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_1209),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_1134),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1119),
.B(n_1161),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1117),
.A2(n_1171),
.B(n_1174),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1160),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1154),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1150),
.A2(n_1149),
.B(n_1138),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1121),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1168),
.Y(n_1277)
);

BUFx2_ASAP7_75t_R g1278 ( 
.A(n_1110),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1177),
.A2(n_1170),
.B(n_1148),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1186),
.A2(n_1213),
.B1(n_1207),
.B2(n_1128),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1124),
.A2(n_1181),
.B1(n_1145),
.B2(n_1150),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1205),
.A2(n_1217),
.B1(n_1096),
.B2(n_1193),
.Y(n_1282)
);

CKINVDCx16_ASAP7_75t_R g1283 ( 
.A(n_1094),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1133),
.B(n_1122),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1121),
.Y(n_1285)
);

OAI222xp33_ASAP7_75t_L g1286 ( 
.A1(n_1159),
.A2(n_1217),
.B1(n_1096),
.B2(n_1182),
.C1(n_1188),
.C2(n_1193),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1094),
.A2(n_1215),
.B1(n_1182),
.B2(n_1188),
.Y(n_1287)
);

BUFx2_ASAP7_75t_R g1288 ( 
.A(n_1123),
.Y(n_1288)
);

NAND2x1p5_ASAP7_75t_L g1289 ( 
.A(n_1195),
.B(n_1215),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1165),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1176),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_SL g1292 ( 
.A(n_1195),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1123),
.B(n_1136),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1148),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1170),
.A2(n_1163),
.B(n_1208),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_SL g1296 ( 
.A1(n_1116),
.A2(n_1216),
.B(n_1173),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1126),
.B(n_1208),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1125),
.Y(n_1298)
);

CKINVDCx11_ASAP7_75t_R g1299 ( 
.A(n_1166),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1116),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1132),
.A2(n_1163),
.B1(n_1152),
.B2(n_1155),
.Y(n_1301)
);

BUFx4f_ASAP7_75t_SL g1302 ( 
.A(n_1115),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1115),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1132),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1163),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1175),
.B(n_1198),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1097),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1135),
.B(n_1156),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1118),
.A2(n_1083),
.B1(n_990),
.B2(n_777),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1097),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1218),
.A2(n_1083),
.B(n_990),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1100),
.Y(n_1312)
);

BUFx12f_ASAP7_75t_L g1313 ( 
.A(n_1095),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1101),
.B(n_986),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1130),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1101),
.A2(n_979),
.B1(n_1083),
.B2(n_990),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1130),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1097),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1130),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1190),
.A2(n_990),
.B1(n_1083),
.B2(n_986),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1135),
.B(n_1156),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1164),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1118),
.A2(n_1083),
.B1(n_990),
.B2(n_777),
.Y(n_1323)
);

CKINVDCx6p67_ASAP7_75t_R g1324 ( 
.A(n_1095),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1264),
.B(n_1314),
.Y(n_1325)
);

NAND3xp33_ASAP7_75t_L g1326 ( 
.A(n_1309),
.B(n_1323),
.C(n_1311),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1233),
.B(n_1245),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1271),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1253),
.Y(n_1329)
);

NOR2x1_ASAP7_75t_R g1330 ( 
.A(n_1231),
.B(n_1312),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1271),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1308),
.B(n_1321),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1252),
.Y(n_1333)
);

INVx4_ASAP7_75t_L g1334 ( 
.A(n_1322),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1236),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1242),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1242),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1294),
.Y(n_1338)
);

BUFx10_ASAP7_75t_L g1339 ( 
.A(n_1231),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1267),
.B(n_1238),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1295),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1308),
.B(n_1321),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1294),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1290),
.B(n_1266),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1262),
.B(n_1275),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_1226),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1265),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1265),
.Y(n_1348)
);

BUFx12f_ASAP7_75t_L g1349 ( 
.A(n_1224),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1284),
.B(n_1251),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1247),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1240),
.B(n_1248),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1235),
.B(n_1316),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1261),
.B(n_1256),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1306),
.B(n_1291),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1256),
.B(n_1232),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1307),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1258),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1320),
.B(n_1315),
.Y(n_1359)
);

INVx5_ASAP7_75t_SL g1360 ( 
.A(n_1263),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1272),
.A2(n_1223),
.B(n_1277),
.Y(n_1361)
);

AO21x2_ASAP7_75t_L g1362 ( 
.A1(n_1279),
.A2(n_1272),
.B(n_1239),
.Y(n_1362)
);

AO21x2_ASAP7_75t_L g1363 ( 
.A1(n_1279),
.A2(n_1305),
.B(n_1257),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1322),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1221),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1222),
.A2(n_1228),
.B(n_1229),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1310),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1246),
.B(n_1260),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1237),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1253),
.Y(n_1370)
);

OR2x6_ASAP7_75t_L g1371 ( 
.A(n_1220),
.B(n_1227),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1243),
.A2(n_1249),
.B(n_1268),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1310),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1318),
.B(n_1219),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1296),
.A2(n_1322),
.B(n_1220),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1286),
.A2(n_1319),
.B(n_1317),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1299),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1293),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1301),
.A2(n_1281),
.B(n_1289),
.Y(n_1379)
);

BUFx5_ASAP7_75t_L g1380 ( 
.A(n_1297),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1254),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1255),
.Y(n_1382)
);

BUFx10_ASAP7_75t_L g1383 ( 
.A(n_1312),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1259),
.Y(n_1384)
);

INVxp33_ASAP7_75t_L g1385 ( 
.A(n_1270),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1273),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1287),
.B(n_1298),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1298),
.B(n_1283),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1300),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1285),
.B(n_1282),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1372),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1328),
.B(n_1280),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1328),
.B(n_1250),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1325),
.B(n_1331),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1331),
.B(n_1263),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1332),
.B(n_1274),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1366),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1375),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1366),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1371),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1366),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1372),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1365),
.Y(n_1403)
);

OAI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1326),
.A2(n_1269),
.B1(n_1304),
.B2(n_1244),
.C(n_1234),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1354),
.B(n_1250),
.Y(n_1405)
);

AND2x2_ASAP7_75t_SL g1406 ( 
.A(n_1356),
.B(n_1288),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1365),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1372),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1332),
.B(n_1276),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1372),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1356),
.A2(n_1292),
.B1(n_1299),
.B2(n_1324),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1375),
.Y(n_1412)
);

INVxp67_ASAP7_75t_SL g1413 ( 
.A(n_1345),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1342),
.B(n_1276),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1357),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1346),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1351),
.B(n_1244),
.Y(n_1417)
);

NOR2x2_ASAP7_75t_L g1418 ( 
.A(n_1371),
.B(n_1302),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1363),
.B(n_1225),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1371),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1367),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1363),
.B(n_1234),
.Y(n_1422)
);

NOR2x1_ASAP7_75t_L g1423 ( 
.A(n_1358),
.B(n_1241),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1342),
.B(n_1234),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1335),
.B(n_1234),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1333),
.B(n_1237),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1363),
.B(n_1324),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1378),
.B(n_1303),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1378),
.B(n_1313),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1409),
.B(n_1367),
.Y(n_1430)
);

OAI221xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1411),
.A2(n_1350),
.B1(n_1353),
.B2(n_1341),
.C(n_1379),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1414),
.B(n_1355),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1406),
.B(n_1427),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1427),
.A2(n_1358),
.B(n_1352),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1395),
.B(n_1341),
.Y(n_1435)
);

NAND3xp33_ASAP7_75t_L g1436 ( 
.A(n_1392),
.B(n_1404),
.C(n_1424),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_L g1437 ( 
.A(n_1392),
.B(n_1344),
.C(n_1347),
.Y(n_1437)
);

NAND3xp33_ASAP7_75t_L g1438 ( 
.A(n_1424),
.B(n_1344),
.C(n_1347),
.Y(n_1438)
);

OAI221xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1395),
.A2(n_1350),
.B1(n_1368),
.B2(n_1340),
.C(n_1348),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1406),
.A2(n_1371),
.B1(n_1340),
.B2(n_1359),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1413),
.B(n_1374),
.Y(n_1441)
);

OAI21xp33_ASAP7_75t_L g1442 ( 
.A1(n_1406),
.A2(n_1390),
.B(n_1359),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_L g1443 ( 
.A(n_1419),
.B(n_1348),
.C(n_1390),
.Y(n_1443)
);

NAND4xp25_ASAP7_75t_L g1444 ( 
.A(n_1396),
.B(n_1327),
.C(n_1384),
.D(n_1374),
.Y(n_1444)
);

AND2x2_ASAP7_75t_SL g1445 ( 
.A(n_1400),
.B(n_1361),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1419),
.B(n_1376),
.C(n_1361),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1423),
.A2(n_1377),
.B(n_1388),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_L g1448 ( 
.A(n_1422),
.B(n_1376),
.C(n_1361),
.Y(n_1448)
);

NAND3xp33_ASAP7_75t_L g1449 ( 
.A(n_1422),
.B(n_1376),
.C(n_1361),
.Y(n_1449)
);

OAI21xp33_ASAP7_75t_L g1450 ( 
.A1(n_1425),
.A2(n_1385),
.B(n_1387),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1417),
.B(n_1373),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1420),
.B(n_1380),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1420),
.B(n_1380),
.Y(n_1453)
);

NAND4xp25_ASAP7_75t_L g1454 ( 
.A(n_1426),
.B(n_1384),
.C(n_1381),
.D(n_1382),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1394),
.B(n_1388),
.Y(n_1455)
);

NAND3xp33_ASAP7_75t_L g1456 ( 
.A(n_1397),
.B(n_1386),
.C(n_1343),
.Y(n_1456)
);

NAND2xp33_ASAP7_75t_SL g1457 ( 
.A(n_1420),
.B(n_1369),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1429),
.A2(n_1349),
.B1(n_1362),
.B2(n_1360),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1403),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1417),
.B(n_1389),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_SL g1461 ( 
.A1(n_1418),
.A2(n_1369),
.B1(n_1313),
.B2(n_1230),
.Y(n_1461)
);

NAND3xp33_ASAP7_75t_L g1462 ( 
.A(n_1397),
.B(n_1401),
.C(n_1399),
.Y(n_1462)
);

NAND3xp33_ASAP7_75t_L g1463 ( 
.A(n_1399),
.B(n_1386),
.C(n_1343),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1405),
.B(n_1338),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1416),
.B(n_1338),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1416),
.B(n_1336),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1393),
.B(n_1337),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1420),
.B(n_1380),
.Y(n_1468)
);

NOR3xp33_ASAP7_75t_L g1469 ( 
.A(n_1417),
.B(n_1334),
.C(n_1364),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1415),
.B(n_1421),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1459),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1462),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1466),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1452),
.B(n_1412),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1467),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1441),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1455),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1465),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1456),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1470),
.B(n_1391),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1463),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1430),
.B(n_1443),
.Y(n_1482)
);

NAND2xp33_ASAP7_75t_R g1483 ( 
.A(n_1435),
.B(n_1428),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1432),
.B(n_1402),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1464),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1452),
.B(n_1408),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1438),
.B(n_1408),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1457),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1454),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1453),
.B(n_1410),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1453),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1468),
.B(n_1410),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1468),
.B(n_1401),
.Y(n_1493)
);

NOR2x1_ASAP7_75t_L g1494 ( 
.A(n_1447),
.B(n_1412),
.Y(n_1494)
);

NAND2x1_ASAP7_75t_L g1495 ( 
.A(n_1437),
.B(n_1398),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1446),
.B(n_1362),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1445),
.B(n_1412),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1460),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1445),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1461),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1435),
.B(n_1450),
.Y(n_1501)
);

INVx5_ASAP7_75t_L g1502 ( 
.A(n_1457),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1451),
.B(n_1398),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1469),
.B(n_1398),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1472),
.B(n_1479),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1486),
.B(n_1499),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1471),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1493),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1471),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1487),
.B(n_1448),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1493),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1487),
.B(n_1472),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1479),
.B(n_1481),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1476),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1481),
.B(n_1449),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1497),
.B(n_1458),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1482),
.B(n_1434),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1497),
.B(n_1458),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1474),
.B(n_1460),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1476),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1490),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_SL g1522 ( 
.A(n_1502),
.B(n_1431),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1475),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1474),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1475),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1490),
.B(n_1444),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1474),
.B(n_1480),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1502),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1492),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1502),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1492),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1496),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1482),
.B(n_1436),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1496),
.Y(n_1534)
);

INVx3_ASAP7_75t_SL g1535 ( 
.A(n_1502),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1491),
.Y(n_1536)
);

INVxp33_ASAP7_75t_L g1537 ( 
.A(n_1501),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1473),
.B(n_1403),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1485),
.B(n_1407),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1507),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1533),
.B(n_1489),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1536),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1527),
.B(n_1494),
.Y(n_1543)
);

OAI32xp33_ASAP7_75t_L g1544 ( 
.A1(n_1533),
.A2(n_1483),
.A3(n_1433),
.B1(n_1500),
.B2(n_1442),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1507),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1528),
.Y(n_1546)
);

AOI21xp33_ASAP7_75t_L g1547 ( 
.A1(n_1515),
.A2(n_1495),
.B(n_1488),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1509),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1509),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1515),
.B(n_1484),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1505),
.B(n_1498),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1505),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1514),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1514),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1520),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1520),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1523),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1513),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1515),
.B(n_1495),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1513),
.B(n_1478),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1537),
.B(n_1517),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1538),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1513),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1535),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1528),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1528),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1517),
.A2(n_1433),
.B(n_1440),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1538),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1539),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1527),
.B(n_1503),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1512),
.B(n_1485),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1539),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1530),
.B(n_1504),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1536),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1527),
.B(n_1503),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1536),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1523),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1525),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1525),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1524),
.B(n_1488),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1526),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1524),
.B(n_1504),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1524),
.B(n_1516),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1512),
.B(n_1477),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1526),
.B(n_1498),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1581),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1543),
.B(n_1524),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1583),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1541),
.B(n_1516),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1540),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1543),
.B(n_1524),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1550),
.B(n_1512),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1540),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1580),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1564),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1553),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1553),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1552),
.B(n_1522),
.C(n_1510),
.Y(n_1598)
);

CKINVDCx16_ASAP7_75t_R g1599 ( 
.A(n_1546),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1561),
.B(n_1567),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1554),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1550),
.B(n_1526),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1554),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1556),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1583),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1551),
.B(n_1558),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1560),
.B(n_1563),
.Y(n_1607)
);

INVxp67_ASAP7_75t_SL g1608 ( 
.A(n_1565),
.Y(n_1608)
);

NAND2xp33_ASAP7_75t_L g1609 ( 
.A(n_1559),
.B(n_1502),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1585),
.B(n_1516),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1570),
.B(n_1518),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1556),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1557),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1570),
.B(n_1518),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1575),
.B(n_1518),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1575),
.B(n_1506),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1557),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1577),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1565),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1577),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1564),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1565),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1545),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1586),
.B(n_1560),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1621),
.Y(n_1625)
);

OAI322xp33_ASAP7_75t_L g1626 ( 
.A1(n_1600),
.A2(n_1510),
.A3(n_1559),
.B1(n_1522),
.B2(n_1534),
.C1(n_1532),
.C2(n_1571),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1595),
.B(n_1580),
.Y(n_1627)
);

OAI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1598),
.A2(n_1599),
.B1(n_1589),
.B2(n_1535),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1621),
.B(n_1562),
.Y(n_1629)
);

OAI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1610),
.A2(n_1609),
.B1(n_1606),
.B2(n_1547),
.C(n_1594),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1599),
.B(n_1500),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1611),
.B(n_1519),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1611),
.B(n_1568),
.Y(n_1633)
);

AO32x1_ASAP7_75t_L g1634 ( 
.A1(n_1619),
.A2(n_1566),
.A3(n_1530),
.B1(n_1582),
.B2(n_1542),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1590),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1590),
.Y(n_1636)
);

OAI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1602),
.A2(n_1535),
.B1(n_1510),
.B2(n_1530),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1593),
.Y(n_1638)
);

NOR2x1_ASAP7_75t_L g1639 ( 
.A(n_1592),
.B(n_1546),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1593),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1588),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1596),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1602),
.A2(n_1544),
.B(n_1573),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1614),
.B(n_1569),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1607),
.A2(n_1544),
.B(n_1573),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1608),
.Y(n_1646)
);

CKINVDCx14_ASAP7_75t_R g1647 ( 
.A(n_1605),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1596),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1614),
.B(n_1572),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_SL g1650 ( 
.A1(n_1607),
.A2(n_1566),
.B(n_1573),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1597),
.Y(n_1651)
);

AOI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1615),
.A2(n_1532),
.B1(n_1534),
.B2(n_1439),
.C(n_1578),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1639),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1641),
.B(n_1592),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1641),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1631),
.B(n_1615),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1635),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1634),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1625),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1624),
.B(n_1623),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1646),
.B(n_1623),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1627),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1636),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1647),
.B(n_1616),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1638),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1646),
.B(n_1616),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1650),
.B(n_1587),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1645),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1632),
.B(n_1587),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1634),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1630),
.B(n_1278),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1643),
.B(n_1591),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1628),
.A2(n_1591),
.B1(n_1584),
.B2(n_1619),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1668),
.A2(n_1628),
.B(n_1626),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1656),
.B(n_1629),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1668),
.A2(n_1634),
.B(n_1637),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1671),
.A2(n_1633),
.B1(n_1649),
.B2(n_1644),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1654),
.Y(n_1678)
);

OAI211xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1662),
.A2(n_1652),
.B(n_1651),
.C(n_1648),
.Y(n_1679)
);

AOI221x1_ASAP7_75t_L g1680 ( 
.A1(n_1658),
.A2(n_1642),
.B1(n_1640),
.B2(n_1622),
.C(n_1620),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1653),
.A2(n_1622),
.B(n_1601),
.Y(n_1681)
);

AOI22x1_ASAP7_75t_L g1682 ( 
.A1(n_1653),
.A2(n_1230),
.B1(n_1620),
.B2(n_1618),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1656),
.B(n_1597),
.Y(n_1683)
);

NAND3xp33_ASAP7_75t_SL g1684 ( 
.A(n_1673),
.B(n_1582),
.C(n_1601),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1654),
.Y(n_1685)
);

NOR3x1_ASAP7_75t_L g1686 ( 
.A(n_1678),
.B(n_1664),
.C(n_1666),
.Y(n_1686)
);

NAND5xp2_ASAP7_75t_L g1687 ( 
.A(n_1674),
.B(n_1672),
.C(n_1667),
.D(n_1655),
.E(n_1669),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1685),
.Y(n_1688)
);

NOR2x1_ASAP7_75t_L g1689 ( 
.A(n_1676),
.B(n_1658),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1679),
.A2(n_1672),
.B1(n_1659),
.B2(n_1669),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1683),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1677),
.B(n_1660),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1675),
.B(n_1660),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_SL g1694 ( 
.A(n_1682),
.B(n_1670),
.Y(n_1694)
);

NOR3xp33_ASAP7_75t_L g1695 ( 
.A(n_1684),
.B(n_1661),
.C(n_1657),
.Y(n_1695)
);

OAI21xp33_ASAP7_75t_L g1696 ( 
.A1(n_1681),
.A2(n_1670),
.B(n_1661),
.Y(n_1696)
);

NOR2x1_ASAP7_75t_L g1697 ( 
.A(n_1689),
.B(n_1663),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1687),
.A2(n_1665),
.B1(n_1663),
.B2(n_1680),
.C(n_1603),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1690),
.B(n_1603),
.Y(n_1699)
);

NOR2xp67_ASAP7_75t_L g1700 ( 
.A(n_1688),
.B(n_1604),
.Y(n_1700)
);

OAI21xp33_ASAP7_75t_L g1701 ( 
.A1(n_1692),
.A2(n_1618),
.B(n_1612),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1693),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1697),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1700),
.B(n_1696),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1702),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1698),
.A2(n_1695),
.B1(n_1694),
.B2(n_1691),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1699),
.B(n_1686),
.Y(n_1707)
);

AND2x2_ASAP7_75t_SL g1708 ( 
.A(n_1701),
.B(n_1224),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_1702),
.Y(n_1709)
);

OAI211xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1706),
.A2(n_1617),
.B(n_1613),
.C(n_1612),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1703),
.Y(n_1711)
);

NOR3xp33_ASAP7_75t_L g1712 ( 
.A(n_1707),
.B(n_1330),
.C(n_1604),
.Y(n_1712)
);

OAI321xp33_ASAP7_75t_L g1713 ( 
.A1(n_1705),
.A2(n_1704),
.A3(n_1709),
.B1(n_1708),
.B2(n_1613),
.C(n_1617),
.Y(n_1713)
);

NAND3xp33_ASAP7_75t_L g1714 ( 
.A(n_1704),
.B(n_1534),
.C(n_1532),
.Y(n_1714)
);

NOR3xp33_ASAP7_75t_L g1715 ( 
.A(n_1707),
.B(n_1370),
.C(n_1329),
.Y(n_1715)
);

OAI22x1_ASAP7_75t_L g1716 ( 
.A1(n_1711),
.A2(n_1542),
.B1(n_1576),
.B2(n_1574),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1714),
.B(n_1584),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1713),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1712),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1717),
.Y(n_1720)
);

XOR2xp5_ASAP7_75t_L g1721 ( 
.A(n_1718),
.B(n_1715),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1710),
.B1(n_1719),
.B2(n_1716),
.Y(n_1722)
);

OAI22x1_ASAP7_75t_L g1723 ( 
.A1(n_1722),
.A2(n_1720),
.B1(n_1574),
.B2(n_1576),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1722),
.Y(n_1724)
);

OAI22xp33_ASAP7_75t_SL g1725 ( 
.A1(n_1724),
.A2(n_1579),
.B1(n_1555),
.B2(n_1549),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1723),
.A2(n_1383),
.B1(n_1339),
.B2(n_1531),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1725),
.A2(n_1548),
.B(n_1571),
.Y(n_1727)
);

AOI222xp33_ASAP7_75t_L g1728 ( 
.A1(n_1727),
.A2(n_1726),
.B1(n_1383),
.B2(n_1339),
.C1(n_1360),
.C2(n_1521),
.Y(n_1728)
);

AOI222xp33_ASAP7_75t_L g1729 ( 
.A1(n_1728),
.A2(n_1339),
.B1(n_1383),
.B2(n_1360),
.C1(n_1531),
.C2(n_1521),
.Y(n_1729)
);

AOI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1729),
.A2(n_1511),
.B1(n_1508),
.B2(n_1529),
.C(n_1531),
.Y(n_1730)
);

AOI211xp5_ASAP7_75t_L g1731 ( 
.A1(n_1730),
.A2(n_1521),
.B(n_1529),
.C(n_1511),
.Y(n_1731)
);


endmodule