module real_jpeg_5695_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_0),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_0),
.Y(n_132)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_0),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_1),
.A2(n_26),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_1),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_1),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_1),
.A2(n_40),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_1),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_1),
.A2(n_153),
.B1(n_216),
.B2(n_219),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_1),
.A2(n_255),
.B(n_258),
.C(n_261),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_1),
.B(n_269),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_1),
.B(n_59),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_1),
.B(n_79),
.C(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_1),
.B(n_116),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_1),
.B(n_112),
.C(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_1),
.B(n_33),
.Y(n_329)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_3),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_3),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_3),
.A2(n_87),
.B1(n_118),
.B2(n_122),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_3),
.A2(n_30),
.B1(n_87),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_3),
.A2(n_87),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_4),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_4),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_4),
.A2(n_93),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_4),
.A2(n_93),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_4),
.A2(n_93),
.B1(n_196),
.B2(n_200),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_6),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_7),
.Y(n_168)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_7),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_7),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_7),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_8),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_14)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_9),
.Y(n_257)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_12),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_12),
.A2(n_28),
.B1(n_145),
.B2(n_148),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_12),
.A2(n_28),
.B1(n_185),
.B2(n_189),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_12),
.A2(n_28),
.B1(n_166),
.B2(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_13),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_13),
.Y(n_81)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_405),
.B(n_407),
.Y(n_19)
);

AO21x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_133),
.B(n_404),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_130),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_22),
.B(n_130),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_124),
.C(n_128),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_23),
.B(n_401),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_56),
.C(n_88),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_24),
.A2(n_179),
.B1(n_180),
.B2(n_191),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_24),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_24),
.B(n_140),
.C(n_180),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_24),
.B(n_236),
.C(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_24),
.A2(n_191),
.B1(n_236),
.B2(n_330),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_24),
.A2(n_191),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B1(n_52),
.B2(n_55),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_25),
.A2(n_32),
.B1(n_52),
.B2(n_55),
.Y(n_224)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_32),
.A2(n_52),
.B1(n_55),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_32),
.A2(n_55),
.B1(n_125),
.B2(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_32),
.A2(n_52),
.B(n_55),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g406 ( 
.A1(n_32),
.A2(n_55),
.B(n_131),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_42),
.Y(n_32)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_34),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_35),
.Y(n_183)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_36),
.Y(n_121)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_40),
.Y(n_260)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_56),
.A2(n_88),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_56),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_56),
.B(n_224),
.C(n_381),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_56),
.A2(n_379),
.B1(n_381),
.B2(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_84),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_57),
.B(n_150),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_72),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_58),
.A2(n_72),
.B1(n_143),
.B2(n_149),
.Y(n_142)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_59),
.A2(n_195),
.B(n_201),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_59),
.B(n_144),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_59),
.A2(n_73),
.B1(n_84),
.B2(n_195),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_70),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_64),
.Y(n_167)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g162 ( 
.A(n_65),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g218 ( 
.A(n_65),
.Y(n_218)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_69),
.Y(n_174)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_73),
.B(n_150),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_80),
.B2(n_82),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_76),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_76),
.Y(n_293)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_86),
.Y(n_200)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_88),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_95),
.B1(n_116),
.B2(n_117),
.Y(n_88)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_89),
.Y(n_382)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_92),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_95),
.B(n_223),
.Y(n_383)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_96),
.B(n_107),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_96),
.A2(n_107),
.B1(n_181),
.B2(n_184),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g236 ( 
.A1(n_96),
.A2(n_107),
.B1(n_181),
.B2(n_184),
.Y(n_236)
);

NAND2x1_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_107),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B1(n_104),
.B2(n_106),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_103),
.Y(n_312)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_107),
.A2(n_382),
.B(n_383),
.Y(n_381)
);

AOI22x1_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_114),
.Y(n_107)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx8_ASAP7_75t_L g314 ( 
.A(n_110),
.Y(n_314)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_124),
.B(n_128),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_129),
.B(n_223),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_130),
.B(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_130),
.B(n_406),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_399),
.B(n_403),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_370),
.B(n_396),
.Y(n_134)
);

OAI211xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_270),
.B(n_364),
.C(n_369),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_241),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g364 ( 
.A1(n_137),
.A2(n_241),
.B(n_365),
.C(n_368),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_225),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_138),
.B(n_225),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_192),
.C(n_208),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_139),
.B(n_192),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_178),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_158),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_141),
.A2(n_142),
.B1(n_158),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_141),
.A2(n_142),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_141),
.A2(n_142),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_142),
.B(n_265),
.C(n_302),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_142),
.B(n_322),
.C(n_324),
.Y(n_335)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_158),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_164),
.B1(n_169),
.B2(n_175),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_160),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_164),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_165),
.A2(n_215),
.B1(n_266),
.B2(n_269),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_165),
.A2(n_215),
.B1(n_266),
.B2(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_166),
.Y(n_281)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_172),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_172),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_179),
.A2(n_180),
.B1(n_220),
.B2(n_291),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_179),
.B(n_291),
.C(n_309),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_179),
.A2(n_180),
.B1(n_340),
.B2(n_341),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_180),
.B(n_224),
.C(n_340),
.Y(n_357)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_182),
.A2(n_256),
.B(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_203),
.B2(n_207),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_203),
.Y(n_232)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_207),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_203),
.A2(n_231),
.B(n_232),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_204),
.B(n_215),
.Y(n_315)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_222),
.C(n_224),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_220),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_211),
.A2(n_220),
.B1(n_291),
.B2(n_356),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_211),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_220),
.A2(n_291),
.B1(n_292),
.B2(n_296),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_220),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_222),
.A2(n_224),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_224),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_224),
.A2(n_248),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_224),
.A2(n_248),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_224),
.A2(n_248),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_224),
.B(n_375),
.C(n_380),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_239),
.B2(n_240),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_233),
.B1(n_234),
.B2(n_238),
.Y(n_227)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_233),
.B(n_238),
.C(n_240),
.Y(n_395)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B(n_237),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_236),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_236),
.A2(n_326),
.B1(n_327),
.B2(n_330),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_236),
.Y(n_330)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_237),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_237),
.A2(n_385),
.B1(n_389),
.B2(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_239),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_242),
.B(n_244),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_250),
.C(n_252),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_246),
.B(n_250),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_252),
.B(n_363),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_253),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_264),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_254),
.A2(n_264),
.B1(n_265),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_254),
.Y(n_347)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_264),
.A2(n_265),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_265),
.B(n_286),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_286),
.Y(n_287)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_349),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_334),
.B(n_348),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_319),
.B(n_333),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_306),
.B(n_318),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_298),
.B(n_305),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_288),
.B(n_297),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_285),
.B(n_287),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_283),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_283),
.A2(n_289),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_290),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_289),
.B(n_328),
.C(n_330),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_296),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_292),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_304),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_304),
.Y(n_305)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_308),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_317),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_315),
.B2(n_316),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_316),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_332),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_332),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_324),
.B1(n_325),
.B2(n_331),
.Y(n_320)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_321),
.Y(n_331)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_336),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_342),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_344),
.C(n_345),
.Y(n_358)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_345),
.B2(n_346),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NOR2x1_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_359),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_358),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_358),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_354),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_352),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_355),
.B(n_357),
.C(n_361),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_359),
.A2(n_366),
.B(n_367),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_360),
.B(n_362),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_391),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_371),
.A2(n_397),
.B(n_398),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_384),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_384),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_380),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_381),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_389),
.C(n_390),
.Y(n_384)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_385),
.Y(n_394)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_390),
.B(n_393),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_395),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_395),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_400),
.B(n_402),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_408),
.Y(n_407)
);


endmodule