module fake_jpeg_21363_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_40),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_0),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_16),
.B1(n_26),
.B2(n_22),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_48),
.B1(n_49),
.B2(n_24),
.Y(n_58)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_27),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_26),
.B1(n_22),
.B2(n_30),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_26),
.B1(n_24),
.B2(n_30),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_19),
.C(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_18),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_64),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_67),
.Y(n_92)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_62),
.A2(n_74),
.B1(n_85),
.B2(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_71),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_38),
.C(n_36),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_21),
.C(n_31),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_80),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_39),
.B1(n_41),
.B2(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_51),
.A2(n_25),
.B1(n_28),
.B2(n_17),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_31),
.CI(n_27),
.CON(n_93),
.SN(n_93)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_19),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_79),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_54),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_36),
.Y(n_99)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_18),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_84),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_38),
.B(n_36),
.C(n_27),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_62),
.B1(n_74),
.B2(n_73),
.Y(n_119)
);

BUFx24_ASAP7_75t_SL g115 ( 
.A(n_93),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_81),
.B1(n_64),
.B2(n_60),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_75),
.B1(n_66),
.B2(n_61),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_38),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_105),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_63),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_32),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_109),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_111),
.B(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_78),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_85),
.B(n_72),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_114),
.B(n_126),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_71),
.B(n_58),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_60),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_107),
.B(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_93),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_91),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_120),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_134),
.B1(n_87),
.B2(n_88),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_91),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_127),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_119),
.B(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_69),
.B(n_80),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_70),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_130),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_84),
.B(n_32),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_109),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_132),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_87),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_133),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_89),
.A2(n_92),
.B1(n_101),
.B2(n_105),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_148),
.B1(n_151),
.B2(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_104),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_115),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_152),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_110),
.B1(n_93),
.B2(n_102),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_113),
.B(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_90),
.A3(n_88),
.B1(n_94),
.B2(n_103),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_127),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_70),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_156),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_165),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_152),
.B1(n_137),
.B2(n_146),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_124),
.C(n_134),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_166),
.C(n_170),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_171),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_124),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_90),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_173),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_118),
.C(n_120),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_86),
.A3(n_94),
.B1(n_103),
.B2(n_21),
.C1(n_108),
.C2(n_11),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_143),
.Y(n_172)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_108),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_168),
.A2(n_151),
.B1(n_150),
.B2(n_149),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_190),
.B1(n_160),
.B2(n_173),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_142),
.C(n_138),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_183),
.C(n_139),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_155),
.C(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_188),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_170),
.C(n_165),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_194),
.C(n_201),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_193),
.A2(n_177),
.B1(n_187),
.B2(n_189),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_166),
.C(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_145),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_176),
.B1(n_169),
.B2(n_159),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_189),
.B1(n_185),
.B2(n_75),
.Y(n_208)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_135),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_182),
.C(n_183),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_4),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_209),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_191),
.B1(n_200),
.B2(n_192),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_14),
.C(n_13),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_0),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_206),
.A2(n_12),
.B(n_11),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_210),
.B(n_204),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_213),
.A2(n_216),
.B1(n_5),
.B2(n_6),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_207),
.B(n_1),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_4),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_1),
.C(n_2),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_217),
.C(n_203),
.Y(n_221)
);

NOR2x1_ASAP7_75t_SL g218 ( 
.A(n_212),
.B(n_202),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_214),
.B(n_6),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_221),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_222),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_224),
.B(n_5),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_219),
.B(n_7),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_226),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_227),
.B(n_225),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_5),
.B(n_7),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g231 ( 
.A(n_230),
.Y(n_231)
);


endmodule