module fake_jpeg_11670_n_28 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_28);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_28;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

INVx1_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_13),
.A2(n_5),
.B(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_16),
.B(n_17),
.Y(n_18)
);

INVx4_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_13),
.C(n_11),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_22),
.B(n_23),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_0),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_0),
.B(n_1),
.Y(n_26)
);

AOI21x1_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_25),
.B(n_2),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_10),
.Y(n_28)
);


endmodule