module fake_netlist_1_1634_n_1340 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1340);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1340;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_533;
wire n_1010;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_409;
wire n_315;
wire n_295;
wire n_1321;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_274;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g273 ( .A(n_108), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_150), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_269), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_231), .Y(n_276) );
INVxp33_ASAP7_75t_SL g277 ( .A(n_201), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_155), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_235), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_258), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_244), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_104), .Y(n_282) );
INVxp67_ASAP7_75t_L g283 ( .A(n_238), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_62), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_188), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_211), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_0), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_142), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_194), .Y(n_289) );
BUFx10_ASAP7_75t_L g290 ( .A(n_245), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_189), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_185), .Y(n_292) );
INVxp33_ASAP7_75t_L g293 ( .A(n_39), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_152), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_66), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_15), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_271), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_105), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_197), .B(n_239), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_166), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_100), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_246), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_263), .Y(n_303) );
CKINVDCx14_ASAP7_75t_R g304 ( .A(n_186), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_41), .Y(n_305) );
INVxp67_ASAP7_75t_L g306 ( .A(n_190), .Y(n_306) );
INVxp67_ASAP7_75t_L g307 ( .A(n_253), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_202), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_124), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_14), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_157), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_38), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_179), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_3), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_181), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_34), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_130), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_174), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_101), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_153), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_134), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_135), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_36), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_184), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_233), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_267), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_270), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_206), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_214), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_170), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_131), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_224), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_87), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_195), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_159), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_12), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_137), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_175), .Y(n_338) );
BUFx5_ASAP7_75t_L g339 ( .A(n_127), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_151), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_193), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_59), .Y(n_342) );
CKINVDCx16_ASAP7_75t_R g343 ( .A(n_232), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_243), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_154), .Y(n_345) );
BUFx10_ASAP7_75t_L g346 ( .A(n_133), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_173), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_119), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_2), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_16), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_145), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_234), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_112), .Y(n_353) );
BUFx2_ASAP7_75t_L g354 ( .A(n_257), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_167), .Y(n_355) );
CKINVDCx16_ASAP7_75t_R g356 ( .A(n_209), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_259), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_143), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_165), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_180), .Y(n_360) );
INVxp67_ASAP7_75t_SL g361 ( .A(n_204), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_96), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_178), .Y(n_363) );
NOR2xp67_ASAP7_75t_L g364 ( .A(n_268), .B(n_121), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_53), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_223), .Y(n_366) );
INVxp33_ASAP7_75t_SL g367 ( .A(n_25), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_1), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_45), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_68), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_203), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_6), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_63), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_67), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_112), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_73), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_78), .Y(n_377) );
INVxp33_ASAP7_75t_L g378 ( .A(n_163), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_164), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_146), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_261), .Y(n_381) );
NOR2xp67_ASAP7_75t_L g382 ( .A(n_215), .B(n_38), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_50), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_111), .Y(n_384) );
CKINVDCx14_ASAP7_75t_R g385 ( .A(n_9), .Y(n_385) );
CKINVDCx16_ASAP7_75t_R g386 ( .A(n_6), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_17), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_191), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_248), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_125), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_252), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_225), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_76), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_200), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_94), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_221), .Y(n_396) );
CKINVDCx14_ASAP7_75t_R g397 ( .A(n_132), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_260), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_168), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_105), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_82), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_255), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g403 ( .A(n_41), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_104), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_78), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_65), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_36), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_210), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_230), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_241), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_207), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_2), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_40), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_218), .Y(n_414) );
BUFx2_ASAP7_75t_SL g415 ( .A(n_266), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_48), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_24), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_187), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_80), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_222), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_192), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_264), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_242), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_103), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_183), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_250), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_25), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_229), .Y(n_428) );
INVxp33_ASAP7_75t_SL g429 ( .A(n_75), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_34), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_240), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_156), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_19), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_247), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_205), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_392), .Y(n_436) );
INVx4_ASAP7_75t_L g437 ( .A(n_392), .Y(n_437) );
INVx4_ASAP7_75t_L g438 ( .A(n_392), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_339), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_305), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_305), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_349), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_349), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_280), .B(n_1), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_339), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_275), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_278), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_339), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_332), .B(n_3), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_339), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_279), .Y(n_451) );
NAND2xp33_ASAP7_75t_R g452 ( .A(n_277), .B(n_126), .Y(n_452) );
AND2x6_ASAP7_75t_L g453 ( .A(n_325), .B(n_128), .Y(n_453) );
OAI22x1_ASAP7_75t_SL g454 ( .A1(n_353), .A2(n_7), .B1(n_4), .B2(n_5), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_290), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_290), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_281), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_339), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_354), .B(n_4), .Y(n_459) );
OAI22xp5_ASAP7_75t_SL g460 ( .A1(n_353), .A2(n_8), .B1(n_5), .B2(n_7), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_285), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_293), .B(n_8), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_288), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_297), .Y(n_464) );
AND2x6_ASAP7_75t_L g465 ( .A(n_325), .B(n_129), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_385), .A2(n_429), .B1(n_367), .B2(n_403), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_339), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_300), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_339), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_340), .Y(n_470) );
INVx3_ASAP7_75t_L g471 ( .A(n_290), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_340), .Y(n_472) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_340), .Y(n_473) );
CKINVDCx8_ASAP7_75t_R g474 ( .A(n_343), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_302), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_385), .Y(n_476) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_340), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_409), .B(n_9), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_436), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_462), .A2(n_293), .B1(n_282), .B2(n_284), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_476), .B(n_378), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_455), .B(n_356), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_455), .B(n_320), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_436), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_436), .B(n_344), .Y(n_485) );
BUFx3_ASAP7_75t_L g486 ( .A(n_453), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_455), .B(n_346), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_437), .Y(n_489) );
INVxp67_ASAP7_75t_SL g490 ( .A(n_462), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_439), .Y(n_491) );
BUFx10_ASAP7_75t_L g492 ( .A(n_476), .Y(n_492) );
BUFx4f_ASAP7_75t_L g493 ( .A(n_453), .Y(n_493) );
NOR2x1p5_ASAP7_75t_L g494 ( .A(n_455), .B(n_298), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_437), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_462), .A2(n_287), .B1(n_295), .B2(n_273), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_439), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_456), .B(n_378), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_445), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_445), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_456), .B(n_346), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_466), .A2(n_370), .B1(n_404), .B2(n_386), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_437), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_473), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_437), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_456), .B(n_351), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_456), .B(n_304), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_471), .B(n_304), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_438), .B(n_276), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_466), .A2(n_429), .B1(n_367), .B2(n_352), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_438), .B(n_276), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_445), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_471), .B(n_283), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_471), .B(n_306), .Y(n_514) );
INVx4_ASAP7_75t_L g515 ( .A(n_438), .Y(n_515) );
INVx8_ASAP7_75t_L g516 ( .A(n_453), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_438), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_446), .B(n_291), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_474), .A2(n_404), .B1(n_370), .B2(n_352), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_471), .B(n_307), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_478), .A2(n_296), .B1(n_310), .B2(n_309), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_446), .B(n_291), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_448), .Y(n_523) );
OR2x6_ASAP7_75t_L g524 ( .A(n_460), .B(n_415), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_490), .A2(n_478), .B1(n_444), .B2(n_459), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_490), .B(n_478), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_485), .B(n_478), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_516), .Y(n_528) );
BUFx12f_ASAP7_75t_L g529 ( .A(n_492), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_485), .B(n_449), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_507), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_498), .B(n_447), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_488), .B(n_501), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_507), .Y(n_534) );
INVxp67_ASAP7_75t_L g535 ( .A(n_481), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_483), .B(n_447), .Y(n_536) );
NOR2x1p5_ASAP7_75t_L g537 ( .A(n_481), .B(n_298), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_483), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_483), .B(n_451), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_483), .B(n_451), .Y(n_540) );
OAI221xp5_ASAP7_75t_L g541 ( .A1(n_480), .A2(n_474), .B1(n_461), .B2(n_464), .C(n_463), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_518), .A2(n_457), .B1(n_463), .B2(n_461), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_506), .B(n_457), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_506), .B(n_464), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_506), .B(n_468), .Y(n_545) );
NOR2xp67_ASAP7_75t_L g546 ( .A(n_510), .B(n_442), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_506), .Y(n_547) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_516), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_489), .Y(n_549) );
NOR2xp67_ASAP7_75t_L g550 ( .A(n_510), .B(n_442), .Y(n_550) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_516), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_494), .A2(n_496), .B1(n_508), .B2(n_521), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_492), .Y(n_553) );
OAI22xp5_ASAP7_75t_SL g554 ( .A1(n_524), .A2(n_460), .B1(n_358), .B2(n_396), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_493), .B(n_448), .Y(n_555) );
NOR2x1p5_ASAP7_75t_L g556 ( .A(n_502), .B(n_301), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_508), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_513), .B(n_468), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_514), .B(n_475), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_520), .B(n_475), .Y(n_560) );
NOR2xp67_ASAP7_75t_L g561 ( .A(n_502), .B(n_443), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_515), .B(n_474), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_489), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_519), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_515), .B(n_443), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_493), .B(n_448), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_509), .Y(n_567) );
CKINVDCx11_ASAP7_75t_R g568 ( .A(n_524), .Y(n_568) );
BUFx3_ASAP7_75t_L g569 ( .A(n_516), .Y(n_569) );
INVx3_ASAP7_75t_L g570 ( .A(n_489), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_492), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_482), .B(n_277), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_509), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_511), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_489), .B(n_294), .Y(n_575) );
INVx2_ASAP7_75t_SL g576 ( .A(n_492), .Y(n_576) );
AO22x1_ASAP7_75t_L g577 ( .A1(n_519), .A2(n_362), .B1(n_372), .B2(n_301), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_517), .B(n_440), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_495), .Y(n_579) );
AND2x6_ASAP7_75t_SL g580 ( .A(n_524), .B(n_454), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_517), .B(n_440), .Y(n_581) );
AOI21x1_ASAP7_75t_L g582 ( .A1(n_511), .A2(n_458), .B(n_450), .Y(n_582) );
NAND2x1p5_ASAP7_75t_L g583 ( .A(n_494), .B(n_312), .Y(n_583) );
NOR2xp67_ASAP7_75t_L g584 ( .A(n_522), .B(n_441), .Y(n_584) );
BUFx12f_ASAP7_75t_L g585 ( .A(n_524), .Y(n_585) );
INVx4_ASAP7_75t_L g586 ( .A(n_516), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_522), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_493), .B(n_450), .Y(n_588) );
INVx5_ASAP7_75t_L g589 ( .A(n_516), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_503), .B(n_321), .Y(n_590) );
INVx3_ASAP7_75t_L g591 ( .A(n_503), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_503), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_505), .Y(n_593) );
NOR3x1_ASAP7_75t_L g594 ( .A(n_524), .B(n_454), .C(n_424), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_505), .B(n_321), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_505), .Y(n_596) );
NAND2xp33_ASAP7_75t_L g597 ( .A(n_517), .B(n_453), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_479), .B(n_324), .Y(n_598) );
NOR2x1p5_ASAP7_75t_L g599 ( .A(n_524), .B(n_362), .Y(n_599) );
BUFx3_ASAP7_75t_L g600 ( .A(n_486), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_484), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_484), .B(n_324), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_487), .B(n_360), .Y(n_603) );
INVx3_ASAP7_75t_L g604 ( .A(n_491), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_497), .A2(n_358), .B1(n_396), .B2(n_311), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_497), .B(n_441), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_499), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_500), .A2(n_465), .B1(n_453), .B2(n_467), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_535), .B(n_311), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_564), .A2(n_383), .B(n_407), .C(n_336), .Y(n_610) );
NOR2xp67_ASAP7_75t_SL g611 ( .A(n_529), .B(n_372), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_576), .B(n_553), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_571), .B(n_371), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_530), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_587), .B(n_371), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_536), .B(n_512), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_538), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_555), .A2(n_523), .B(n_512), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_539), .B(n_523), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_538), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_540), .B(n_405), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_547), .Y(n_622) );
O2A1O1Ixp33_ASAP7_75t_L g623 ( .A1(n_541), .A2(n_412), .B(n_433), .C(n_387), .Y(n_623) );
INVx3_ASAP7_75t_L g624 ( .A(n_604), .Y(n_624) );
BUFx12f_ASAP7_75t_L g625 ( .A(n_568), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_547), .B(n_398), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_543), .B(n_405), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_537), .A2(n_546), .B1(n_550), .B2(n_552), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_572), .B(n_398), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_526), .A2(n_333), .B(n_342), .C(n_314), .Y(n_630) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_544), .A2(n_350), .B(n_365), .C(n_348), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_555), .A2(n_469), .B(n_299), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_584), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_567), .A2(n_425), .B1(n_397), .B2(n_381), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_573), .A2(n_425), .B1(n_397), .B2(n_381), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_566), .A2(n_361), .B(n_504), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_570), .Y(n_637) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_545), .A2(n_373), .B(n_374), .C(n_368), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_561), .A2(n_452), .B1(n_316), .B2(n_319), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_574), .A2(n_525), .B1(n_527), .B2(n_542), .Y(n_640) );
A2O1A1Ixp33_ASAP7_75t_L g641 ( .A1(n_578), .A2(n_376), .B(n_390), .C(n_384), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_570), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g643 ( .A(n_605), .B(n_377), .C(n_369), .Y(n_643) );
NOR2xp33_ASAP7_75t_R g644 ( .A(n_585), .B(n_380), .Y(n_644) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_528), .Y(n_645) );
BUFx3_ASAP7_75t_L g646 ( .A(n_583), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_583), .B(n_323), .Y(n_647) );
INVx4_ASAP7_75t_L g648 ( .A(n_589), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_582), .A2(n_465), .B(n_453), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_542), .A2(n_395), .B1(n_400), .B2(n_393), .Y(n_650) );
OAI22x1_ASAP7_75t_L g651 ( .A1(n_556), .A2(n_413), .B1(n_402), .B2(n_380), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g652 ( .A1(n_578), .A2(n_406), .B(n_416), .C(n_401), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_532), .A2(n_419), .B1(n_427), .B2(n_417), .Y(n_653) );
CKINVDCx11_ASAP7_75t_R g654 ( .A(n_580), .Y(n_654) );
AND3x1_ASAP7_75t_SL g655 ( .A(n_599), .B(n_430), .C(n_315), .Y(n_655) );
A2O1A1Ixp33_ASAP7_75t_L g656 ( .A1(n_581), .A2(n_382), .B(n_364), .C(n_317), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_591), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_533), .B(n_418), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_591), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_593), .Y(n_660) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_528), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_577), .Y(n_662) );
O2A1O1Ixp33_ASAP7_75t_L g663 ( .A1(n_531), .A2(n_326), .B(n_327), .C(n_322), .Y(n_663) );
CKINVDCx8_ASAP7_75t_R g664 ( .A(n_594), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_534), .A2(n_557), .B1(n_559), .B2(n_558), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_569), .B(n_328), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_560), .A2(n_330), .B(n_331), .C(n_329), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_606), .A2(n_337), .B1(n_338), .B2(n_335), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_606), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_607), .B(n_346), .Y(n_670) );
INVxp67_ASAP7_75t_L g671 ( .A(n_605), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_565), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_603), .B(n_375), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_533), .B(n_274), .Y(n_674) );
INVx4_ASAP7_75t_L g675 ( .A(n_589), .Y(n_675) );
INVx3_ASAP7_75t_L g676 ( .A(n_586), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_554), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_598), .B(n_375), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_602), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_588), .A2(n_596), .B(n_592), .Y(n_680) );
BUFx2_ASAP7_75t_L g681 ( .A(n_575), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_601), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_562), .A2(n_359), .B(n_363), .C(n_357), .Y(n_683) );
NOR2xp33_ASAP7_75t_R g684 ( .A(n_597), .B(n_318), .Y(n_684) );
NOR2xp33_ASAP7_75t_R g685 ( .A(n_569), .B(n_334), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_563), .Y(n_686) );
CKINVDCx5p33_ASAP7_75t_R g687 ( .A(n_590), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g688 ( .A1(n_595), .A2(n_420), .B1(n_426), .B2(n_411), .Y(n_688) );
BUFx12f_ASAP7_75t_L g689 ( .A(n_528), .Y(n_689) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_549), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_579), .Y(n_691) );
NOR3xp33_ASAP7_75t_SL g692 ( .A(n_608), .B(n_434), .C(n_428), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_600), .B(n_286), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_608), .A2(n_389), .B1(n_391), .B2(n_388), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_528), .B(n_289), .Y(n_695) );
NAND2x1p5_ASAP7_75t_L g696 ( .A(n_548), .B(n_347), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g697 ( .A(n_548), .B(n_313), .C(n_308), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_548), .A2(n_399), .B(n_394), .Y(n_698) );
O2A1O1Ixp5_ASAP7_75t_L g699 ( .A1(n_548), .A2(n_303), .B(n_341), .C(n_292), .Y(n_699) );
BUFx2_ASAP7_75t_L g700 ( .A(n_551), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_551), .A2(n_423), .B(n_408), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_551), .A2(n_432), .B1(n_379), .B2(n_414), .Y(n_702) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_578), .A2(n_303), .B(n_341), .C(n_292), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_535), .B(n_10), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_535), .B(n_10), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_587), .B(n_345), .Y(n_706) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_553), .B(n_431), .Y(n_707) );
AO31x2_ASAP7_75t_L g708 ( .A1(n_606), .A2(n_410), .A3(n_435), .B(n_422), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_587), .Y(n_709) );
BUFx12f_ASAP7_75t_L g710 ( .A(n_568), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_526), .A2(n_410), .B1(n_435), .B2(n_422), .Y(n_711) );
INVx5_ASAP7_75t_L g712 ( .A(n_529), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_535), .B(n_11), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_553), .B(n_421), .Y(n_714) );
BUFx3_ASAP7_75t_L g715 ( .A(n_529), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_587), .A2(n_472), .B1(n_470), .B2(n_366), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_587), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_604), .Y(n_718) );
OAI22x1_ASAP7_75t_L g719 ( .A1(n_556), .A2(n_13), .B1(n_11), .B2(n_12), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g720 ( .A1(n_578), .A2(n_472), .B(n_470), .C(n_366), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_553), .B(n_355), .Y(n_721) );
O2A1O1Ixp33_ASAP7_75t_L g722 ( .A1(n_535), .A2(n_15), .B(n_13), .C(n_14), .Y(n_722) );
INVx1_ASAP7_75t_SL g723 ( .A(n_553), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_587), .B(n_465), .Y(n_724) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_529), .Y(n_725) );
BUFx2_ASAP7_75t_L g726 ( .A(n_529), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g727 ( .A1(n_567), .A2(n_465), .B(n_473), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_605), .B(n_17), .Y(n_728) );
AND2x4_ASAP7_75t_L g729 ( .A(n_576), .B(n_465), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_587), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_614), .Y(n_731) );
CKINVDCx16_ASAP7_75t_R g732 ( .A(n_715), .Y(n_732) );
CKINVDCx6p67_ASAP7_75t_R g733 ( .A(n_712), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_665), .B(n_18), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_610), .A2(n_477), .B1(n_19), .B2(n_20), .C(n_21), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_709), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_682), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_686), .Y(n_738) );
AO31x2_ASAP7_75t_L g739 ( .A1(n_703), .A2(n_477), .A3(n_21), .B(n_18), .Y(n_739) );
BUFx3_ASAP7_75t_L g740 ( .A(n_712), .Y(n_740) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_665), .A2(n_671), .B1(n_653), .B2(n_643), .C(n_623), .Y(n_741) );
AO31x2_ASAP7_75t_L g742 ( .A1(n_656), .A2(n_477), .A3(n_23), .B(n_20), .Y(n_742) );
OAI22xp33_ASAP7_75t_L g743 ( .A1(n_728), .A2(n_24), .B1(n_22), .B2(n_23), .Y(n_743) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_712), .A2(n_27), .B1(n_22), .B2(n_26), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_609), .B(n_26), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_626), .B(n_27), .Y(n_746) );
BUFx12f_ASAP7_75t_L g747 ( .A(n_712), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_640), .A2(n_477), .B1(n_30), .B2(n_28), .Y(n_748) );
OAI22x1_ASAP7_75t_L g749 ( .A1(n_662), .A2(n_30), .B1(n_28), .B2(n_29), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_629), .B(n_29), .Y(n_750) );
AO21x1_ASAP7_75t_L g751 ( .A1(n_694), .A2(n_138), .B(n_136), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_723), .Y(n_752) );
INVxp67_ASAP7_75t_L g753 ( .A(n_723), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g754 ( .A(n_625), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_632), .A2(n_140), .B(n_139), .Y(n_755) );
INVx3_ASAP7_75t_L g756 ( .A(n_689), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_717), .B(n_31), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_730), .Y(n_758) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_645), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_620), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_628), .B(n_32), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_669), .B(n_32), .Y(n_762) );
OR2x2_ASAP7_75t_L g763 ( .A(n_726), .B(n_33), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_617), .B(n_33), .Y(n_764) );
NOR2x1_ASAP7_75t_L g765 ( .A(n_648), .B(n_35), .Y(n_765) );
O2A1O1Ixp33_ASAP7_75t_L g766 ( .A1(n_641), .A2(n_39), .B(n_35), .C(n_37), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_691), .Y(n_767) );
OAI21xp5_ASAP7_75t_L g768 ( .A1(n_618), .A2(n_144), .B(n_141), .Y(n_768) );
INVx3_ASAP7_75t_L g769 ( .A(n_675), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_704), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_677), .A2(n_42), .B1(n_37), .B2(n_40), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g772 ( .A(n_710), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_662), .A2(n_42), .B1(n_43), .B2(n_44), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_705), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_678), .Y(n_775) );
AO31x2_ASAP7_75t_L g776 ( .A1(n_711), .A2(n_43), .A3(n_44), .B(n_45), .Y(n_776) );
NAND2xp33_ASAP7_75t_L g777 ( .A(n_684), .B(n_147), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_649), .A2(n_149), .B(n_148), .Y(n_778) );
A2O1A1Ixp33_ASAP7_75t_L g779 ( .A1(n_683), .A2(n_46), .B(n_47), .C(n_48), .Y(n_779) );
INVx1_ASAP7_75t_SL g780 ( .A(n_646), .Y(n_780) );
A2O1A1Ixp33_ASAP7_75t_L g781 ( .A1(n_667), .A2(n_46), .B(n_47), .C(n_49), .Y(n_781) );
OR2x2_ASAP7_75t_L g782 ( .A(n_634), .B(n_49), .Y(n_782) );
NOR2xp33_ASAP7_75t_SL g783 ( .A(n_725), .B(n_50), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_673), .Y(n_784) );
AOI221xp5_ASAP7_75t_SL g785 ( .A1(n_630), .A2(n_51), .B1(n_52), .B2(n_53), .C(n_54), .Y(n_785) );
A2O1A1Ixp33_ASAP7_75t_L g786 ( .A1(n_631), .A2(n_51), .B(n_52), .C(n_54), .Y(n_786) );
INVx4_ASAP7_75t_L g787 ( .A(n_612), .Y(n_787) );
AO31x2_ASAP7_75t_L g788 ( .A1(n_711), .A2(n_55), .A3(n_56), .B(n_57), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_696), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_652), .B(n_55), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_690), .Y(n_791) );
BUFx2_ASAP7_75t_L g792 ( .A(n_612), .Y(n_792) );
AO31x2_ASAP7_75t_L g793 ( .A1(n_720), .A2(n_56), .A3(n_57), .B(n_58), .Y(n_793) );
OAI22xp33_ASAP7_75t_L g794 ( .A1(n_635), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_794) );
BUFx2_ASAP7_75t_L g795 ( .A(n_685), .Y(n_795) );
INVx3_ASAP7_75t_L g796 ( .A(n_675), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_616), .A2(n_619), .B1(n_672), .B2(n_622), .Y(n_797) );
BUFx3_ASAP7_75t_L g798 ( .A(n_654), .Y(n_798) );
O2A1O1Ixp5_ASAP7_75t_SL g799 ( .A1(n_714), .A2(n_171), .B(n_265), .C(n_262), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_713), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_650), .A2(n_61), .B1(n_63), .B2(n_64), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_650), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_696), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g804 ( .A1(n_680), .A2(n_160), .B(n_158), .Y(n_804) );
A2O1A1Ixp33_ASAP7_75t_L g805 ( .A1(n_638), .A2(n_67), .B(n_68), .C(n_69), .Y(n_805) );
AO31x2_ASAP7_75t_L g806 ( .A1(n_694), .A2(n_69), .A3(n_70), .B(n_71), .Y(n_806) );
BUFx2_ASAP7_75t_L g807 ( .A(n_644), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_664), .Y(n_808) );
OAI222xp33_ASAP7_75t_L g809 ( .A1(n_722), .A2(n_70), .B1(n_71), .B2(n_72), .C1(n_73), .C2(n_74), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g810 ( .A1(n_680), .A2(n_162), .B(n_161), .Y(n_810) );
O2A1O1Ixp33_ASAP7_75t_L g811 ( .A1(n_663), .A2(n_653), .B(n_668), .C(n_621), .Y(n_811) );
BUFx2_ASAP7_75t_L g812 ( .A(n_687), .Y(n_812) );
OR2x2_ASAP7_75t_L g813 ( .A(n_627), .B(n_72), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_679), .A2(n_76), .B1(n_77), .B2(n_79), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_633), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_670), .Y(n_816) );
INVx2_ASAP7_75t_SL g817 ( .A(n_613), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_666), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_681), .A2(n_77), .B1(n_79), .B2(n_80), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_658), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_820) );
AND2x2_ASAP7_75t_SL g821 ( .A(n_697), .B(n_81), .Y(n_821) );
AO31x2_ASAP7_75t_L g822 ( .A1(n_668), .A2(n_83), .A3(n_84), .B(n_85), .Y(n_822) );
AO31x2_ASAP7_75t_L g823 ( .A1(n_719), .A2(n_84), .A3(n_85), .B(n_86), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_624), .A2(n_86), .B1(n_87), .B2(n_88), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_647), .B(n_88), .Y(n_825) );
OAI21xp5_ASAP7_75t_L g826 ( .A1(n_727), .A2(n_196), .B(n_256), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_651), .B(n_89), .Y(n_827) );
OR2x2_ASAP7_75t_L g828 ( .A(n_706), .B(n_89), .Y(n_828) );
OAI22xp33_ASAP7_75t_L g829 ( .A1(n_639), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_611), .B(n_90), .Y(n_830) );
BUFx6f_ASAP7_75t_L g831 ( .A(n_645), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_666), .B(n_91), .Y(n_832) );
INVx4_ASAP7_75t_L g833 ( .A(n_645), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_655), .Y(n_834) );
AO31x2_ASAP7_75t_L g835 ( .A1(n_636), .A2(n_93), .A3(n_95), .B(n_96), .Y(n_835) );
OAI21xp5_ASAP7_75t_L g836 ( .A1(n_699), .A2(n_199), .B(n_254), .Y(n_836) );
AOI221xp5_ASAP7_75t_L g837 ( .A1(n_702), .A2(n_95), .B1(n_97), .B2(n_98), .C(n_99), .Y(n_837) );
OR2x6_ASAP7_75t_L g838 ( .A(n_707), .B(n_97), .Y(n_838) );
INVx8_ASAP7_75t_L g839 ( .A(n_661), .Y(n_839) );
O2A1O1Ixp33_ASAP7_75t_SL g840 ( .A1(n_721), .A2(n_198), .B(n_251), .C(n_249), .Y(n_840) );
A2O1A1Ixp33_ASAP7_75t_L g841 ( .A1(n_698), .A2(n_100), .B(n_101), .C(n_102), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_615), .B(n_102), .Y(n_842) );
AO31x2_ASAP7_75t_L g843 ( .A1(n_708), .A2(n_103), .A3(n_106), .B(n_107), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_674), .B(n_106), .Y(n_844) );
O2A1O1Ixp33_ASAP7_75t_L g845 ( .A1(n_688), .A2(n_107), .B(n_108), .C(n_109), .Y(n_845) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_693), .B(n_109), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_718), .B(n_110), .Y(n_847) );
BUFx2_ASAP7_75t_L g848 ( .A(n_700), .Y(n_848) );
A2O1A1Ixp33_ASAP7_75t_L g849 ( .A1(n_701), .A2(n_113), .B(n_114), .C(n_115), .Y(n_849) );
NOR2xp33_ASAP7_75t_SL g850 ( .A(n_661), .B(n_114), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_692), .B(n_115), .Y(n_851) );
OAI22xp5_ASAP7_75t_SL g852 ( .A1(n_729), .A2(n_676), .B1(n_642), .B2(n_657), .Y(n_852) );
AOI221xp5_ASAP7_75t_L g853 ( .A1(n_695), .A2(n_116), .B1(n_117), .B2(n_118), .C(n_119), .Y(n_853) );
AO22x1_ASAP7_75t_L g854 ( .A1(n_729), .A2(n_116), .B1(n_117), .B2(n_118), .Y(n_854) );
BUFx2_ASAP7_75t_L g855 ( .A(n_661), .Y(n_855) );
AOI22xp5_ASAP7_75t_L g856 ( .A1(n_637), .A2(n_120), .B1(n_121), .B2(n_122), .Y(n_856) );
INVx1_ASAP7_75t_SL g857 ( .A(n_659), .Y(n_857) );
INVx4_ASAP7_75t_L g858 ( .A(n_660), .Y(n_858) );
INVx2_ASAP7_75t_SL g859 ( .A(n_708), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_708), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_716), .A2(n_120), .B1(n_122), .B2(n_123), .Y(n_861) );
A2O1A1Ixp33_ASAP7_75t_L g862 ( .A1(n_683), .A2(n_123), .B(n_124), .C(n_125), .Y(n_862) );
INVxp67_ASAP7_75t_SL g863 ( .A(n_614), .Y(n_863) );
BUFx8_ASAP7_75t_L g864 ( .A(n_726), .Y(n_864) );
BUFx12f_ASAP7_75t_L g865 ( .A(n_712), .Y(n_865) );
AOI21xp5_ASAP7_75t_L g866 ( .A1(n_724), .A2(n_169), .B(n_172), .Y(n_866) );
INVx3_ASAP7_75t_L g867 ( .A(n_689), .Y(n_867) );
A2O1A1Ixp33_ASAP7_75t_L g868 ( .A1(n_683), .A2(n_176), .B(n_177), .C(n_182), .Y(n_868) );
INVx3_ASAP7_75t_L g869 ( .A(n_689), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_682), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_682), .Y(n_871) );
BUFx2_ASAP7_75t_L g872 ( .A(n_614), .Y(n_872) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_614), .Y(n_873) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_872), .Y(n_874) );
AOI21xp5_ASAP7_75t_L g875 ( .A1(n_797), .A2(n_208), .B(n_212), .Y(n_875) );
INVxp67_ASAP7_75t_L g876 ( .A(n_863), .Y(n_876) );
INVx1_ASAP7_75t_SL g877 ( .A(n_752), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_731), .Y(n_878) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_873), .B(n_213), .Y(n_879) );
INVx2_ASAP7_75t_L g880 ( .A(n_737), .Y(n_880) );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_741), .A2(n_216), .B1(n_217), .B2(n_219), .C(n_220), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_870), .Y(n_882) );
BUFx8_ASAP7_75t_L g883 ( .A(n_747), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_734), .A2(n_226), .B1(n_227), .B2(n_228), .Y(n_884) );
AND2x4_ASAP7_75t_L g885 ( .A(n_740), .B(n_787), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_753), .B(n_236), .Y(n_886) );
AND2x4_ASAP7_75t_L g887 ( .A(n_787), .B(n_237), .Y(n_887) );
AOI221xp5_ASAP7_75t_L g888 ( .A1(n_816), .A2(n_272), .B1(n_743), .B2(n_770), .C(n_774), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_871), .Y(n_889) );
OAI21xp5_ASAP7_75t_L g890 ( .A1(n_762), .A2(n_764), .B(n_844), .Y(n_890) );
INVx1_ASAP7_75t_SL g891 ( .A(n_733), .Y(n_891) );
OR2x6_ASAP7_75t_L g892 ( .A(n_865), .B(n_795), .Y(n_892) );
BUFx2_ASAP7_75t_L g893 ( .A(n_864), .Y(n_893) );
INVxp67_ASAP7_75t_SL g894 ( .A(n_864), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_760), .Y(n_895) );
CKINVDCx5p33_ASAP7_75t_R g896 ( .A(n_754), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_791), .Y(n_897) );
BUFx4f_ASAP7_75t_SL g898 ( .A(n_798), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_736), .Y(n_899) );
A2O1A1Ixp33_ASAP7_75t_L g900 ( .A1(n_846), .A2(n_845), .B(n_825), .C(n_766), .Y(n_900) );
NAND2xp5_ASAP7_75t_SL g901 ( .A(n_812), .B(n_850), .Y(n_901) );
OR2x2_ASAP7_75t_L g902 ( .A(n_732), .B(n_780), .Y(n_902) );
AOI222xp33_ASAP7_75t_L g903 ( .A1(n_821), .A2(n_735), .B1(n_834), .B2(n_807), .C1(n_749), .C2(n_827), .Y(n_903) );
CKINVDCx11_ASAP7_75t_R g904 ( .A(n_732), .Y(n_904) );
HB1xp67_ASAP7_75t_L g905 ( .A(n_756), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_758), .Y(n_906) );
NOR2xp33_ASAP7_75t_L g907 ( .A(n_792), .B(n_817), .Y(n_907) );
HB1xp67_ASAP7_75t_L g908 ( .A(n_756), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_818), .B(n_746), .Y(n_909) );
INVx3_ASAP7_75t_L g910 ( .A(n_839), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_767), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_801), .Y(n_912) );
OAI221xp5_ASAP7_75t_L g913 ( .A1(n_761), .A2(n_838), .B1(n_782), .B2(n_763), .C(n_842), .Y(n_913) );
OAI22xp33_ASAP7_75t_L g914 ( .A1(n_838), .A2(n_783), .B1(n_802), .B2(n_801), .Y(n_914) );
AO31x2_ASAP7_75t_L g915 ( .A1(n_751), .A2(n_748), .A3(n_868), .B(n_810), .Y(n_915) );
INVx3_ASAP7_75t_L g916 ( .A(n_839), .Y(n_916) );
AND2x4_ASAP7_75t_L g917 ( .A(n_867), .B(n_869), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_738), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_848), .B(n_867), .Y(n_919) );
OR2x6_ASAP7_75t_L g920 ( .A(n_869), .B(n_854), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_745), .B(n_813), .Y(n_921) );
AO21x2_ASAP7_75t_L g922 ( .A1(n_836), .A2(n_826), .B(n_768), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_802), .Y(n_923) );
OAI22x1_ASAP7_75t_L g924 ( .A1(n_800), .A2(n_856), .B1(n_765), .B2(n_820), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_800), .A2(n_828), .B1(n_856), .B2(n_784), .Y(n_925) );
AO31x2_ASAP7_75t_L g926 ( .A1(n_804), .A2(n_781), .A3(n_779), .B(n_862), .Y(n_926) );
AOI22xp33_ASAP7_75t_SL g927 ( .A1(n_830), .A2(n_814), .B1(n_777), .B2(n_824), .Y(n_927) );
AOI22xp5_ASAP7_75t_L g928 ( .A1(n_794), .A2(n_829), .B1(n_790), .B2(n_785), .Y(n_928) );
INVx3_ASAP7_75t_L g929 ( .A(n_769), .Y(n_929) );
HB1xp67_ASAP7_75t_L g930 ( .A(n_765), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_757), .B(n_815), .Y(n_931) );
OAI221xp5_ASAP7_75t_L g932 ( .A1(n_786), .A2(n_805), .B1(n_832), .B2(n_819), .C(n_851), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_822), .Y(n_933) );
AOI211xp5_ASAP7_75t_L g934 ( .A1(n_744), .A2(n_809), .B(n_837), .C(n_853), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_822), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_775), .B(n_857), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_776), .Y(n_937) );
OR2x6_ASAP7_75t_L g938 ( .A(n_769), .B(n_796), .Y(n_938) );
HB1xp67_ASAP7_75t_L g939 ( .A(n_796), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_776), .Y(n_940) );
AOI21xp33_ASAP7_75t_L g941 ( .A1(n_847), .A2(n_803), .B(n_789), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_776), .Y(n_942) );
CKINVDCx11_ASAP7_75t_R g943 ( .A(n_772), .Y(n_943) );
OAI21xp5_ASAP7_75t_L g944 ( .A1(n_841), .A2(n_849), .B(n_866), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_771), .B(n_808), .Y(n_945) );
BUFx6f_ASAP7_75t_L g946 ( .A(n_759), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_788), .Y(n_947) );
OAI21xp33_ASAP7_75t_L g948 ( .A1(n_773), .A2(n_861), .B(n_755), .Y(n_948) );
OR2x6_ASAP7_75t_L g949 ( .A(n_852), .B(n_833), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_858), .B(n_855), .Y(n_950) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_858), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_788), .B(n_806), .Y(n_952) );
OR2x2_ASAP7_75t_L g953 ( .A(n_806), .B(n_788), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_835), .Y(n_954) );
OR2x2_ASAP7_75t_L g955 ( .A(n_806), .B(n_742), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g956 ( .A1(n_840), .A2(n_831), .B(n_799), .Y(n_956) );
AOI22xp33_ASAP7_75t_SL g957 ( .A1(n_823), .A2(n_742), .B1(n_739), .B2(n_835), .Y(n_957) );
AOI21xp5_ASAP7_75t_L g958 ( .A1(n_739), .A2(n_793), .B(n_843), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_823), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_823), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_843), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_793), .B(n_614), .Y(n_962) );
OAI21xp5_ASAP7_75t_L g963 ( .A1(n_859), .A2(n_860), .B(n_665), .Y(n_963) );
OR2x6_ASAP7_75t_SL g964 ( .A(n_754), .B(n_519), .Y(n_964) );
OR2x2_ASAP7_75t_L g965 ( .A(n_872), .B(n_863), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_741), .B(n_614), .Y(n_966) );
AND2x2_ASAP7_75t_L g967 ( .A(n_863), .B(n_614), .Y(n_967) );
AO31x2_ASAP7_75t_L g968 ( .A1(n_860), .A2(n_751), .A3(n_748), .B(n_778), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_731), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_863), .B(n_614), .Y(n_970) );
OR2x2_ASAP7_75t_L g971 ( .A(n_872), .B(n_863), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_731), .Y(n_972) );
OR2x6_ASAP7_75t_L g973 ( .A(n_747), .B(n_865), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_731), .Y(n_974) );
A2O1A1Ixp33_ASAP7_75t_L g975 ( .A1(n_811), .A2(n_750), .B(n_846), .C(n_845), .Y(n_975) );
NAND2xp5_ASAP7_75t_SL g976 ( .A(n_797), .B(n_723), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_797), .A2(n_665), .B1(n_605), .B2(n_734), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_731), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_863), .B(n_614), .Y(n_979) );
CKINVDCx16_ASAP7_75t_R g980 ( .A(n_747), .Y(n_980) );
CKINVDCx6p67_ASAP7_75t_R g981 ( .A(n_747), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_741), .A2(n_556), .B1(n_561), .B2(n_554), .Y(n_982) );
BUFx3_ASAP7_75t_L g983 ( .A(n_747), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_741), .B(n_614), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_737), .Y(n_985) );
OAI221xp5_ASAP7_75t_L g986 ( .A1(n_741), .A2(n_628), .B1(n_561), .B2(n_863), .C(n_510), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_872), .B(n_863), .Y(n_987) );
OAI221xp5_ASAP7_75t_L g988 ( .A1(n_741), .A2(n_628), .B1(n_561), .B2(n_863), .C(n_510), .Y(n_988) );
A2O1A1Ixp33_ASAP7_75t_L g989 ( .A1(n_811), .A2(n_750), .B(n_846), .C(n_845), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_863), .B(n_614), .Y(n_990) );
A2O1A1Ixp33_ASAP7_75t_L g991 ( .A1(n_811), .A2(n_750), .B(n_846), .C(n_845), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_741), .B(n_614), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_741), .B(n_614), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_731), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_731), .Y(n_995) );
INVx3_ASAP7_75t_L g996 ( .A(n_747), .Y(n_996) );
INVx2_ASAP7_75t_L g997 ( .A(n_737), .Y(n_997) );
INVx2_ASAP7_75t_L g998 ( .A(n_737), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_741), .A2(n_556), .B1(n_561), .B2(n_554), .Y(n_999) );
OAI21xp5_ASAP7_75t_L g1000 ( .A1(n_859), .A2(n_860), .B(n_665), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_872), .Y(n_1001) );
CKINVDCx5p33_ASAP7_75t_R g1002 ( .A(n_747), .Y(n_1002) );
OR2x2_ASAP7_75t_L g1003 ( .A(n_872), .B(n_863), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_741), .B(n_614), .Y(n_1004) );
OR2x6_ASAP7_75t_L g1005 ( .A(n_747), .B(n_865), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_731), .Y(n_1006) );
HB1xp67_ASAP7_75t_L g1007 ( .A(n_872), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_731), .Y(n_1008) );
NOR2xp33_ASAP7_75t_L g1009 ( .A(n_872), .B(n_564), .Y(n_1009) );
CKINVDCx5p33_ASAP7_75t_R g1010 ( .A(n_883), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_966), .B(n_984), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_992), .B(n_993), .Y(n_1012) );
OA21x2_ASAP7_75t_L g1013 ( .A1(n_958), .A2(n_961), .B(n_954), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_918), .B(n_880), .Y(n_1014) );
OAI211xp5_ASAP7_75t_SL g1015 ( .A1(n_982), .A2(n_999), .B(n_903), .C(n_913), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_1004), .B(n_967), .Y(n_1016) );
AOI221xp5_ASAP7_75t_L g1017 ( .A1(n_986), .A2(n_988), .B1(n_977), .B2(n_914), .C(n_1009), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_970), .B(n_979), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_882), .B(n_985), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_940), .Y(n_1020) );
AO21x2_ASAP7_75t_L g1021 ( .A1(n_942), .A2(n_947), .B(n_963), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g1022 ( .A(n_965), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_903), .A2(n_923), .B1(n_912), .B2(n_888), .Y(n_1023) );
AND2x4_ASAP7_75t_L g1024 ( .A(n_963), .B(n_1000), .Y(n_1024) );
AOI221xp5_ASAP7_75t_L g1025 ( .A1(n_925), .A2(n_921), .B1(n_924), .B2(n_975), .C(n_989), .Y(n_1025) );
AND2x4_ASAP7_75t_L g1026 ( .A(n_1000), .B(n_949), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_933), .Y(n_1027) );
AND2x4_ASAP7_75t_L g1028 ( .A(n_949), .B(n_946), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_935), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_997), .B(n_998), .Y(n_1030) );
INVx2_ASAP7_75t_SL g1031 ( .A(n_973), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_952), .Y(n_1032) );
NOR2x1_ASAP7_75t_L g1033 ( .A(n_920), .B(n_949), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_953), .Y(n_1034) );
INVx2_ASAP7_75t_SL g1035 ( .A(n_973), .Y(n_1035) );
BUFx2_ASAP7_75t_L g1036 ( .A(n_951), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_990), .B(n_878), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_955), .Y(n_1038) );
NOR2x1_ASAP7_75t_L g1039 ( .A(n_920), .B(n_959), .Y(n_1039) );
BUFx3_ASAP7_75t_L g1040 ( .A(n_885), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_960), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_962), .Y(n_1042) );
BUFx4f_ASAP7_75t_L g1043 ( .A(n_887), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_889), .B(n_911), .Y(n_1044) );
HB1xp67_ASAP7_75t_L g1045 ( .A(n_971), .Y(n_1045) );
BUFx3_ASAP7_75t_L g1046 ( .A(n_885), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_899), .Y(n_1047) );
AO21x2_ASAP7_75t_L g1048 ( .A1(n_922), .A2(n_944), .B(n_956), .Y(n_1048) );
BUFx3_ASAP7_75t_L g1049 ( .A(n_910), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_906), .B(n_895), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_1008), .B(n_969), .Y(n_1051) );
NOR2xp33_ASAP7_75t_L g1052 ( .A(n_964), .B(n_945), .Y(n_1052) );
OR2x2_ASAP7_75t_L g1053 ( .A(n_877), .B(n_987), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_930), .Y(n_1054) );
AO21x2_ASAP7_75t_L g1055 ( .A1(n_991), .A2(n_890), .B(n_948), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_897), .B(n_877), .Y(n_1056) );
AO21x2_ASAP7_75t_L g1057 ( .A1(n_941), .A2(n_900), .B(n_928), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_957), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_920), .A2(n_976), .B1(n_927), .B2(n_932), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_1003), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_936), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_972), .Y(n_1062) );
AOI21xp5_ASAP7_75t_SL g1063 ( .A1(n_887), .A2(n_884), .B(n_875), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_974), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_978), .B(n_1006), .Y(n_1065) );
OAI31xp33_ASAP7_75t_L g1066 ( .A1(n_876), .A2(n_874), .A3(n_1001), .B(n_1007), .Y(n_1066) );
OAI21xp5_ASAP7_75t_L g1067 ( .A1(n_934), .A2(n_881), .B(n_909), .Y(n_1067) );
HB1xp67_ASAP7_75t_L g1068 ( .A(n_919), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_994), .Y(n_1069) );
OAI21x1_ASAP7_75t_L g1070 ( .A1(n_929), .A2(n_901), .B(n_950), .Y(n_1070) );
HB1xp67_ASAP7_75t_L g1071 ( .A(n_902), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_995), .B(n_939), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_938), .B(n_931), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_938), .B(n_886), .Y(n_1074) );
AO21x2_ASAP7_75t_L g1075 ( .A1(n_968), .A2(n_915), .B(n_926), .Y(n_1075) );
INVx2_ASAP7_75t_L g1076 ( .A(n_968), .Y(n_1076) );
INVx3_ASAP7_75t_L g1077 ( .A(n_926), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_926), .Y(n_1078) );
AO21x2_ASAP7_75t_L g1079 ( .A1(n_915), .A2(n_879), .B(n_934), .Y(n_1079) );
AO21x2_ASAP7_75t_L g1080 ( .A1(n_907), .A2(n_905), .B(n_908), .Y(n_1080) );
OAI21xp33_ASAP7_75t_L g1081 ( .A1(n_891), .A2(n_892), .B(n_1005), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_910), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_916), .B(n_891), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_917), .B(n_892), .Y(n_1084) );
INVx2_ASAP7_75t_L g1085 ( .A(n_917), .Y(n_1085) );
OA21x2_ASAP7_75t_L g1086 ( .A1(n_894), .A2(n_893), .B(n_1002), .Y(n_1086) );
AND2x4_ASAP7_75t_L g1087 ( .A(n_892), .B(n_973), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_996), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_996), .B(n_980), .Y(n_1089) );
INVx2_ASAP7_75t_L g1090 ( .A(n_1005), .Y(n_1090) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_1005), .B(n_983), .Y(n_1091) );
OA21x2_ASAP7_75t_L g1092 ( .A1(n_896), .A2(n_904), .B(n_981), .Y(n_1092) );
NOR2xp33_ASAP7_75t_L g1093 ( .A(n_883), .B(n_898), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_943), .B(n_966), .Y(n_1094) );
NAND3xp33_ASAP7_75t_L g1095 ( .A(n_957), .B(n_903), .C(n_958), .Y(n_1095) );
INVx4_ASAP7_75t_L g1096 ( .A(n_887), .Y(n_1096) );
OR2x6_ASAP7_75t_L g1097 ( .A(n_949), .B(n_963), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_914), .A2(n_903), .B1(n_988), .B2(n_986), .Y(n_1098) );
BUFx2_ASAP7_75t_L g1099 ( .A(n_963), .Y(n_1099) );
AOI22xp33_ASAP7_75t_SL g1100 ( .A1(n_977), .A2(n_821), .B1(n_783), .B2(n_519), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_937), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_918), .B(n_880), .Y(n_1102) );
BUFx2_ASAP7_75t_L g1103 ( .A(n_963), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1104 ( .A(n_965), .Y(n_1104) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_912), .B(n_923), .Y(n_1105) );
HB1xp67_ASAP7_75t_L g1106 ( .A(n_1036), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1032), .B(n_1042), .Y(n_1107) );
HB1xp67_ASAP7_75t_L g1108 ( .A(n_1036), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1020), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1032), .B(n_1042), .Y(n_1110) );
INVx2_ASAP7_75t_SL g1111 ( .A(n_1043), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1058), .B(n_1034), .Y(n_1112) );
BUFx3_ASAP7_75t_L g1113 ( .A(n_1040), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1058), .B(n_1034), .Y(n_1114) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_1096), .Y(n_1115) );
HB1xp67_ASAP7_75t_L g1116 ( .A(n_1022), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g1117 ( .A(n_1045), .Y(n_1117) );
NAND2x1_ASAP7_75t_L g1118 ( .A(n_1096), .B(n_1033), .Y(n_1118) );
BUFx2_ASAP7_75t_L g1119 ( .A(n_1096), .Y(n_1119) );
OAI33xp33_ASAP7_75t_L g1120 ( .A1(n_1015), .A2(n_1054), .A3(n_1095), .B1(n_1053), .B2(n_1069), .B3(n_1064), .Y(n_1120) );
NAND2x1_ASAP7_75t_L g1121 ( .A(n_1096), .B(n_1033), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_1060), .Y(n_1122) );
BUFx2_ASAP7_75t_L g1123 ( .A(n_1043), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1038), .B(n_1024), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1038), .B(n_1024), .Y(n_1125) );
NAND4xp25_ASAP7_75t_L g1126 ( .A(n_1098), .B(n_1017), .C(n_1100), .D(n_1025), .Y(n_1126) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_1104), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1011), .B(n_1012), .Y(n_1128) );
AND2x4_ASAP7_75t_SL g1129 ( .A(n_1087), .B(n_1091), .Y(n_1129) );
AND2x4_ASAP7_75t_L g1130 ( .A(n_1039), .B(n_1026), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1024), .B(n_1055), .Y(n_1131) );
OR2x2_ASAP7_75t_L g1132 ( .A(n_1105), .B(n_1053), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1016), .B(n_1050), .Y(n_1133) );
NAND2x1_ASAP7_75t_L g1134 ( .A(n_1097), .B(n_1039), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1024), .B(n_1055), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_1050), .B(n_1061), .Y(n_1136) );
INVx5_ASAP7_75t_SL g1137 ( .A(n_1087), .Y(n_1137) );
OR2x2_ASAP7_75t_L g1138 ( .A(n_1095), .B(n_1041), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1055), .B(n_1041), .Y(n_1139) );
INVx2_ASAP7_75t_SL g1140 ( .A(n_1043), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1044), .B(n_1027), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1044), .B(n_1029), .Y(n_1142) );
INVx3_ASAP7_75t_L g1143 ( .A(n_1043), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1065), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1065), .Y(n_1145) );
AND2x4_ASAP7_75t_L g1146 ( .A(n_1026), .B(n_1028), .Y(n_1146) );
OR2x6_ASAP7_75t_L g1147 ( .A(n_1097), .B(n_1026), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1101), .B(n_1047), .Y(n_1148) );
HB1xp67_ASAP7_75t_L g1149 ( .A(n_1068), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1047), .B(n_1014), .Y(n_1150) );
OR2x6_ASAP7_75t_L g1151 ( .A(n_1097), .B(n_1026), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1014), .B(n_1019), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1062), .Y(n_1153) );
HB1xp67_ASAP7_75t_L g1154 ( .A(n_1056), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1019), .B(n_1030), .Y(n_1155) );
AOI22xp33_ASAP7_75t_SL g1156 ( .A1(n_1087), .A2(n_1052), .B1(n_1097), .B2(n_1040), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1080), .B(n_1097), .Y(n_1157) );
NAND2x1p5_ASAP7_75t_L g1158 ( .A(n_1040), .B(n_1046), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1080), .B(n_1061), .Y(n_1159) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1080), .B(n_1099), .Y(n_1160) );
INVx1_ASAP7_75t_SL g1161 ( .A(n_1089), .Y(n_1161) );
INVx5_ASAP7_75t_SL g1162 ( .A(n_1087), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1023), .B(n_1037), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1062), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1102), .B(n_1099), .Y(n_1165) );
HB1xp67_ASAP7_75t_L g1166 ( .A(n_1056), .Y(n_1166) );
OR2x2_ASAP7_75t_L g1167 ( .A(n_1154), .B(n_1103), .Y(n_1167) );
INVx1_ASAP7_75t_SL g1168 ( .A(n_1161), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1141), .B(n_1064), .Y(n_1169) );
NOR2xp33_ASAP7_75t_L g1170 ( .A(n_1133), .B(n_1094), .Y(n_1170) );
CKINVDCx16_ASAP7_75t_R g1171 ( .A(n_1123), .Y(n_1171) );
NAND2xp5_ASAP7_75t_SL g1172 ( .A(n_1156), .B(n_1081), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1124), .B(n_1077), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1125), .B(n_1077), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1141), .B(n_1069), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1131), .B(n_1077), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1131), .B(n_1078), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1135), .B(n_1078), .Y(n_1178) );
NAND2xp33_ASAP7_75t_L g1179 ( .A(n_1111), .B(n_1081), .Y(n_1179) );
HB1xp67_ASAP7_75t_L g1180 ( .A(n_1106), .Y(n_1180) );
INVxp67_ASAP7_75t_L g1181 ( .A(n_1149), .Y(n_1181) );
OAI21xp33_ASAP7_75t_L g1182 ( .A1(n_1126), .A2(n_1059), .B(n_1067), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1135), .B(n_1021), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1109), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1185 ( .A(n_1166), .B(n_1021), .Y(n_1185) );
BUFx3_ASAP7_75t_L g1186 ( .A(n_1113), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1165), .B(n_1021), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1142), .B(n_1152), .Y(n_1188) );
NOR2x1_ASAP7_75t_L g1189 ( .A(n_1113), .B(n_1046), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1109), .Y(n_1190) );
NOR2xp67_ASAP7_75t_L g1191 ( .A(n_1138), .B(n_1076), .Y(n_1191) );
HB1xp67_ASAP7_75t_L g1192 ( .A(n_1108), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1107), .B(n_1013), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1110), .B(n_1013), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1132), .B(n_1076), .Y(n_1195) );
BUFx2_ASAP7_75t_L g1196 ( .A(n_1115), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1110), .B(n_1075), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1112), .B(n_1075), .Y(n_1198) );
INVxp67_ASAP7_75t_SL g1199 ( .A(n_1116), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1152), .B(n_1072), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1155), .B(n_1071), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1114), .B(n_1048), .Y(n_1202) );
NOR2x1_ASAP7_75t_L g1203 ( .A(n_1118), .B(n_1028), .Y(n_1203) );
HB1xp67_ASAP7_75t_L g1204 ( .A(n_1117), .Y(n_1204) );
OR2x6_ASAP7_75t_L g1205 ( .A(n_1147), .B(n_1063), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1148), .B(n_1048), .Y(n_1206) );
NAND2x1_ASAP7_75t_SL g1207 ( .A(n_1143), .B(n_1028), .Y(n_1207) );
INVx2_ASAP7_75t_SL g1208 ( .A(n_1186), .Y(n_1208) );
NOR2xp67_ASAP7_75t_SL g1209 ( .A(n_1171), .B(n_1063), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1193), .B(n_1139), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1204), .Y(n_1211) );
HB1xp67_ASAP7_75t_L g1212 ( .A(n_1180), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1188), .B(n_1122), .Y(n_1213) );
INVxp33_ASAP7_75t_L g1214 ( .A(n_1170), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1184), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1190), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1190), .Y(n_1217) );
INVxp67_ASAP7_75t_L g1218 ( .A(n_1199), .Y(n_1218) );
INVxp67_ASAP7_75t_L g1219 ( .A(n_1192), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1193), .B(n_1139), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1197), .B(n_1127), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1197), .B(n_1144), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1194), .B(n_1151), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1194), .B(n_1151), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1176), .B(n_1151), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1169), .B(n_1145), .Y(n_1226) );
NAND2xp33_ASAP7_75t_L g1227 ( .A(n_1172), .B(n_1111), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1176), .B(n_1151), .Y(n_1228) );
AND2x4_ASAP7_75t_L g1229 ( .A(n_1205), .B(n_1146), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1175), .B(n_1150), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1177), .B(n_1146), .Y(n_1231) );
AND2x4_ASAP7_75t_L g1232 ( .A(n_1205), .B(n_1146), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1177), .B(n_1148), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1178), .B(n_1130), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1167), .B(n_1159), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1200), .B(n_1150), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1178), .B(n_1130), .Y(n_1237) );
BUFx2_ASAP7_75t_L g1238 ( .A(n_1196), .Y(n_1238) );
AND2x4_ASAP7_75t_L g1239 ( .A(n_1205), .B(n_1130), .Y(n_1239) );
NOR3xp33_ASAP7_75t_L g1240 ( .A(n_1182), .B(n_1120), .C(n_1128), .Y(n_1240) );
AND2x4_ASAP7_75t_L g1241 ( .A(n_1205), .B(n_1157), .Y(n_1241) );
INVxp67_ASAP7_75t_SL g1242 ( .A(n_1196), .Y(n_1242) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1167), .B(n_1195), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1195), .B(n_1159), .Y(n_1244) );
INVxp67_ASAP7_75t_L g1245 ( .A(n_1168), .Y(n_1245) );
INVx1_ASAP7_75t_SL g1246 ( .A(n_1238), .Y(n_1246) );
NOR2x1_ASAP7_75t_L g1247 ( .A(n_1227), .B(n_1179), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1215), .Y(n_1248) );
NAND2x1p5_ASAP7_75t_L g1249 ( .A(n_1209), .B(n_1115), .Y(n_1249) );
OR2x2_ASAP7_75t_L g1250 ( .A(n_1243), .B(n_1185), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1210), .B(n_1183), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1210), .B(n_1187), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1233), .B(n_1181), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1215), .Y(n_1254) );
HB1xp67_ASAP7_75t_L g1255 ( .A(n_1238), .Y(n_1255) );
INVxp67_ASAP7_75t_L g1256 ( .A(n_1212), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1220), .B(n_1187), .Y(n_1257) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1216), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1223), .B(n_1206), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1211), .B(n_1202), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1221), .B(n_1206), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_1243), .B(n_1185), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1216), .Y(n_1263) );
OAI21xp33_ASAP7_75t_L g1264 ( .A1(n_1240), .A2(n_1138), .B(n_1201), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1223), .B(n_1173), .Y(n_1265) );
NOR2x1_ASAP7_75t_L g1266 ( .A(n_1227), .B(n_1189), .Y(n_1266) );
INVxp67_ASAP7_75t_SL g1267 ( .A(n_1242), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1224), .B(n_1173), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1217), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1224), .B(n_1174), .Y(n_1270) );
HB1xp67_ASAP7_75t_L g1271 ( .A(n_1218), .Y(n_1271) );
INVx2_ASAP7_75t_SL g1272 ( .A(n_1208), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1222), .B(n_1198), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1217), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1250), .Y(n_1275) );
NAND2xp5_ASAP7_75t_SL g1276 ( .A(n_1247), .B(n_1208), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1264), .B(n_1219), .Y(n_1277) );
NAND3xp33_ASAP7_75t_L g1278 ( .A(n_1264), .B(n_1245), .C(n_1209), .Y(n_1278) );
OR2x2_ASAP7_75t_L g1279 ( .A(n_1250), .B(n_1235), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_1251), .B(n_1213), .Y(n_1280) );
INVxp67_ASAP7_75t_SL g1281 ( .A(n_1255), .Y(n_1281) );
NAND4xp25_ASAP7_75t_L g1282 ( .A(n_1247), .B(n_1066), .C(n_1163), .D(n_1093), .Y(n_1282) );
AOI222xp33_ASAP7_75t_L g1283 ( .A1(n_1256), .A2(n_1214), .B1(n_1031), .B2(n_1035), .C1(n_1226), .C2(n_1136), .Y(n_1283) );
NOR2x1_ASAP7_75t_L g1284 ( .A(n_1266), .B(n_1092), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1262), .Y(n_1285) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_1249), .A2(n_1230), .B1(n_1236), .B2(n_1162), .Y(n_1286) );
OAI221xp5_ASAP7_75t_L g1287 ( .A1(n_1249), .A2(n_1271), .B1(n_1267), .B2(n_1272), .C(n_1246), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1248), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1252), .B(n_1235), .Y(n_1289) );
A2O1A1Ixp33_ASAP7_75t_L g1290 ( .A1(n_1272), .A2(n_1129), .B(n_1091), .C(n_1121), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1252), .B(n_1198), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1248), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1254), .Y(n_1293) );
NAND5xp2_ASAP7_75t_L g1294 ( .A(n_1283), .B(n_1089), .C(n_1158), .D(n_1123), .E(n_1084), .Y(n_1294) );
OAI211xp5_ASAP7_75t_SL g1295 ( .A1(n_1284), .A2(n_1253), .B(n_1260), .C(n_1090), .Y(n_1295) );
AOI32xp33_ASAP7_75t_L g1296 ( .A1(n_1276), .A2(n_1257), .A3(n_1268), .B1(n_1265), .B2(n_1270), .Y(n_1296) );
INVxp67_ASAP7_75t_L g1297 ( .A(n_1277), .Y(n_1297) );
OAI21xp5_ASAP7_75t_L g1298 ( .A1(n_1276), .A2(n_1092), .B(n_1191), .Y(n_1298) );
AOI221xp5_ASAP7_75t_L g1299 ( .A1(n_1282), .A2(n_1261), .B1(n_1273), .B2(n_1257), .C(n_1259), .Y(n_1299) );
OAI211xp5_ASAP7_75t_L g1300 ( .A1(n_1278), .A2(n_1092), .B(n_1086), .C(n_1207), .Y(n_1300) );
AOI221xp5_ASAP7_75t_L g1301 ( .A1(n_1287), .A2(n_1091), .B1(n_1274), .B2(n_1269), .C(n_1254), .Y(n_1301) );
AOI22xp5_ASAP7_75t_L g1302 ( .A1(n_1286), .A2(n_1241), .B1(n_1229), .B2(n_1232), .Y(n_1302) );
AOI222xp33_ASAP7_75t_L g1303 ( .A1(n_1281), .A2(n_1091), .B1(n_1259), .B2(n_1274), .C1(n_1263), .C2(n_1269), .Y(n_1303) );
A2O1A1Ixp33_ASAP7_75t_L g1304 ( .A1(n_1290), .A2(n_1129), .B(n_1232), .C(n_1229), .Y(n_1304) );
AOI222xp33_ASAP7_75t_L g1305 ( .A1(n_1275), .A2(n_1258), .B1(n_1263), .B2(n_1191), .C1(n_1241), .C2(n_1090), .Y(n_1305) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1279), .Y(n_1306) );
INVx2_ASAP7_75t_L g1307 ( .A(n_1285), .Y(n_1307) );
OR2x2_ASAP7_75t_L g1308 ( .A(n_1306), .B(n_1289), .Y(n_1308) );
AOI221xp5_ASAP7_75t_L g1309 ( .A1(n_1299), .A2(n_1293), .B1(n_1292), .B2(n_1288), .C(n_1280), .Y(n_1309) );
NAND3xp33_ASAP7_75t_SL g1310 ( .A(n_1300), .B(n_1010), .C(n_1119), .Y(n_1310) );
NAND2xp5_ASAP7_75t_SL g1311 ( .A(n_1296), .B(n_1186), .Y(n_1311) );
AOI221xp5_ASAP7_75t_L g1312 ( .A1(n_1297), .A2(n_1291), .B1(n_1258), .B2(n_1270), .C(n_1088), .Y(n_1312) );
OAI321xp33_ASAP7_75t_L g1313 ( .A1(n_1298), .A2(n_1160), .A3(n_1225), .B1(n_1228), .B2(n_1244), .C(n_1158), .Y(n_1313) );
NOR3xp33_ASAP7_75t_L g1314 ( .A(n_1301), .B(n_1088), .C(n_1083), .Y(n_1314) );
AOI221xp5_ASAP7_75t_SL g1315 ( .A1(n_1301), .A2(n_1231), .B1(n_1234), .B2(n_1237), .C(n_1083), .Y(n_1315) );
OAI211xp5_ASAP7_75t_SL g1316 ( .A1(n_1303), .A2(n_1018), .B(n_1203), .C(n_1143), .Y(n_1316) );
NAND4xp25_ASAP7_75t_L g1317 ( .A(n_1294), .B(n_1084), .C(n_1203), .D(n_1239), .Y(n_1317) );
NOR2x1_ASAP7_75t_L g1318 ( .A(n_1310), .B(n_1311), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1308), .Y(n_1319) );
NOR3xp33_ASAP7_75t_L g1320 ( .A(n_1313), .B(n_1295), .C(n_1304), .Y(n_1320) );
AOI22xp5_ASAP7_75t_L g1321 ( .A1(n_1315), .A2(n_1302), .B1(n_1305), .B2(n_1307), .Y(n_1321) );
NOR3xp33_ASAP7_75t_L g1322 ( .A(n_1316), .B(n_1082), .C(n_1051), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1312), .Y(n_1323) );
NOR3xp33_ASAP7_75t_L g1324 ( .A(n_1309), .B(n_1082), .C(n_1070), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1319), .Y(n_1325) );
NAND2xp5_ASAP7_75t_SL g1326 ( .A(n_1318), .B(n_1314), .Y(n_1326) );
NOR2xp67_ASAP7_75t_L g1327 ( .A(n_1321), .B(n_1317), .Y(n_1327) );
NAND5xp2_ASAP7_75t_L g1328 ( .A(n_1320), .B(n_1074), .C(n_1158), .D(n_1073), .E(n_1086), .Y(n_1328) );
NOR4xp25_ASAP7_75t_L g1329 ( .A(n_1323), .B(n_1085), .C(n_1153), .D(n_1164), .Y(n_1329) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1325), .B(n_1328), .Y(n_1330) );
NAND4xp25_ASAP7_75t_L g1331 ( .A(n_1327), .B(n_1324), .C(n_1322), .D(n_1143), .Y(n_1331) );
AOI22xp33_ASAP7_75t_SL g1332 ( .A1(n_1326), .A2(n_1137), .B1(n_1162), .B2(n_1119), .Y(n_1332) );
INVx3_ASAP7_75t_L g1333 ( .A(n_1330), .Y(n_1333) );
OAI22xp5_ASAP7_75t_L g1334 ( .A1(n_1332), .A2(n_1328), .B1(n_1329), .B2(n_1134), .Y(n_1334) );
OAI22xp5_ASAP7_75t_L g1335 ( .A1(n_1333), .A2(n_1331), .B1(n_1140), .B2(n_1160), .Y(n_1335) );
CKINVDCx20_ASAP7_75t_R g1336 ( .A(n_1334), .Y(n_1336) );
AOI21xp5_ASAP7_75t_L g1337 ( .A1(n_1336), .A2(n_1049), .B(n_1085), .Y(n_1337) );
XNOR2x1_ASAP7_75t_L g1338 ( .A(n_1337), .B(n_1335), .Y(n_1338) );
INVx3_ASAP7_75t_L g1339 ( .A(n_1338), .Y(n_1339) );
AOI22xp5_ASAP7_75t_L g1340 ( .A1(n_1339), .A2(n_1079), .B1(n_1028), .B2(n_1057), .Y(n_1340) );
endmodule