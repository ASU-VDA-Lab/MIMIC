module real_aes_17300_n_7 (n_4, n_0, n_3, n_5, n_2, n_6, n_1, n_7);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_6;
input n_1;
output n_7;
wire n_16;
wire n_17;
wire n_13;
wire n_15;
wire n_8;
wire n_9;
wire n_12;
wire n_14;
wire n_10;
wire n_11;
INVx2_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
A2O1A1Ixp33_ASAP7_75t_L g7 ( .A1(n_1), .A2(n_8), .B(n_13), .C(n_16), .Y(n_7) );
AND2x4_ASAP7_75t_L g16 ( .A(n_2), .B(n_17), .Y(n_16) );
INVx1_ASAP7_75t_L g12 ( .A(n_3), .Y(n_12) );
O2A1O1Ixp33_ASAP7_75t_L g13 ( .A1(n_4), .A2(n_8), .B(n_14), .C(n_15), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_4), .B(n_14), .Y(n_15) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx1_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
AND2x2_ASAP7_75t_L g8 ( .A(n_9), .B(n_11), .Y(n_8) );
INVx3_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
BUFx2_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
endmodule