module fake_netlist_5_435_n_202 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_32, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_202);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_32;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;

output n_202;

wire n_137;
wire n_168;
wire n_164;
wire n_91;
wire n_82;
wire n_122;
wire n_194;
wire n_142;
wire n_176;
wire n_140;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_184;
wire n_78;
wire n_65;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_189;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_197;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_195;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_193;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_192;
wire n_53;
wire n_160;
wire n_198;
wire n_188;
wire n_190;
wire n_201;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_154;
wire n_71;
wire n_148;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_183;
wire n_185;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_196;
wire n_99;
wire n_181;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_178;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_200;
wire n_87;
wire n_170;
wire n_150;
wire n_162;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_186;
wire n_199;
wire n_134;
wire n_187;
wire n_41;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_191;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_23),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVxp67_ASAP7_75t_SL g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVxp33_ASAP7_75t_SL g50 ( 
.A(n_21),
.Y(n_50)
);

INVxp67_ASAP7_75t_SL g51 ( 
.A(n_25),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_18),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_1),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_3),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_3),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_6),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_7),
.Y(n_75)
);

INVxp67_ASAP7_75t_SL g76 ( 
.A(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_8),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_13),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AOI21x1_ASAP7_75t_L g82 ( 
.A1(n_41),
.A2(n_17),
.B(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_45),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_40),
.Y(n_85)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_56),
.B1(n_57),
.B2(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_81),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_63),
.B(n_56),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_57),
.B1(n_51),
.B2(n_48),
.Y(n_98)
);

AND2x4_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_34),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_52),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_22),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_27),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_75),
.Y(n_104)
);

OR2x6_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_30),
.Y(n_105)
);

OAI21x1_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_82),
.B(n_79),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_68),
.Y(n_107)
);

OAI21x1_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_68),
.B(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_62),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_104),
.B(n_73),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_76),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_68),
.B(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_71),
.Y(n_118)
);

NOR2xp67_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_95),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_71),
.B(n_66),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

OAI21x1_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_67),
.B(n_31),
.Y(n_124)
);

NOR2xp67_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_101),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

NOR2xp67_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_98),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_89),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_96),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_89),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_105),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_90),
.B(n_87),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_105),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_96),
.Y(n_136)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_106),
.B(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_103),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_122),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_92),
.B(n_67),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_92),
.Y(n_141)
);

NOR2x1_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_86),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_86),
.B(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_123),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_125),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_113),
.Y(n_147)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_145),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_132),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_123),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_123),
.Y(n_154)
);

BUFx2_ASAP7_75t_SL g155 ( 
.A(n_127),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_120),
.B(n_121),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_139),
.B1(n_146),
.B2(n_127),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_135),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_135),
.B1(n_128),
.B2(n_127),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_127),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_131),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_134),
.B1(n_144),
.B2(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_139),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_134),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_172),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_154),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

OAI221xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_161),
.B1(n_148),
.B2(n_159),
.C(n_158),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_154),
.C(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_150),
.C(n_153),
.Y(n_190)
);

OAI321xp33_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_179),
.A3(n_150),
.B1(n_153),
.B2(n_162),
.C(n_147),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_SL g192 ( 
.A(n_186),
.B(n_187),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_147),
.C(n_182),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_148),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_193),
.B(n_191),
.Y(n_195)
);

OAI221xp5_ASAP7_75t_L g196 ( 
.A1(n_194),
.A2(n_189),
.B1(n_188),
.B2(n_142),
.C(n_182),
.Y(n_196)
);

NAND4xp75_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_143),
.C(n_178),
.D(n_175),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_178),
.A3(n_169),
.B1(n_168),
.B2(n_165),
.C1(n_166),
.C2(n_143),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

OAI22x1_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_196),
.B1(n_177),
.B2(n_137),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_155),
.B1(n_168),
.B2(n_169),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_137),
.B1(n_155),
.B2(n_199),
.Y(n_202)
);


endmodule