module real_aes_7110_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_13;
wire n_7;
wire n_8;
wire n_12;
wire n_9;
wire n_10;
wire n_11;
CKINVDCx20_ASAP7_75t_R g8 ( .A(n_0), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_1), .B(n_13), .Y(n_12) );
AOI221xp5_ASAP7_75t_L g6 ( .A1(n_2), .A2(n_4), .B1(n_7), .B2(n_11), .C(n_12), .Y(n_6) );
INVx1_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
INVx2_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
CKINVDCx16_ASAP7_75t_R g11 ( .A(n_7), .Y(n_11) );
NOR2xp33_ASAP7_75t_SL g7 ( .A(n_8), .B(n_9), .Y(n_7) );
INVx1_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
endmodule