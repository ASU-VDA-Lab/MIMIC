module real_aes_1226_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_824, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_822, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_823, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_824;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_822;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_823;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_746;
wire n_316;
wire n_284;
wire n_532;
wire n_656;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_725;
wire n_504;
wire n_455;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_358;
wire n_275;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_475;
wire n_554;
wire n_798;
wire n_668;
wire n_797;
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_0), .A2(n_199), .B1(n_482), .B2(n_513), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_1), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_2), .A2(n_245), .B1(n_596), .B2(n_801), .Y(n_800) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_3), .A2(n_197), .B1(n_489), .B2(n_490), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_4), .A2(n_11), .B1(n_539), .B2(n_707), .Y(n_706) );
OA22x2_ASAP7_75t_L g723 ( .A1(n_5), .A2(n_724), .B1(n_725), .B2(n_726), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_5), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_6), .B(n_341), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_7), .A2(n_213), .B1(n_741), .B2(n_742), .Y(n_740) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_8), .A2(n_198), .B1(n_296), .B2(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g753 ( .A(n_8), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_9), .A2(n_169), .B1(n_477), .B2(n_478), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_10), .A2(n_85), .B1(n_729), .B2(n_730), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_12), .A2(n_50), .B1(n_316), .B2(n_320), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_13), .A2(n_125), .B1(n_326), .B2(n_330), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_14), .A2(n_180), .B1(n_438), .B2(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_15), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_16), .A2(n_20), .B1(n_513), .B2(n_714), .Y(n_778) );
NAND2xp5_ASAP7_75t_SL g795 ( .A(n_17), .B(n_730), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_18), .A2(n_256), .B1(n_290), .B2(n_310), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_19), .A2(n_133), .B1(n_408), .B2(n_411), .Y(n_461) );
AOI22x1_ASAP7_75t_L g407 ( .A1(n_21), .A2(n_121), .B1(n_312), .B2(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_22), .A2(n_237), .B1(n_401), .B2(n_402), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_23), .A2(n_119), .B1(n_520), .B2(n_521), .Y(n_519) );
AO22x2_ASAP7_75t_L g295 ( .A1(n_24), .A2(n_68), .B1(n_296), .B2(n_297), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_24), .B(n_752), .Y(n_751) );
AO222x2_ASAP7_75t_L g565 ( .A1(n_25), .A2(n_67), .B1(n_219), .B2(n_384), .C1(n_394), .C2(n_397), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_26), .A2(n_127), .B1(n_347), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_27), .A2(n_220), .B1(n_401), .B2(n_402), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_28), .A2(n_760), .B1(n_783), .B2(n_784), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_28), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_29), .A2(n_250), .B1(n_410), .B2(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_30), .A2(n_268), .B1(n_518), .B2(n_551), .Y(n_782) );
XNOR2xp5_ASAP7_75t_L g378 ( .A(n_31), .B(n_379), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_32), .A2(n_226), .B1(n_430), .B2(n_480), .Y(n_514) );
AOI222xp33_ASAP7_75t_L g554 ( .A1(n_33), .A2(n_59), .B1(n_158), .B2(n_384), .C1(n_451), .C2(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_34), .A2(n_230), .B1(n_492), .B2(n_493), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_35), .A2(n_162), .B1(n_423), .B2(n_594), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_36), .A2(n_214), .B1(n_334), .B2(n_337), .Y(n_333) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_37), .A2(n_234), .B1(n_387), .B2(n_390), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_38), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_39), .A2(n_242), .B1(n_338), .B2(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_40), .A2(n_252), .B1(n_393), .B2(n_394), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_41), .A2(n_109), .B1(n_404), .B2(n_405), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_42), .B(n_496), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_43), .A2(n_163), .B1(n_405), .B2(n_576), .Y(n_582) );
OA22x2_ASAP7_75t_L g626 ( .A1(n_44), .A2(n_627), .B1(n_628), .B2(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_44), .Y(n_627) );
AOI222xp33_ASAP7_75t_L g418 ( .A1(n_45), .A2(n_142), .B1(n_269), .B2(n_419), .C1(n_420), .C2(n_421), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_46), .A2(n_184), .B1(n_394), .B2(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g794 ( .A(n_47), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g804 ( .A1(n_47), .A2(n_48), .B(n_729), .Y(n_804) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_47), .A2(n_807), .B1(n_812), .B2(n_824), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_48), .Y(n_813) );
AOI222xp33_ASAP7_75t_SL g810 ( .A1(n_49), .A2(n_56), .B1(n_171), .B2(n_341), .C1(n_347), .C2(n_349), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_51), .A2(n_247), .B1(n_330), .B2(n_809), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_52), .A2(n_130), .B1(n_437), .B2(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_SL g567 ( .A1(n_53), .A2(n_110), .B1(n_396), .B2(n_456), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_54), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_55), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_57), .A2(n_264), .B1(n_363), .B2(n_367), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_58), .A2(n_145), .B1(n_363), .B2(n_367), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_60), .A2(n_210), .B1(n_390), .B2(n_674), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_61), .A2(n_100), .B1(n_798), .B2(n_799), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_62), .A2(n_150), .B1(n_548), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_63), .A2(n_258), .B1(n_326), .B2(n_714), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_64), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_65), .A2(n_179), .B1(n_478), .B2(n_553), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_66), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_69), .A2(n_106), .B1(n_396), .B2(n_397), .Y(n_395) );
AOI22xp33_ASAP7_75t_SL g619 ( .A1(n_70), .A2(n_212), .B1(n_437), .B2(n_620), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_71), .A2(n_118), .B1(n_482), .B2(n_483), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_72), .A2(n_175), .B1(n_408), .B2(n_410), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_73), .A2(n_243), .B1(n_405), .B2(n_465), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g270 ( .A1(n_74), .A2(n_271), .B1(n_281), .B2(n_755), .C(n_758), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_75), .A2(n_141), .B1(n_441), .B2(n_443), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_76), .A2(n_194), .B1(n_443), .B2(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_77), .A2(n_123), .B1(n_396), .B2(n_454), .Y(n_453) );
OAI22x1_ASAP7_75t_L g534 ( .A1(n_78), .A2(n_535), .B1(n_556), .B2(n_557), .Y(n_534) );
CKINVDCx16_ASAP7_75t_R g557 ( .A(n_78), .Y(n_557) );
INVx1_ASAP7_75t_L g719 ( .A(n_79), .Y(n_719) );
INVx3_ASAP7_75t_L g296 ( .A(n_80), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_81), .A2(n_159), .B1(n_411), .B2(n_576), .Y(n_575) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_82), .A2(n_285), .B(n_372), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_82), .B(n_287), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_83), .A2(n_88), .B1(n_354), .B2(n_357), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_84), .A2(n_192), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_86), .A2(n_261), .B1(n_431), .B2(n_685), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_87), .A2(n_89), .B1(n_334), .B2(n_732), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_90), .A2(n_193), .B1(n_489), .B2(n_490), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_91), .A2(n_181), .B1(n_538), .B2(n_539), .Y(n_537) );
OA22x2_ASAP7_75t_L g472 ( .A1(n_92), .A2(n_473), .B1(n_474), .B2(n_497), .Y(n_472) );
INVxp67_ASAP7_75t_L g497 ( .A(n_92), .Y(n_497) );
OA22x2_ASAP7_75t_L g526 ( .A1(n_92), .A2(n_473), .B1(n_474), .B2(n_497), .Y(n_526) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_93), .A2(n_177), .B1(n_430), .B2(n_618), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_94), .A2(n_211), .B1(n_658), .B2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_95), .A2(n_236), .B1(n_347), .B2(n_493), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_96), .A2(n_126), .B1(n_326), .B2(n_620), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_97), .A2(n_200), .B1(n_317), .B2(n_480), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_98), .A2(n_251), .B1(n_423), .B2(n_424), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_99), .A2(n_182), .B1(n_402), .B2(n_460), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g643 ( .A(n_101), .Y(n_643) );
INVx1_ASAP7_75t_SL g305 ( .A(n_102), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_102), .B(n_134), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_103), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_104), .Y(n_385) );
INVx2_ASAP7_75t_L g280 ( .A(n_105), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_107), .A2(n_183), .B1(n_547), .B2(n_548), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_108), .A2(n_152), .B1(n_433), .B2(n_435), .Y(n_432) );
OA22x2_ASAP7_75t_L g499 ( .A1(n_111), .A2(n_500), .B1(n_523), .B2(n_524), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_111), .Y(n_523) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_112), .A2(n_120), .B1(n_427), .B2(n_490), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_113), .A2(n_147), .B1(n_354), .B2(n_357), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_114), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_115), .A2(n_195), .B1(n_437), .B2(n_482), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_116), .A2(n_143), .B1(n_426), .B2(n_427), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_117), .B(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_122), .A2(n_223), .B1(n_312), .B2(n_334), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_124), .A2(n_167), .B1(n_338), .B2(n_486), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_128), .A2(n_225), .B1(n_648), .B2(n_781), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_129), .A2(n_218), .B1(n_427), .B2(n_490), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_131), .A2(n_267), .B1(n_393), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_132), .A2(n_138), .B1(n_430), .B2(n_480), .Y(n_479) );
AO22x2_ASAP7_75t_L g308 ( .A1(n_134), .A2(n_207), .B1(n_296), .B2(n_309), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_135), .A2(n_260), .B1(n_424), .B2(n_596), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_136), .A2(n_231), .B1(n_687), .B2(n_688), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_137), .A2(n_140), .B1(n_435), .B2(n_477), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_139), .A2(n_206), .B1(n_411), .B2(n_584), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_144), .A2(n_165), .B1(n_489), .B2(n_490), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_146), .A2(n_257), .B1(n_594), .B2(n_596), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_148), .A2(n_224), .B1(n_363), .B2(n_539), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_149), .A2(n_161), .B1(n_437), .B2(n_438), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_151), .B(n_738), .Y(n_737) );
XNOR2x1_ASAP7_75t_L g579 ( .A(n_153), .B(n_580), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_154), .A2(n_217), .B1(n_420), .B2(n_421), .Y(n_509) );
INVx1_ASAP7_75t_L g306 ( .A(n_155), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_156), .A2(n_189), .B1(n_430), .B2(n_431), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_157), .A2(n_229), .B1(n_387), .B2(n_451), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_160), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_164), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_166), .A2(n_209), .B1(n_592), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_168), .A2(n_244), .B1(n_312), .B2(n_553), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_170), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_172), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_173), .A2(n_238), .B1(n_346), .B2(n_349), .Y(n_345) );
INVx1_ASAP7_75t_L g668 ( .A(n_174), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_176), .A2(n_188), .B1(n_423), .B2(n_424), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_178), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_185), .A2(n_204), .B1(n_424), .B2(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_186), .A2(n_190), .B1(n_443), .B2(n_517), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_187), .A2(n_262), .B1(n_317), .B2(n_480), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_191), .A2(n_239), .B1(n_349), .B2(n_592), .Y(n_591) );
CKINVDCx16_ASAP7_75t_R g466 ( .A(n_196), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_201), .A2(n_235), .B1(n_687), .B2(n_717), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_202), .A2(n_222), .B1(n_410), .B2(n_411), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_203), .A2(n_263), .B1(n_363), .B2(n_367), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_205), .A2(n_562), .B1(n_563), .B2(n_577), .Y(n_561) );
INVx1_ASAP7_75t_L g577 ( .A(n_205), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_208), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_215), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g749 ( .A(n_215), .Y(n_749) );
OA22x2_ASAP7_75t_L g413 ( .A1(n_216), .A2(n_414), .B1(n_415), .B2(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_216), .Y(n_414) );
INVx1_ASAP7_75t_L g602 ( .A(n_221), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_227), .A2(n_259), .B1(n_346), .B2(n_349), .Y(n_639) );
INVx1_ASAP7_75t_L g276 ( .A(n_228), .Y(n_276) );
AND2x2_ASAP7_75t_R g786 ( .A(n_228), .B(n_749), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_232), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_233), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_240), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_241), .Y(n_772) );
INVxp67_ASAP7_75t_L g278 ( .A(n_246), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_248), .A2(n_266), .B1(n_404), .B2(n_405), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_249), .B(n_384), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_253), .A2(n_265), .B1(n_354), .B2(n_703), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_254), .B(n_341), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_255), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_SL g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g820 ( .A(n_275), .B(n_277), .Y(n_820) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_276), .B(n_749), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AOI21xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_597), .B(n_746), .Y(n_281) );
INVx1_ASAP7_75t_L g756 ( .A(n_282), .Y(n_756) );
XOR2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_530), .Y(n_282) );
XNOR2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_373), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_339), .Y(n_287) );
NAND4xp25_ASAP7_75t_SL g288 ( .A(n_289), .B(n_315), .C(n_325), .D(n_333), .Y(n_288) );
INVx4_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_SL g430 ( .A(n_291), .Y(n_430) );
INVx2_ASAP7_75t_L g553 ( .A(n_291), .Y(n_553) );
INVx2_ASAP7_75t_SL g648 ( .A(n_291), .Y(n_648) );
INVx3_ASAP7_75t_SL g687 ( .A(n_291), .Y(n_687) );
INVx8_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_301), .Y(n_292) );
AND2x2_ASAP7_75t_L g318 ( .A(n_293), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g335 ( .A(n_293), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g343 ( .A(n_293), .B(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g384 ( .A(n_293), .B(n_344), .Y(n_384) );
AND2x2_ASAP7_75t_L g404 ( .A(n_293), .B(n_336), .Y(n_404) );
AND2x6_ASAP7_75t_L g408 ( .A(n_293), .B(n_319), .Y(n_408) );
AND2x2_ASAP7_75t_L g410 ( .A(n_293), .B(n_301), .Y(n_410) );
AND2x2_ASAP7_75t_L g576 ( .A(n_293), .B(n_336), .Y(n_576) );
AND2x4_ASAP7_75t_L g293 ( .A(n_294), .B(n_298), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g314 ( .A(n_295), .B(n_298), .Y(n_314) );
INVx1_ASAP7_75t_L g324 ( .A(n_295), .Y(n_324) );
AND2x2_ASAP7_75t_L g332 ( .A(n_295), .B(n_299), .Y(n_332) );
INVx2_ASAP7_75t_L g297 ( .A(n_296), .Y(n_297) );
INVx1_ASAP7_75t_L g300 ( .A(n_296), .Y(n_300) );
OAI22x1_ASAP7_75t_L g303 ( .A1(n_296), .A2(n_304), .B1(n_305), .B2(n_306), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_296), .Y(n_304) );
INVx1_ASAP7_75t_L g309 ( .A(n_296), .Y(n_309) );
INVxp67_ASAP7_75t_L g352 ( .A(n_298), .Y(n_352) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g323 ( .A(n_299), .B(n_324), .Y(n_323) );
AND2x4_ASAP7_75t_L g313 ( .A(n_301), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g322 ( .A(n_301), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g338 ( .A(n_301), .B(n_332), .Y(n_338) );
AND2x4_ASAP7_75t_L g405 ( .A(n_301), .B(n_332), .Y(n_405) );
AND2x6_ASAP7_75t_L g411 ( .A(n_301), .B(n_323), .Y(n_411) );
AND2x2_ASAP7_75t_L g465 ( .A(n_301), .B(n_314), .Y(n_465) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_307), .Y(n_301) );
AND2x2_ASAP7_75t_L g319 ( .A(n_302), .B(n_308), .Y(n_319) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g336 ( .A(n_303), .B(n_307), .Y(n_336) );
AND2x2_ASAP7_75t_L g344 ( .A(n_303), .B(n_308), .Y(n_344) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_303), .Y(n_361) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx2_ASAP7_75t_L g331 ( .A(n_308), .Y(n_331) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_311), .A2(n_442), .B1(n_642), .B2(n_643), .Y(n_641) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx3_ASAP7_75t_L g435 ( .A(n_313), .Y(n_435) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_313), .Y(n_478) );
INVx2_ASAP7_75t_L g522 ( .A(n_313), .Y(n_522) );
AND2x4_ASAP7_75t_L g348 ( .A(n_314), .B(n_319), .Y(n_348) );
AND2x2_ASAP7_75t_L g356 ( .A(n_314), .B(n_336), .Y(n_356) );
AND2x4_ASAP7_75t_L g387 ( .A(n_314), .B(n_336), .Y(n_387) );
AND2x2_ASAP7_75t_L g393 ( .A(n_314), .B(n_319), .Y(n_393) );
AND2x2_ASAP7_75t_L g456 ( .A(n_314), .B(n_319), .Y(n_456) );
BUFx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx3_ASAP7_75t_L g434 ( .A(n_318), .Y(n_434) );
BUFx2_ASAP7_75t_L g547 ( .A(n_318), .Y(n_547) );
AND2x2_ASAP7_75t_L g329 ( .A(n_319), .B(n_323), .Y(n_329) );
AND2x2_ASAP7_75t_SL g401 ( .A(n_319), .B(n_323), .Y(n_401) );
AND2x2_ASAP7_75t_L g460 ( .A(n_319), .B(n_323), .Y(n_460) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_SL g431 ( .A(n_321), .Y(n_431) );
INVx2_ASAP7_75t_L g480 ( .A(n_321), .Y(n_480) );
INVx2_ASAP7_75t_L g548 ( .A(n_321), .Y(n_548) );
INVx1_ASAP7_75t_SL g618 ( .A(n_321), .Y(n_618) );
INVx2_ASAP7_75t_L g658 ( .A(n_321), .Y(n_658) );
INVx8_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g366 ( .A(n_323), .B(n_336), .Y(n_366) );
AND2x4_ASAP7_75t_L g396 ( .A(n_323), .B(n_336), .Y(n_396) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_324), .Y(n_371) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g484 ( .A(n_328), .Y(n_484) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_329), .Y(n_437) );
BUFx3_ASAP7_75t_L g513 ( .A(n_329), .Y(n_513) );
INVx5_ASAP7_75t_SL g439 ( .A(n_330), .Y(n_439) );
BUFx2_ASAP7_75t_L g482 ( .A(n_330), .Y(n_482) );
BUFx2_ASAP7_75t_L g545 ( .A(n_330), .Y(n_545) );
BUFx3_ASAP7_75t_L g714 ( .A(n_330), .Y(n_714) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
AND2x4_ASAP7_75t_L g402 ( .A(n_331), .B(n_332), .Y(n_402) );
AND2x2_ASAP7_75t_L g360 ( .A(n_332), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_SL g390 ( .A(n_332), .B(n_361), .Y(n_390) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_332), .B(n_361), .Y(n_451) );
BUFx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx6_ASAP7_75t_L g442 ( .A(n_335), .Y(n_442) );
BUFx3_ASAP7_75t_L g551 ( .A(n_335), .Y(n_551) );
BUFx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g444 ( .A(n_338), .Y(n_444) );
BUFx3_ASAP7_75t_L g518 ( .A(n_338), .Y(n_518) );
BUFx2_ASAP7_75t_SL g651 ( .A(n_338), .Y(n_651) );
BUFx3_ASAP7_75t_L g688 ( .A(n_338), .Y(n_688) );
NAND4xp25_ASAP7_75t_SL g339 ( .A(n_340), .B(n_345), .C(n_353), .D(n_362), .Y(n_339) );
INVx3_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx4_ASAP7_75t_SL g419 ( .A(n_342), .Y(n_419) );
INVx3_ASAP7_75t_L g496 ( .A(n_342), .Y(n_496) );
INVx4_ASAP7_75t_SL g612 ( .A(n_342), .Y(n_612) );
INVx3_ASAP7_75t_SL g634 ( .A(n_342), .Y(n_634) );
INVx6_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g351 ( .A(n_344), .B(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g369 ( .A(n_344), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g394 ( .A(n_344), .B(n_352), .Y(n_394) );
AND2x2_ASAP7_75t_L g397 ( .A(n_344), .B(n_370), .Y(n_397) );
AND2x2_ASAP7_75t_L g454 ( .A(n_344), .B(n_370), .Y(n_454) );
AND2x2_ASAP7_75t_L g542 ( .A(n_344), .B(n_352), .Y(n_542) );
BUFx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_L g741 ( .A(n_347), .Y(n_741) );
INVx1_ASAP7_75t_L g773 ( .A(n_347), .Y(n_773) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx3_ASAP7_75t_L g421 ( .A(n_348), .Y(n_421) );
BUFx2_ASAP7_75t_L g492 ( .A(n_348), .Y(n_492) );
BUFx2_ASAP7_75t_L g592 ( .A(n_348), .Y(n_592) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_SL g420 ( .A(n_350), .Y(n_420) );
INVx1_ASAP7_75t_L g493 ( .A(n_350), .Y(n_493) );
INVx2_ASAP7_75t_L g678 ( .A(n_350), .Y(n_678) );
INVx2_ASAP7_75t_SL g709 ( .A(n_350), .Y(n_709) );
INVx2_ASAP7_75t_L g742 ( .A(n_350), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_350), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_771) );
INVx6_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx5_ASAP7_75t_L g424 ( .A(n_356), .Y(n_424) );
INVx2_ASAP7_75t_L g595 ( .A(n_356), .Y(n_595) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g423 ( .A(n_359), .Y(n_423) );
INVx2_ASAP7_75t_L g504 ( .A(n_359), .Y(n_504) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx12f_ASAP7_75t_L g596 ( .A(n_360), .Y(n_596) );
BUFx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g489 ( .A(n_365), .Y(n_489) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_366), .Y(n_427) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_366), .Y(n_538) );
BUFx6f_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx4f_ASAP7_75t_L g426 ( .A(n_369), .Y(n_426) );
BUFx6f_ASAP7_75t_SL g490 ( .A(n_369), .Y(n_490) );
INVx2_ASAP7_75t_L g540 ( .A(n_369), .Y(n_540) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
XNOR2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_468), .Y(n_373) );
OAI22x1_ASAP7_75t_SL g374 ( .A1(n_375), .A2(n_376), .B1(n_412), .B2(n_467), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2x1p5_ASAP7_75t_L g379 ( .A(n_380), .B(n_398), .Y(n_379) );
NOR2x1_ASAP7_75t_L g380 ( .A(n_381), .B(n_391), .Y(n_380) );
OAI222xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B1(n_385), .B2(n_386), .C1(n_388), .C2(n_389), .Y(n_381) );
OAI21xp5_ASAP7_75t_SL g671 ( .A1(n_383), .A2(n_672), .B(n_673), .Y(n_671) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g674 ( .A(n_386), .Y(n_674) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_387), .Y(n_555) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_395), .Y(n_391) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_406), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_403), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g585 ( .A(n_408), .Y(n_585) );
INVx2_ASAP7_75t_L g467 ( .A(n_412), .Y(n_467) );
XNOR2x1_ASAP7_75t_L g412 ( .A(n_413), .B(n_445), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_428), .Y(n_416) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_422), .C(n_425), .Y(n_417) );
INVx1_ASAP7_75t_L g768 ( .A(n_427), .Y(n_768) );
NAND4xp25_ASAP7_75t_L g428 ( .A(n_429), .B(n_432), .C(n_436), .D(n_440), .Y(n_428) );
BUFx2_ASAP7_75t_L g729 ( .A(n_430), .Y(n_729) );
INVx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g477 ( .A(n_434), .Y(n_477) );
INVx2_ASAP7_75t_L g520 ( .A(n_434), .Y(n_520) );
INVx3_ASAP7_75t_L g685 ( .A(n_434), .Y(n_685) );
BUFx2_ASAP7_75t_L g730 ( .A(n_435), .Y(n_730) );
INVx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g620 ( .A(n_439), .Y(n_620) );
OAI22xp33_ASAP7_75t_SL g660 ( .A1(n_439), .A2(n_661), .B1(n_664), .B2(n_665), .Y(n_660) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx3_ASAP7_75t_L g486 ( .A(n_442), .Y(n_486) );
INVx2_ASAP7_75t_L g517 ( .A(n_442), .Y(n_517) );
INVx1_ASAP7_75t_SL g798 ( .A(n_442), .Y(n_798) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_SL g732 ( .A(n_444), .Y(n_732) );
INVx2_ASAP7_75t_L g527 ( .A(n_445), .Y(n_527) );
INVx1_ASAP7_75t_L g529 ( .A(n_445), .Y(n_529) );
XOR2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_466), .Y(n_445) );
NAND2x1p5_ASAP7_75t_L g446 ( .A(n_447), .B(n_457), .Y(n_446) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_452), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_462), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
AOI22xp5_ASAP7_75t_SL g468 ( .A1(n_469), .A2(n_470), .B1(n_527), .B2(n_528), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_498), .B1(n_499), .B2(n_526), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_487), .Y(n_474) );
NAND4xp25_ASAP7_75t_SL g475 ( .A(n_476), .B(n_479), .C(n_481), .D(n_485), .Y(n_475) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_478), .Y(n_717) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g663 ( .A(n_484), .Y(n_663) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_484), .Y(n_809) );
NAND4xp25_ASAP7_75t_L g487 ( .A(n_488), .B(n_491), .C(n_494), .D(n_495), .Y(n_487) );
INVxp67_ASAP7_75t_L g770 ( .A(n_490), .Y(n_770) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
NOR3xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_506), .C(n_508), .Y(n_501) );
NOR4xp25_ASAP7_75t_L g524 ( .A(n_502), .B(n_511), .C(n_515), .D(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_505), .Y(n_502) );
INVxp67_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_507), .B(n_509), .Y(n_525) );
INVxp67_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_514), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .Y(n_515) );
BUFx2_ASAP7_75t_L g655 ( .A(n_520), .Y(n_655) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g781 ( .A(n_522), .Y(n_781) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AO22x2_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B1(n_558), .B2(n_559), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NAND4xp25_ASAP7_75t_SL g535 ( .A(n_536), .B(n_543), .C(n_549), .D(n_554), .Y(n_535) );
AND4x1_ASAP7_75t_L g556 ( .A(n_536), .B(n_543), .C(n_549), .D(n_554), .Y(n_556) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
BUFx6f_ASAP7_75t_SL g707 ( .A(n_538), .Y(n_707) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
INVx2_ASAP7_75t_L g793 ( .A(n_547), .Y(n_793) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OA22x2_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_578), .B2(n_579), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_564), .B(n_569), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
NOR2x1_ASAP7_75t_L g580 ( .A(n_581), .B(n_588), .Y(n_580) );
NAND4xp25_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .C(n_586), .D(n_587), .Y(n_581) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND4xp25_ASAP7_75t_SL g588 ( .A(n_589), .B(n_590), .C(n_591), .D(n_593), .Y(n_588) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_594), .Y(n_699) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g801 ( .A(n_595), .Y(n_801) );
BUFx3_ASAP7_75t_L g703 ( .A(n_596), .Y(n_703) );
INVx1_ASAP7_75t_L g757 ( .A(n_597), .Y(n_757) );
AOI22xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_721), .B1(n_722), .B2(n_745), .Y(n_597) );
INVx1_ASAP7_75t_L g745 ( .A(n_598), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_693), .B1(n_694), .B2(n_720), .Y(n_598) );
INVx1_ASAP7_75t_L g720 ( .A(n_599), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_625), .B1(n_691), .B2(n_692), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_601), .Y(n_691) );
OAI21x1_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B(n_624), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_602), .B(n_605), .Y(n_624) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_615), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_610), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .B(n_614), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_621), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g692 ( .A(n_625), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_666), .B1(n_689), .B2(n_690), .Y(n_625) );
INVx1_ASAP7_75t_SL g689 ( .A(n_626), .Y(n_689) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND3x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_640), .C(n_652), .Y(n_629) );
NOR2xp67_ASAP7_75t_SL g630 ( .A(n_631), .B(n_637), .Y(n_630) );
OAI21xp5_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_635), .B(n_636), .Y(n_631) );
OAI222xp33_ASAP7_75t_L g697 ( .A1(n_632), .A2(n_698), .B1(n_700), .B2(n_701), .C1(n_702), .C2(n_704), .Y(n_697) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g739 ( .A(n_634), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_638), .B(n_639), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_644), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_649), .B2(n_650), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_660), .Y(n_652) );
OAI22xp33_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_656), .B1(n_657), .B2(n_659), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g690 ( .A(n_666), .Y(n_690) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
XNOR2x1_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NAND2x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_679), .Y(n_669) );
NOR2xp67_ASAP7_75t_L g670 ( .A(n_671), .B(n_675), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_683), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
BUFx6f_ASAP7_75t_L g799 ( .A(n_688), .Y(n_799) );
INVx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
XOR2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_719), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_696), .B(n_710), .Y(n_695) );
NOR2x1_ASAP7_75t_L g696 ( .A(n_697), .B(n_705), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_715), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NOR3x1_ASAP7_75t_SL g726 ( .A(n_727), .B(n_733), .C(n_736), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_731), .Y(n_727) );
INVx1_ASAP7_75t_L g814 ( .A(n_729), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
NAND4xp25_ASAP7_75t_SL g736 ( .A(n_737), .B(n_740), .C(n_743), .D(n_744), .Y(n_736) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_750), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_748), .B(n_751), .Y(n_817) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
OAI222xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_785), .B1(n_787), .B2(n_794), .C1(n_815), .C2(n_818), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_760), .Y(n_784) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_775), .Y(n_761) );
NOR3xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_766), .C(n_771), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B1(n_769), .B2(n_770), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_779), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_782), .Y(n_779) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OR2x2_ASAP7_75t_L g787 ( .A(n_788), .B(n_802), .Y(n_787) );
OAI222xp33_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_794), .B1(n_795), .B2(n_796), .C1(n_822), .C2(n_823), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_789), .B(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g803 ( .A(n_795), .B(n_796), .C(n_804), .Y(n_803) );
AND2x2_ASAP7_75t_SL g796 ( .A(n_797), .B(n_800), .Y(n_796) );
OAI21xp5_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_805), .B(n_811), .Y(n_802) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_810), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
CKINVDCx6p67_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
endmodule