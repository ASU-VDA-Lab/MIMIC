module fake_jpeg_11226_n_193 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_193);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_42),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_31),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_16),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_9),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_90),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_89),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_81),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_100),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_65),
.B(n_80),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_99),
.C(n_103),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_63),
.B1(n_55),
.B2(n_71),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g101 ( 
.A(n_82),
.Y(n_101)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_81),
.B1(n_57),
.B2(n_63),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_106),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_84),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_98),
.A2(n_81),
.B1(n_57),
.B2(n_55),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_119),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

OR2x2_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_75),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_5),
.Y(n_151)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_78),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_122),
.Y(n_138)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_64),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_123),
.B(n_124),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_69),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_76),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_77),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_61),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_115),
.C(n_128),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_151),
.C(n_134),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_117),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_141),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_122),
.A2(n_71),
.B1(n_60),
.B2(n_59),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_145),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_73),
.B1(n_70),
.B2(n_72),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_66),
.B1(n_65),
.B2(n_79),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_54),
.Y(n_141)
);

AOI32xp33_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_54),
.B1(n_3),
.B2(n_4),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_113),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_148),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_2),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_149),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_151),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_162)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_156),
.B(n_159),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_158),
.C(n_160),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_166),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_133),
.B1(n_140),
.B2(n_132),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_50),
.B(n_14),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_35),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_147),
.A3(n_19),
.B1(n_22),
.B2(n_23),
.C1(n_27),
.C2(n_28),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_150),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_12),
.B(n_30),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_155),
.C(n_153),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_175),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_40),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_177),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_34),
.B(n_37),
.C(n_39),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_154),
.B1(n_166),
.B2(n_167),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_179),
.A2(n_170),
.B1(n_166),
.B2(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_182),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_179),
.C(n_180),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_173),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_185),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_185),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_183),
.B(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_191),
.B(n_181),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_176),
.Y(n_193)
);


endmodule