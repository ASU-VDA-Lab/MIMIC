module fake_jpeg_27508_n_117 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_117);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_4),
.B(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

OR2x2_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_54),
.Y(n_64)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_1),
.Y(n_54)
);

CKINVDCx12_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_2),
.Y(n_57)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_43),
.B1(n_46),
.B2(n_50),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_62),
.B1(n_69),
.B2(n_7),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_46),
.B1(n_49),
.B2(n_41),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_68),
.B1(n_2),
.B2(n_5),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_43),
.B1(n_40),
.B2(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_44),
.B1(n_3),
.B2(n_4),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_44),
.B1(n_5),
.B2(n_7),
.Y(n_69)
);

O2A1O1Ixp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_21),
.B(n_36),
.C(n_35),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_82),
.Y(n_88)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_77),
.B1(n_58),
.B2(n_9),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_23),
.B(n_34),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_78),
.B(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_78),
.Y(n_87)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_8),
.Y(n_78)
);

AND2x6_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_18),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_8),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g83 ( 
.A(n_66),
.Y(n_83)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_9),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_13),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_81),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_93),
.B1(n_95),
.B2(n_25),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_96),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_14),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_74),
.B1(n_86),
.B2(n_71),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_98),
.B(n_104),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_101),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_16),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_103),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_17),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_95),
.B1(n_90),
.B2(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_100),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_110),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_103),
.B(n_92),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_105),
.B(n_106),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_112),
.B(n_107),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_26),
.B(n_27),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_114),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_90),
.B(n_29),
.C(n_30),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_28),
.Y(n_117)
);


endmodule