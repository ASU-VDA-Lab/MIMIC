module real_jpeg_24706_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_215;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_167;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_182;
wire n_273;
wire n_253;
wire n_269;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_1),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_1),
.A2(n_22),
.B1(n_24),
.B2(n_31),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_1),
.A2(n_31),
.B1(n_53),
.B2(n_54),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_1),
.A2(n_31),
.B1(n_67),
.B2(n_68),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_5),
.A2(n_18),
.B1(n_27),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_5),
.A2(n_22),
.B1(n_24),
.B2(n_33),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_5),
.A2(n_33),
.B1(n_53),
.B2(n_54),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_5),
.A2(n_33),
.B1(n_67),
.B2(n_68),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_6),
.A2(n_18),
.B1(n_20),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_22),
.B1(n_24),
.B2(n_45),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_6),
.A2(n_45),
.B1(n_53),
.B2(n_54),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_6),
.A2(n_45),
.B1(n_67),
.B2(n_68),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_6),
.B(n_17),
.C(n_22),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_6),
.B(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_6),
.B(n_52),
.C(n_54),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_6),
.B(n_65),
.C(n_68),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_6),
.B(n_58),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_6),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_6),
.B(n_123),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_38),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_37),
.Y(n_12)
);

OR2x2_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_34),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_14),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_14),
.B(n_40),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_21),
.B1(n_25),
.B2(n_32),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_21),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_15),
.A2(n_21),
.B1(n_25),
.B2(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_21),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_16)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

OA22x2_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_21)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_18),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_21),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_22),
.A2(n_24),
.B1(n_52),
.B2(n_56),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_22),
.B(n_195),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_44),
.Y(n_43)
);

AO21x1_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_77),
.B(n_273),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_73),
.C(n_75),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_42),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.C(n_60),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_43),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_43),
.A2(n_86),
.B1(n_102),
.B2(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_43),
.B(n_119),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_43),
.A2(n_86),
.B1(n_118),
.B2(n_119),
.Y(n_141)
);

AOI211xp5_ASAP7_75t_L g163 ( 
.A1(n_43),
.A2(n_132),
.B(n_135),
.C(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_43),
.A2(n_86),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_43),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_43),
.A2(n_86),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_43),
.A2(n_100),
.B(n_103),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_44),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_47),
.B1(n_60),
.B2(n_61),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_58),
.B2(n_59),
.Y(n_47)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_51),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_50),
.A2(n_51),
.B1(n_90),
.B2(n_92),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_51)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_71)
);

INVx5_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_54),
.B(n_206),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_60),
.A2(n_61),
.B1(n_89),
.B2(n_261),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_86),
.C(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_72),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_63),
.B(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_64),
.A2(n_70),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_68),
.B(n_216),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_75),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_74),
.B(n_91),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_93),
.B(n_272),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_79),
.B(n_82),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.C(n_88),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_118),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_88),
.B(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_89),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI31xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_253),
.A3(n_264),
.B(n_269),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_154),
.B(n_252),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_137),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_96),
.B(n_137),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_126),
.B1(n_127),
.B2(n_136),
.Y(n_96)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_116),
.B2(n_117),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_99),
.B(n_116),
.C(n_126),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_114),
.B2(n_115),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_110),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_103),
.B1(n_110),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_107),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_106),
.B(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_107),
.A2(n_130),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_109),
.Y(n_217)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_120),
.B(n_125),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_118),
.B(n_120),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_162),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_118),
.A2(n_119),
.B1(n_132),
.B2(n_162),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_118),
.A2(n_119),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_119),
.B(n_167),
.C(n_182),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_119),
.A2(n_132),
.B(n_164),
.C(n_227),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_125),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_125),
.A2(n_258),
.B1(n_262),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_133),
.B(n_134),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_129),
.A2(n_132),
.B1(n_162),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_129),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_148),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_132),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_132),
.B(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_132),
.A2(n_162),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_132),
.A2(n_162),
.B1(n_204),
.B2(n_205),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_132),
.A2(n_162),
.B1(n_192),
.B2(n_233),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_133),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_133),
.A2(n_134),
.B(n_166),
.Y(n_244)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_146),
.B(n_153),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.C(n_145),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_138),
.A2(n_139),
.B1(n_143),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_141),
.B1(n_166),
.B2(n_173),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_140),
.A2(n_141),
.B1(n_146),
.B2(n_147),
.Y(n_241)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_143),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_145),
.B(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_246),
.B(n_251),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_185),
.B(n_237),
.C(n_245),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_175),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_157),
.B(n_175),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_165),
.B2(n_174),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_160),
.B(n_163),
.C(n_174),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_189),
.C(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_162),
.B(n_168),
.C(n_211),
.Y(n_224)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_166),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_168),
.B1(n_182),
.B2(n_183),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_167),
.A2(n_168),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_167),
.B(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_167),
.A2(n_168),
.B1(n_193),
.B2(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_168),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_168),
.B(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.C(n_180),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_177),
.A2(n_178),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_198),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_179),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_236),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_199),
.B(n_235),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_196),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_188),
.B(n_196),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_229),
.B(n_234),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_223),
.B(n_228),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_212),
.B(n_222),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_203),
.B(n_207),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_220),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_224),
.B(n_225),
.Y(n_228)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_230),
.B(n_231),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_239),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_242),
.C(n_244),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_250),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_257),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.C(n_263),
.Y(n_257)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_266),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_268),
.Y(n_270)
);


endmodule