module real_jpeg_32684_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_11;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_150;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_0),
.Y(n_138)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_1),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_2),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_2),
.Y(n_171)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_4),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_4),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_5),
.A2(n_78),
.B1(n_81),
.B2(n_82),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_5),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_5),
.A2(n_81),
.B1(n_126),
.B2(n_130),
.Y(n_125)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_6),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_6),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_34),
.B1(n_39),
.B2(n_45),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_7),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_8),
.A2(n_23),
.B1(n_26),
.B2(n_30),
.Y(n_22)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_8),
.A2(n_30),
.B1(n_174),
.B2(n_177),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_151),
.Y(n_9)
);

HB1xp67_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

AOI21x1_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_115),
.B(n_150),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_46),
.Y(n_12)
);

NOR2xp67_ASAP7_75t_L g150 ( 
.A(n_13),
.B(n_46),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_21),
.B1(n_31),
.B2(n_32),
.Y(n_13)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_14),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_14),
.B(n_125),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_18),
.Y(n_14)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_15),
.Y(n_31)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_17),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_17),
.Y(n_147)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_20),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp33_ASAP7_75t_SL g145 ( 
.A1(n_22),
.A2(n_146),
.B(n_148),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_25),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVxp33_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_33),
.A2(n_118),
.B(n_119),
.Y(n_156)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22x1_ASAP7_75t_L g85 ( 
.A1(n_37),
.A2(n_86),
.B1(n_89),
.B2(n_92),
.Y(n_85)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_44),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_75),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_47),
.B(n_75),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_54),
.B1(n_64),
.B2(n_70),
.Y(n_47)
);

INVxp67_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_49),
.A2(n_50),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_50),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_50),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_50),
.B(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_53),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_71),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_94),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_84),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_77),
.B(n_102),
.Y(n_181)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_84),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_102),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_110),
.B2(n_113),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_142),
.B(n_149),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_132),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_139),
.Y(n_132)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_143),
.B(n_145),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_173),
.B(n_181),
.Y(n_172)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_182),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NOR2xp67_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_155),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_172),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_164),
.B1(n_167),
.B2(n_169),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx5_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);


endmodule