module fake_jpeg_2466_n_525 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_525);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_52),
.Y(n_117)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_67),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_20),
.B(n_10),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_54),
.B(n_76),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_59),
.Y(n_144)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_63),
.Y(n_161)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_29),
.B(n_10),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_69),
.Y(n_153)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_74),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_84),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_18),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_34),
.B(n_10),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_25),
.B(n_10),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_90),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_87),
.B(n_88),
.Y(n_156)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_25),
.B(n_11),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_11),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_93),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_28),
.B(n_32),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_38),
.A2(n_9),
.B1(n_17),
.B2(n_2),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_94),
.A2(n_30),
.B1(n_32),
.B2(n_37),
.Y(n_139)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_97),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_99),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_39),
.CON(n_133),
.SN(n_133)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_28),
.B(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_102),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_98),
.A2(n_43),
.B1(n_44),
.B2(n_41),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_104),
.A2(n_139),
.B1(n_141),
.B2(n_146),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_26),
.B1(n_36),
.B2(n_43),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_97),
.B1(n_96),
.B2(n_59),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_110),
.A2(n_42),
.B1(n_21),
.B2(n_1),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_26),
.B1(n_36),
.B2(n_43),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_113),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_52),
.A2(n_50),
.B(n_30),
.C(n_45),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_115),
.B(n_63),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_62),
.A2(n_36),
.B1(n_46),
.B2(n_40),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_68),
.A2(n_36),
.B1(n_46),
.B2(n_40),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_125),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_64),
.B(n_50),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_132),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_45),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_133),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_55),
.B(n_27),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_86),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_80),
.B(n_37),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_145),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_66),
.A2(n_36),
.B1(n_27),
.B2(n_41),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_56),
.B(n_23),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_58),
.A2(n_89),
.B1(n_77),
.B2(n_73),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_69),
.A2(n_41),
.B1(n_44),
.B2(n_39),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_155),
.B1(n_23),
.B2(n_78),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_69),
.A2(n_44),
.B1(n_39),
.B2(n_42),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_162),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_156),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_163),
.B(n_166),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g262 ( 
.A(n_164),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_165),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_61),
.C(n_81),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_172),
.B(n_150),
.C(n_112),
.Y(n_239)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_203),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_178),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_0),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_180),
.B(n_184),
.Y(n_240)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_117),
.Y(n_181)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_182),
.B(n_191),
.Y(n_231)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_121),
.B(n_0),
.Y(n_184)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_185),
.Y(n_247)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_189),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_109),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_193),
.A2(n_215),
.B1(n_128),
.B2(n_142),
.Y(n_257)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_194),
.Y(n_261)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_121),
.B(n_0),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_197),
.B(n_205),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_103),
.B(n_78),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_198),
.B(n_199),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_118),
.B(n_23),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_200),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_202),
.Y(n_267)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_126),
.B(n_71),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_133),
.B(n_153),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_0),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_139),
.A2(n_57),
.B1(n_42),
.B2(n_21),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_206),
.A2(n_207),
.B1(n_218),
.B2(n_123),
.Y(n_238)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_210),
.Y(n_228)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_209),
.Y(n_255)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_136),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_214),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_108),
.B(n_12),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_213),
.B(n_219),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_153),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_157),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_216),
.B(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_146),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_150),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_104),
.B1(n_126),
.B2(n_115),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_225),
.A2(n_232),
.B1(n_241),
.B2(n_236),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_173),
.A2(n_112),
.B1(n_135),
.B2(n_120),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_236),
.B(n_242),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_238),
.B(n_14),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_239),
.B(n_259),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_173),
.A2(n_120),
.B1(n_135),
.B2(n_130),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_175),
.A2(n_108),
.A3(n_152),
.B1(n_147),
.B2(n_154),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_179),
.A2(n_107),
.B1(n_149),
.B2(n_158),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_243),
.A2(n_244),
.B1(n_42),
.B2(n_209),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_179),
.A2(n_212),
.B1(n_176),
.B2(n_177),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_177),
.A2(n_158),
.B1(n_144),
.B2(n_130),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_246),
.A2(n_253),
.B1(n_167),
.B2(n_162),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_207),
.A2(n_136),
.B1(n_147),
.B2(n_142),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_215),
.B1(n_214),
.B2(n_164),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_180),
.A2(n_116),
.B1(n_106),
.B2(n_152),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_SL g281 ( 
.A1(n_257),
.A2(n_192),
.B(n_183),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_SL g258 ( 
.A(n_205),
.B(n_111),
.C(n_128),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_258),
.B(n_170),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_184),
.B(n_154),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_197),
.B(n_138),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_269),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_186),
.B(n_149),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_204),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_271),
.B(n_277),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_220),
.A2(n_212),
.B(n_176),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_272),
.A2(n_310),
.B(n_235),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_273),
.A2(n_280),
.B1(n_293),
.B2(n_303),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_274),
.A2(n_314),
.B1(n_235),
.B2(n_254),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_275),
.B(n_276),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_236),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_240),
.B(n_172),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_225),
.A2(n_204),
.B1(n_116),
.B2(n_106),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_278),
.A2(n_297),
.B1(n_298),
.B2(n_308),
.Y(n_316)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_281),
.A2(n_260),
.B1(n_268),
.B2(n_249),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_229),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_282),
.B(n_283),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_221),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_204),
.C(n_202),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g345 ( 
.A(n_284),
.B(n_288),
.C(n_305),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_285),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_239),
.A2(n_210),
.B(n_194),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_286),
.A2(n_255),
.B(n_226),
.Y(n_329)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_168),
.C(n_216),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_231),
.B(n_211),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_291),
.B(n_261),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_252),
.B(n_200),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_296),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_227),
.A2(n_203),
.B1(n_195),
.B2(n_171),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_241),
.B(n_187),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_294),
.Y(n_335)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_237),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_222),
.A2(n_185),
.B1(n_189),
.B2(n_178),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_228),
.Y(n_299)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_299),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_248),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_306),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_232),
.B(n_188),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_301),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_266),
.B(n_111),
.C(n_2),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_269),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_222),
.A2(n_18),
.B1(n_3),
.B2(n_4),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_307),
.A2(n_313),
.B1(n_263),
.B2(n_264),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_222),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_256),
.B(n_4),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_312),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_223),
.A2(n_6),
.B(n_8),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_242),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_267),
.B1(n_265),
.B2(n_224),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_256),
.B(n_233),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_253),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_315),
.B(n_337),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_276),
.A2(n_272),
.B(n_289),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_319),
.A2(n_329),
.B(n_330),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_223),
.C(n_234),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_336),
.C(n_355),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_304),
.B(n_258),
.Y(n_327)
);

XNOR2x1_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_350),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_289),
.A2(n_255),
.B1(n_247),
.B2(n_234),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_328),
.A2(n_341),
.B1(n_297),
.B2(n_301),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_289),
.A2(n_267),
.B(n_233),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_333),
.B(n_294),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_278),
.A2(n_247),
.B1(n_224),
.B2(n_264),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_334),
.A2(n_290),
.B1(n_296),
.B2(n_283),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_277),
.B(n_230),
.C(n_254),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_312),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_273),
.B(n_261),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_338),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_340),
.B(n_301),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_306),
.A2(n_265),
.B1(n_226),
.B2(n_230),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_343),
.Y(n_371)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_287),
.Y(n_344)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_344),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_346),
.A2(n_352),
.B(n_353),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_270),
.B(n_249),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_310),
.A2(n_250),
.B(n_15),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_286),
.A2(n_250),
.B(n_15),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_354),
.A2(n_307),
.B(n_294),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_288),
.B(n_14),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_338),
.A2(n_270),
.B1(n_298),
.B2(n_271),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_356),
.A2(n_362),
.B1(n_368),
.B2(n_383),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_288),
.C(n_284),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_372),
.C(n_385),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_317),
.B(n_292),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_359),
.B(n_364),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_348),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_363),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_338),
.A2(n_300),
.B1(n_314),
.B2(n_282),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_348),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_317),
.B(n_323),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_323),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_369),
.B(n_373),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_370),
.A2(n_328),
.B1(n_347),
.B2(n_335),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_284),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_337),
.B(n_291),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_331),
.B(n_299),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_377),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_331),
.B(n_309),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_378),
.Y(n_404)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_322),
.Y(n_379)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_379),
.Y(n_392)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_322),
.Y(n_380)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_380),
.Y(n_403)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_382),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_316),
.A2(n_318),
.B1(n_330),
.B2(n_319),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_340),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_384),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_336),
.B(n_345),
.C(n_350),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_386),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_318),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_387),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_316),
.A2(n_314),
.B1(n_313),
.B2(n_305),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_388),
.A2(n_308),
.B1(n_274),
.B2(n_326),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_389),
.A2(n_346),
.B(n_353),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_321),
.B(n_305),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_390),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_327),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_391),
.B(n_400),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_365),
.A2(n_351),
.B1(n_321),
.B2(n_349),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_395),
.A2(n_405),
.B1(n_413),
.B2(n_414),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_357),
.B(n_345),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_355),
.C(n_329),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_409),
.C(n_410),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_365),
.A2(n_334),
.B1(n_333),
.B2(n_347),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_406),
.A2(n_417),
.B1(n_419),
.B2(n_369),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_358),
.B(n_372),
.C(n_366),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_366),
.B(n_332),
.C(n_354),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_411),
.A2(n_367),
.B(n_381),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_364),
.B(n_332),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_412),
.B(n_416),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_383),
.A2(n_342),
.B1(n_344),
.B2(n_324),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_361),
.A2(n_342),
.B1(n_324),
.B2(n_325),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_359),
.B(n_325),
.C(n_326),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_362),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_390),
.B(n_341),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_361),
.A2(n_281),
.B1(n_315),
.B2(n_311),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_376),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_426),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_422),
.A2(n_428),
.B1(n_430),
.B2(n_440),
.Y(n_448)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_418),
.Y(n_423)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_423),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_384),
.Y(n_425)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_425),
.Y(n_458)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_394),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_408),
.A2(n_360),
.B1(n_363),
.B2(n_375),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_394),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_431),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_408),
.A2(n_368),
.B1(n_382),
.B2(n_373),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_398),
.B(n_374),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_433),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_402),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_436),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_407),
.B(n_377),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_367),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_445),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_414),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_442),
.Y(n_465)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_392),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_419),
.A2(n_356),
.B1(n_374),
.B2(n_353),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_441),
.A2(n_443),
.B1(n_417),
.B2(n_406),
.Y(n_454)
);

NOR3xp33_ASAP7_75t_SL g442 ( 
.A(n_392),
.B(n_381),
.C(n_386),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_420),
.A2(n_388),
.B1(n_370),
.B2(n_380),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_403),
.Y(n_444)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_444),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_399),
.B(n_415),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_396),
.C(n_409),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_447),
.C(n_453),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_396),
.C(n_401),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_391),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_456),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_399),
.C(n_412),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_454),
.A2(n_430),
.B1(n_443),
.B2(n_424),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_437),
.B(n_410),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_427),
.B(n_413),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_459),
.B(n_461),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_416),
.C(n_407),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_462),
.C(n_432),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_439),
.B(n_411),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_395),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_428),
.B(n_397),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_397),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_467),
.A2(n_476),
.B1(n_479),
.B2(n_480),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_469),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_449),
.A2(n_423),
.B1(n_426),
.B2(n_429),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_466),
.Y(n_471)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_471),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_465),
.A2(n_424),
.B1(n_425),
.B2(n_393),
.Y(n_472)
);

INVxp33_ASAP7_75t_L g493 ( 
.A(n_472),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_295),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_474),
.B(n_463),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_481),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_448),
.A2(n_442),
.B1(n_393),
.B2(n_440),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_405),
.Y(n_477)
);

XNOR2x1_ASAP7_75t_L g489 ( 
.A(n_477),
.B(n_450),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_457),
.A2(n_444),
.B1(n_403),
.B2(n_371),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_452),
.A2(n_379),
.B1(n_371),
.B2(n_389),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_455),
.A2(n_339),
.B1(n_302),
.B2(n_17),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_455),
.Y(n_482)
);

AOI21x1_ASAP7_75t_L g492 ( 
.A1(n_482),
.A2(n_461),
.B(n_302),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_480),
.A2(n_459),
.B(n_447),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_484),
.B(n_490),
.Y(n_506)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_485),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_446),
.C(n_451),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_SL g501 ( 
.A(n_487),
.B(n_488),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_477),
.A2(n_450),
.B(n_462),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_491),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_453),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_473),
.B(n_339),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_492),
.A2(n_482),
.B1(n_477),
.B2(n_479),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_456),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_470),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_496),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_467),
.C(n_478),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_500),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_478),
.C(n_470),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_493),
.A2(n_496),
.B1(n_483),
.B2(n_488),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_503),
.B(n_505),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_504),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_493),
.A2(n_481),
.B(n_16),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_510),
.B(n_511),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_501),
.A2(n_494),
.B(n_490),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_495),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_512),
.B(n_513),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_486),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_509),
.B(n_498),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_514),
.C(n_506),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_507),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_517),
.A2(n_507),
.B(n_502),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_518),
.B(n_515),
.C(n_516),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_519),
.A2(n_497),
.B(n_505),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_520),
.B(n_521),
.C(n_500),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_489),
.C(n_16),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_14),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_17),
.B(n_517),
.Y(n_525)
);


endmodule