module fake_jpeg_11268_n_191 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_191);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_29),
.B(n_9),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx11_ASAP7_75t_SL g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_27),
.Y(n_76)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_10),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_88),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_1),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_91),
.Y(n_102)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_2),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_85),
.A2(n_78),
.B1(n_58),
.B2(n_65),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_97),
.B1(n_61),
.B2(n_56),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_80),
.B(n_64),
.C(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_103),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_78),
.B1(n_54),
.B2(n_58),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_101),
.B1(n_71),
.B2(n_57),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_90),
.A2(n_79),
.B1(n_61),
.B2(n_57),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_60),
.B(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_2),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_79),
.B1(n_71),
.B2(n_56),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_76),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_112),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_99),
.Y(n_109)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_55),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_119),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_120),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_126),
.Y(n_132)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_75),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_97),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_122),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_123),
.A2(n_74),
.B(n_5),
.Y(n_137)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_63),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_3),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_73),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_11),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_3),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_148),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_145),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_77),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_139),
.A2(n_15),
.B(n_17),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_77),
.B1(n_25),
.B2(n_28),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_21),
.B(n_50),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_150),
.B(n_43),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_6),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_35),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_8),
.B(n_11),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_116),
.B1(n_110),
.B2(n_109),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_155),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_142),
.B1(n_129),
.B2(n_139),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_122),
.B1(n_13),
.B2(n_12),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_168),
.B(n_147),
.C(n_45),
.D(n_47),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_161)
);

XOR2x2_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_140),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_163),
.C(n_164),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_18),
.B1(n_19),
.B2(n_33),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_167),
.C(n_145),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_34),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_36),
.B(n_40),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_171),
.C(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

INVxp33_ASAP7_75t_SL g178 ( 
.A(n_176),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_181),
.C(n_182),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_157),
.C(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_180),
.B(n_172),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_154),
.B(n_166),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_172),
.B(n_178),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_183),
.B1(n_179),
.B2(n_164),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_175),
.B1(n_174),
.B2(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_187),
.B(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_189),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_146),
.Y(n_191)
);


endmodule