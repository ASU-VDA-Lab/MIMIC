module fake_jpeg_7307_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_38),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_51),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_22),
.B1(n_33),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_60),
.B1(n_63),
.B2(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_22),
.B1(n_33),
.B2(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_31),
.B1(n_26),
.B2(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_69),
.A2(n_93),
.B1(n_18),
.B2(n_20),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_70),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_126)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_73),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_56),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_22),
.B1(n_36),
.B2(n_35),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_90),
.B1(n_97),
.B2(n_23),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_40),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_79),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_28),
.B1(n_26),
.B2(n_32),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_77),
.A2(n_86),
.B1(n_100),
.B2(n_20),
.Y(n_130)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_40),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

FAx1_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_35),
.CI(n_37),
.CON(n_82),
.SN(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_28),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_94),
.C(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_26),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_29),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_59),
.A2(n_32),
.B1(n_41),
.B2(n_17),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_95),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_44),
.B1(n_42),
.B2(n_16),
.Y(n_90)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_0),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_54),
.A2(n_34),
.B1(n_30),
.B2(n_23),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_34),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_30),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_54),
.A2(n_17),
.B1(n_34),
.B2(n_30),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_24),
.A3(n_18),
.B1(n_20),
.B2(n_16),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_18),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_0),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_72),
.B1(n_78),
.B2(n_69),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_106),
.Y(n_136)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_110),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_12),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_68),
.B1(n_67),
.B2(n_23),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_91),
.B1(n_96),
.B2(n_75),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_71),
.B(n_11),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_117),
.B(n_0),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_44),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_129),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_126),
.B1(n_130),
.B2(n_96),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_71),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_13),
.B1(n_24),
.B2(n_2),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_44),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_92),
.C(n_102),
.Y(n_132)
);

AO22x1_ASAP7_75t_L g128 ( 
.A1(n_84),
.A2(n_42),
.B1(n_29),
.B2(n_27),
.Y(n_128)
);

AO22x1_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_82),
.B1(n_25),
.B2(n_29),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_73),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_147),
.C(n_160),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_138),
.A2(n_145),
.B1(n_150),
.B2(n_158),
.Y(n_195)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_139),
.B(n_144),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_141),
.B1(n_162),
.B2(n_104),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_94),
.B(n_84),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_148),
.B(n_154),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_94),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_75),
.B(n_81),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_103),
.A2(n_87),
.B1(n_82),
.B2(n_88),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_157),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_80),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_156),
.Y(n_173)
);

AO22x1_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_131),
.B1(n_21),
.B2(n_105),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_29),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_116),
.A2(n_27),
.B1(n_21),
.B2(n_13),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_27),
.C(n_21),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_114),
.A2(n_27),
.B1(n_21),
.B2(n_3),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_105),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_174),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_107),
.B1(n_128),
.B2(n_110),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_166),
.A2(n_171),
.B(n_179),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_128),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_169),
.C(n_184),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_117),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_21),
.B(n_120),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_175),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_155),
.A2(n_131),
.B1(n_104),
.B2(n_113),
.Y(n_176)
);

OAI22x1_ASAP7_75t_L g223 ( 
.A1(n_176),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_154),
.B1(n_162),
.B2(n_134),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_1),
.Y(n_178)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

XOR2x1_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_21),
.Y(n_179)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_180),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_1),
.Y(n_181)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_136),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_182),
.B(n_185),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_113),
.C(n_2),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_188),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_113),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_192),
.B(n_4),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_1),
.Y(n_189)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_191),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_134),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_142),
.A2(n_1),
.B(n_2),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_3),
.Y(n_193)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_4),
.C(n_5),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_159),
.C(n_151),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_170),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_207),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_220),
.C(n_224),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_152),
.B1(n_163),
.B2(n_135),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_205),
.B1(n_210),
.B2(n_217),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_139),
.B1(n_145),
.B2(n_133),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_170),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_209),
.A2(n_194),
.B1(n_181),
.B2(n_189),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_198),
.A2(n_149),
.B1(n_5),
.B2(n_6),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_149),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_213),
.B(n_169),
.Y(n_241)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_193),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_198),
.A2(n_186),
.B1(n_187),
.B2(n_166),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_219),
.A2(n_183),
.B1(n_192),
.B2(n_178),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_167),
.B(n_7),
.C(n_8),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_223),
.A2(n_180),
.B1(n_191),
.B2(n_171),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_167),
.B(n_10),
.C(n_168),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_225),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_165),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_184),
.C(n_165),
.Y(n_244)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_230),
.A2(n_251),
.B1(n_252),
.B2(n_210),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_172),
.B(n_182),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_238),
.B1(n_248),
.B2(n_249),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_195),
.B1(n_164),
.B2(n_174),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_240),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_227),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_216),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_253),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_196),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_211),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_219),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_205),
.A2(n_164),
.B1(n_174),
.B2(n_185),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_214),
.Y(n_255)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_173),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_263),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_224),
.C(n_199),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_266),
.C(n_267),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_262),
.B1(n_274),
.B2(n_249),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_204),
.B1(n_222),
.B2(n_206),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_232),
.B(n_226),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_238),
.B(n_226),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_263),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_199),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_220),
.C(n_173),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_229),
.Y(n_271)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_202),
.C(n_201),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_231),
.C(n_233),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_230),
.A2(n_206),
.B1(n_200),
.B2(n_207),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_246),
.B(n_248),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_276),
.A2(n_286),
.B(n_290),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_242),
.B1(n_233),
.B2(n_250),
.Y(n_277)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_282),
.Y(n_297)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_291),
.C(n_276),
.Y(n_294)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_273),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_231),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_283),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_285),
.C(n_288),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_236),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_262),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_256),
.B(n_234),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_267),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_236),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_234),
.Y(n_289)
);

AOI21xp33_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_209),
.B(n_212),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_257),
.A2(n_252),
.B1(n_208),
.B2(n_237),
.Y(n_290)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_254),
.CI(n_272),
.CON(n_292),
.SN(n_292)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_293),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_294),
.B(n_300),
.Y(n_318)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_270),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_299),
.C(n_305),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_258),
.C(n_261),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_269),
.B(n_208),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_301),
.A2(n_290),
.B1(n_218),
.B2(n_278),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_221),
.C(n_212),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_221),
.C(n_218),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_305),
.C(n_300),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_314),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_309),
.B(n_310),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_285),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_295),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_281),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_314),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_180),
.C(n_298),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_292),
.Y(n_315)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_315),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_292),
.A2(n_299),
.B1(n_293),
.B2(n_294),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_326),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_307),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_324),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_313),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_319),
.Y(n_328)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_328),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_330),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_308),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_327),
.Y(n_334)
);

A2O1A1O1Ixp25_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_326),
.B(n_323),
.C(n_332),
.D(n_307),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_311),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_329),
.C(n_312),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_331),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_318),
.Y(n_339)
);


endmodule