module fake_jpeg_24120_n_82 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_82);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_82;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_49),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_49),
.B(n_45),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_39),
.B1(n_33),
.B2(n_38),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_34),
.B1(n_44),
.B2(n_41),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_56),
.B1(n_0),
.B2(n_2),
.Y(n_60)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_55),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_59),
.Y(n_63)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_4),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_57),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_58),
.B(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_65),
.Y(n_69)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_3),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_54),
.B(n_7),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_17),
.Y(n_73)
);

AOI22x1_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_73),
.B(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_69),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_71),
.B1(n_19),
.B2(n_20),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_30),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_23),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_25),
.Y(n_82)
);


endmodule