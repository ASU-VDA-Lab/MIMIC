module fake_aes_8086_n_29 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_29);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx2_ASAP7_75t_L g8 ( .A(n_3), .Y(n_8) );
INVx4_ASAP7_75t_L g9 ( .A(n_1), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_2), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g13 ( .A(n_0), .B(n_6), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
AOI21xp5_ASAP7_75t_L g15 ( .A1(n_10), .A2(n_0), .B(n_1), .Y(n_15) );
AOI21xp5_ASAP7_75t_L g16 ( .A1(n_10), .A2(n_1), .B(n_2), .Y(n_16) );
OAI21xp5_ASAP7_75t_L g17 ( .A1(n_8), .A2(n_3), .B(n_4), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_14), .B(n_9), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_18), .B(n_15), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_20), .B(n_9), .Y(n_22) );
OAI221xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_19), .B1(n_16), .B2(n_13), .C(n_11), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_22), .B(n_19), .Y(n_24) );
AOI32xp33_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_4), .A3(n_5), .B1(n_7), .B2(n_24), .Y(n_25) );
NOR3xp33_ASAP7_75t_L g26 ( .A(n_23), .B(n_5), .C(n_7), .Y(n_26) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_25), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_27), .B(n_28), .Y(n_29) );
endmodule