module fake_jpeg_17142_n_176 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_34),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_30),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_1),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_76),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

BUFx2_ASAP7_75t_SL g85 ( 
.A(n_78),
.Y(n_85)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_64),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_67),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_70),
.B1(n_59),
.B2(n_60),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_50),
.B1(n_49),
.B2(n_62),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_93),
.Y(n_102)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_61),
.Y(n_100)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_97),
.B(n_100),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_52),
.B(n_58),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_103),
.B1(n_119),
.B2(n_121),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_106),
.Y(n_124)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_69),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_50),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_48),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_48),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_69),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_86),
.B(n_54),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_86),
.B(n_54),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_0),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_122),
.A2(n_62),
.B1(n_63),
.B2(n_4),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_65),
.B1(n_57),
.B2(n_25),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_123),
.B(n_127),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_1),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_23),
.B1(n_46),
.B2(n_44),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_21),
.B1(n_41),
.B2(n_39),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_134),
.B(n_135),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_13),
.B1(n_38),
.B2(n_37),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_133),
.B(n_100),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_139),
.A2(n_143),
.B(n_131),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_102),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_145),
.B(n_147),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_127),
.B1(n_111),
.B2(n_120),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_146),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_140),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_131),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_136),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_148),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_125),
.B(n_130),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_132),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_156),
.B1(n_141),
.B2(n_151),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_158),
.A2(n_150),
.B1(n_126),
.B2(n_112),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_157),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_149),
.B1(n_137),
.B2(n_129),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_162),
.B(n_159),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_137),
.B1(n_26),
.B2(n_27),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_164),
.B(n_22),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_101),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_11),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_24),
.C(n_31),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_9),
.C(n_8),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_32),
.B(n_47),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_7),
.C(n_36),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_33),
.C(n_4),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_3),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_3),
.B(n_5),
.Y(n_176)
);


endmodule