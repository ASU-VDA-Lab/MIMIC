module fake_jpeg_30701_n_477 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_477);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_477;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_10),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_9),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_2),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_7),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_57),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_7),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_59),
.B(n_63),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_60),
.B(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_8),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_76),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_8),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_31),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_64),
.B(n_86),
.Y(n_131)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_6),
.C(n_14),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_70),
.B(n_78),
.Y(n_146)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_31),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_6),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_83),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_17),
.B(n_6),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_17),
.B(n_9),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_85),
.B(n_91),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_25),
.B(n_5),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_44),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_23),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_41),
.B1(n_40),
.B2(n_26),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_30),
.B1(n_25),
.B2(n_40),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_59),
.A2(n_30),
.B1(n_28),
.B2(n_42),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_41),
.B1(n_34),
.B2(n_32),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_51),
.A2(n_41),
.B1(n_28),
.B2(n_42),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_112),
.A2(n_137),
.B1(n_147),
.B2(n_33),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_68),
.A2(n_47),
.B1(n_24),
.B2(n_35),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_149),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_49),
.A2(n_34),
.B1(n_35),
.B2(n_47),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_50),
.A2(n_34),
.B1(n_32),
.B2(n_27),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_75),
.A2(n_27),
.B1(n_29),
.B2(n_34),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_56),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_78),
.Y(n_174)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_52),
.A2(n_53),
.B1(n_58),
.B2(n_66),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_69),
.A2(n_34),
.B1(n_29),
.B2(n_20),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_151),
.Y(n_225)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_153),
.B(n_155),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_134),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_160),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_116),
.B(n_74),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_98),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_157),
.B(n_176),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_39),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_158),
.B(n_161),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

HAxp5_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_78),
.CON(n_160),
.SN(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_39),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_16),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_164),
.B(n_171),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_108),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_166),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_99),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_167),
.B(n_180),
.Y(n_220)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_168),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_101),
.A2(n_82),
.B1(n_88),
.B2(n_81),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_169),
.A2(n_130),
.B1(n_127),
.B2(n_117),
.Y(n_232)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_106),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_189),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_174),
.Y(n_233)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_97),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_113),
.Y(n_177)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_92),
.B(n_71),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_145),
.B(n_39),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_114),
.A2(n_62),
.B1(n_95),
.B2(n_90),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_185),
.B1(n_149),
.B2(n_123),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

BUFx2_ASAP7_75t_SL g224 ( 
.A(n_182),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_183),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_194),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_114),
.A2(n_62),
.B1(n_87),
.B2(n_93),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_129),
.Y(n_187)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_115),
.B(n_16),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_132),
.A2(n_23),
.B1(n_20),
.B2(n_39),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_191),
.B(n_16),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_104),
.B(n_120),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_111),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_100),
.B(n_56),
.C(n_23),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_138),
.C(n_143),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_138),
.B(n_39),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_96),
.Y(n_195)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_196),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_134),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_16),
.Y(n_227)
);

BUFx2_ASAP7_75t_SL g198 ( 
.A(n_99),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_198),
.Y(n_213)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_199),
.Y(n_238)
);

AO22x1_ASAP7_75t_L g200 ( 
.A1(n_126),
.A2(n_16),
.B1(n_39),
.B2(n_20),
.Y(n_200)
);

AO22x1_ASAP7_75t_SL g218 ( 
.A1(n_200),
.A2(n_117),
.B1(n_127),
.B2(n_132),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_209),
.B(n_141),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_211),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_218),
.A2(n_162),
.B1(n_187),
.B2(n_182),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_221),
.B(n_229),
.Y(n_251)
);

NAND2xp33_ASAP7_75t_SL g226 ( 
.A(n_200),
.B(n_143),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_226),
.A2(n_183),
.B(n_151),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_109),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_158),
.B(n_125),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_189),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_172),
.B(n_109),
.C(n_118),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_236),
.C(n_193),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_232),
.A2(n_191),
.B1(n_130),
.B2(n_110),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_172),
.B(n_133),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_166),
.B1(n_163),
.B2(n_164),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_161),
.B(n_150),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_243),
.B(n_244),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_173),
.B(n_141),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_159),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_245),
.B(n_252),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_246),
.B(n_247),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_156),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_249),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_250),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_164),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_171),
.B1(n_178),
.B2(n_200),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_253),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_257),
.B1(n_261),
.B2(n_276),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_206),
.A2(n_160),
.B1(n_175),
.B2(n_170),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_189),
.B1(n_186),
.B2(n_179),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_228),
.A2(n_206),
.B1(n_242),
.B2(n_236),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_205),
.A2(n_199),
.B1(n_196),
.B2(n_152),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_221),
.B(n_195),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_264),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_224),
.Y(n_264)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_266),
.A2(n_278),
.B(n_255),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_197),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_269),
.Y(n_290)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_217),
.Y(n_268)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_204),
.B(n_168),
.Y(n_270)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_202),
.Y(n_271)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_271),
.Y(n_295)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_272),
.Y(n_311)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_202),
.Y(n_273)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_273),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_210),
.B(n_154),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_274),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_220),
.B(n_23),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_275),
.A2(n_208),
.B1(n_235),
.B2(n_225),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_232),
.A2(n_177),
.B1(n_184),
.B2(n_165),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_226),
.A2(n_190),
.B1(n_184),
.B2(n_2),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_256),
.B1(n_261),
.B2(n_276),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_222),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_205),
.B(n_0),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_248),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_239),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_207),
.B1(n_213),
.B2(n_237),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_218),
.A2(n_201),
.B1(n_214),
.B2(n_223),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_281),
.A2(n_283),
.B1(n_207),
.B2(n_225),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_209),
.B(n_0),
.C(n_1),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_231),
.C(n_203),
.Y(n_289)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_234),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_286),
.B(n_289),
.Y(n_337)
);

OAI32xp33_ASAP7_75t_L g291 ( 
.A1(n_247),
.A2(n_218),
.A3(n_203),
.B1(n_223),
.B2(n_215),
.Y(n_291)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_249),
.C(n_259),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_301),
.C(n_308),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_296),
.A2(n_300),
.B1(n_304),
.B2(n_316),
.Y(n_350)
);

NAND2x1_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_203),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_297),
.A2(n_299),
.B(n_303),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_212),
.B1(n_238),
.B2(n_241),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_252),
.B(n_212),
.C(n_241),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_266),
.A2(n_253),
.B(n_267),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_257),
.A2(n_208),
.B1(n_214),
.B2(n_234),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_251),
.B(n_279),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_317),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_312),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_246),
.A2(n_235),
.B(n_240),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_314),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_278),
.A2(n_240),
.B1(n_3),
.B2(n_1),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_258),
.A2(n_4),
.B(n_5),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_255),
.A2(n_260),
.B(n_264),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_15),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_250),
.A2(n_4),
.B1(n_12),
.B2(n_13),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_320),
.A2(n_263),
.B1(n_268),
.B2(n_272),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_287),
.B(n_282),
.C(n_254),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_332),
.C(n_342),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_285),
.B(n_270),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_327),
.B(n_346),
.Y(n_375)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_295),
.Y(n_328)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_328),
.Y(n_357)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_309),
.Y(n_330)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_315),
.A2(n_250),
.B1(n_265),
.B2(n_263),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_331),
.A2(n_347),
.B1(n_298),
.B2(n_294),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_287),
.B(n_293),
.C(n_286),
.Y(n_332)
);

OA22x2_ASAP7_75t_L g333 ( 
.A1(n_296),
.A2(n_273),
.B1(n_271),
.B2(n_283),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_345),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_334),
.A2(n_344),
.B(n_338),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_292),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_335),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_12),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_336),
.Y(n_367)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_313),
.Y(n_339)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_339),
.Y(n_365)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_340),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_316),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_341),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_1),
.C(n_3),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_343),
.A2(n_317),
.B(n_304),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_3),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_305),
.B(n_15),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_306),
.B(n_319),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_312),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_348),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_301),
.B(n_314),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_351),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_337),
.B(n_290),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_356),
.B(n_379),
.Y(n_392)
);

NOR3xp33_ASAP7_75t_SL g358 ( 
.A(n_336),
.B(n_297),
.C(n_303),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_358),
.B(n_327),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_289),
.C(n_315),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_371),
.C(n_324),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_350),
.A2(n_318),
.B1(n_291),
.B2(n_288),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_362),
.A2(n_373),
.B1(n_331),
.B2(n_321),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_326),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_329),
.A2(n_300),
.B(n_288),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_366),
.A2(n_326),
.B(n_324),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_368),
.A2(n_378),
.B1(n_341),
.B2(n_322),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_308),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_345),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_334),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_333),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_323),
.B(n_297),
.C(n_294),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_323),
.B(n_311),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_329),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_350),
.A2(n_298),
.B1(n_311),
.B2(n_322),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_349),
.B(n_325),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_381),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_382),
.A2(n_388),
.B(n_389),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_400),
.C(n_376),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_398),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_343),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_385),
.B(n_397),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_386),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_347),
.Y(n_387)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_387),
.Y(n_407)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_365),
.Y(n_390)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_365),
.Y(n_391)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_391),
.Y(n_411)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_375),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_393),
.B(n_353),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_335),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_395),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_356),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_402),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_321),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_374),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_401),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_353),
.B(n_342),
.C(n_333),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_379),
.B(n_346),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_371),
.B(n_333),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_377),
.Y(n_408)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_408),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_392),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_397),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_382),
.A2(n_366),
.B(n_352),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_413),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_396),
.C(n_400),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_419),
.C(n_355),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_402),
.B(n_352),
.C(n_373),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_403),
.A2(n_370),
.B1(n_362),
.B2(n_354),
.Y(n_421)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_421),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_417),
.B(n_380),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_426),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_413),
.A2(n_399),
.B1(n_381),
.B2(n_385),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_423),
.A2(n_418),
.B1(n_406),
.B2(n_405),
.Y(n_444)
);

NOR2xp67_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_358),
.Y(n_424)
);

OAI321xp33_ASAP7_75t_L g442 ( 
.A1(n_424),
.A2(n_425),
.A3(n_423),
.B1(n_404),
.B2(n_420),
.C(n_412),
.Y(n_442)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_408),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_410),
.A2(n_386),
.B1(n_354),
.B2(n_363),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_433),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_429),
.B(n_435),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_411),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_431),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_392),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_434),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_417),
.B(n_357),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_416),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_435),
.Y(n_437)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_437),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_426),
.A2(n_410),
.B(n_415),
.Y(n_438)
);

O2A1O1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_448),
.B(n_441),
.C(n_436),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_428),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_427),
.Y(n_450)
);

AOI211xp5_ASAP7_75t_L g441 ( 
.A1(n_425),
.A2(n_405),
.B(n_419),
.C(n_411),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_SL g457 ( 
.A(n_441),
.B(n_442),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_444),
.B(n_445),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_414),
.C(n_406),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_453),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_445),
.B(n_414),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_451),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_446),
.B(n_444),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_452),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_432),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_447),
.B(n_420),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_455),
.B(n_458),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_456),
.A2(n_364),
.B(n_361),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_439),
.A2(n_355),
.B(n_364),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_438),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_459),
.B(n_333),
.Y(n_464)
);

NOR3xp33_ASAP7_75t_L g462 ( 
.A(n_457),
.B(n_437),
.C(n_328),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_SL g467 ( 
.A(n_462),
.B(n_463),
.C(n_464),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_465),
.A2(n_449),
.B(n_454),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_468),
.A2(n_469),
.B(n_470),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_460),
.A2(n_456),
.B(n_459),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_461),
.Y(n_470)
);

OAI21x1_ASAP7_75t_L g471 ( 
.A1(n_467),
.A2(n_452),
.B(n_453),
.Y(n_471)
);

A2O1A1Ixp33_ASAP7_75t_L g474 ( 
.A1(n_471),
.A2(n_466),
.B(n_378),
.C(n_351),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_472),
.A2(n_466),
.B(n_340),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_473),
.B(n_474),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_475),
.A2(n_361),
.B(n_339),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_476),
.B(n_330),
.Y(n_477)
);


endmodule