module real_jpeg_17343_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_0),
.A2(n_207),
.B1(n_212),
.B2(n_214),
.Y(n_206)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_0),
.Y(n_215)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_1),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_3),
.A2(n_51),
.B1(n_120),
.B2(n_123),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_3),
.A2(n_51),
.B1(n_151),
.B2(n_154),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_3),
.A2(n_51),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_4),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_4),
.A2(n_27),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_4),
.B(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_4),
.A2(n_27),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_4),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_4),
.B(n_125),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_4),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_4),
.B(n_196),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_5),
.Y(n_146)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_5),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_5),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_6),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_6),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_7),
.A2(n_338),
.B1(n_343),
.B2(n_344),
.Y(n_337)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_7),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_8),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_10),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_10),
.Y(n_153)
);

BUFx4f_ASAP7_75t_L g342 ( 
.A(n_10),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_319),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_219),
.B(n_317),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_181),
.Y(n_16)
);

NOR2x1_ASAP7_75t_L g318 ( 
.A(n_17),
.B(n_181),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.C(n_167),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_18),
.B(n_224),
.Y(n_223)
);

XOR2x1_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_55),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_21),
.B(n_57),
.C(n_82),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_21),
.A2(n_22),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_31),
.B1(n_41),
.B2(n_49),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_23),
.A2(n_31),
.B1(n_41),
.B2(n_49),
.Y(n_185)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_39),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_27),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_27),
.B(n_54),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_27),
.B(n_281),
.Y(n_280)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21x1_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_38),
.B(n_41),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_32),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_41),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_42),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_42),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_82),
.B2(n_83),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_67),
.B(n_76),
.Y(n_57)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_58),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_58),
.A2(n_67),
.B1(n_76),
.B2(n_198),
.Y(n_233)
);

NAND2x1p5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_62),
.Y(n_248)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_66),
.Y(n_283)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_67),
.Y(n_196)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_70),
.Y(n_211)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_74),
.Y(n_277)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_76),
.Y(n_194)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_82),
.A2(n_83),
.B1(n_193),
.B2(n_218),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_82),
.Y(n_310)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22x1_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_107),
.B1(n_119),
.B2(n_125),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_84),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_84),
.A2(n_107),
.B(n_125),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_100),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_91),
.B1(n_95),
.B2(n_99),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_96),
.Y(n_241)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g168 ( 
.A1(n_100),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_168)
);

OA22x2_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_102),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g271 ( 
.A(n_102),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_107),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_111),
.Y(n_237)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g235 ( 
.A1(n_113),
.A2(n_236),
.A3(n_238),
.B1(n_239),
.B2(n_242),
.Y(n_235)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_126),
.B(n_167),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_142),
.B2(n_143),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_142),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_139),
.B2(n_141),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_142),
.A2(n_143),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_143),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_143),
.B(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_143),
.B(n_295),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_150),
.B1(n_157),
.B2(n_161),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_144),
.B(n_252),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_144),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_153),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_153),
.Y(n_344)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_159),
.Y(n_254)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g250 ( 
.A(n_161),
.Y(n_250)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_163),
.Y(n_279)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_172),
.C(n_174),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_184)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_172),
.A2(n_174),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

NOR2xp67_ASAP7_75t_SL g285 ( 
.A(n_174),
.B(n_286),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_179),
.B(n_180),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_206),
.B(n_216),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_188),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_182),
.B(n_189),
.C(n_192),
.Y(n_322)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_183),
.B(n_185),
.C(n_232),
.Y(n_324)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_228),
.B1(n_229),
.B2(n_232),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_204),
.B1(n_205),
.B2(n_218),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_193),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_193),
.A2(n_218),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

NAND2xp33_ASAP7_75t_R g299 ( 
.A(n_193),
.B(n_269),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_193),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_193),
.B(n_205),
.Y(n_331)
);

AO22x2_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_206),
.A2(n_336),
.B1(n_337),
.B2(n_345),
.Y(n_335)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_213),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_255),
.B(n_316),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_223),
.B(n_225),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_233),
.C(n_234),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_226),
.A2(n_227),
.B1(n_312),
.B2(n_314),
.Y(n_311)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp67_ASAP7_75t_SL g266 ( 
.A(n_231),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_231),
.B(n_267),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_262),
.C(n_263),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_233),
.A2(n_263),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_233),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_233),
.A2(n_234),
.B1(n_303),
.B2(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_233),
.A2(n_303),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_249),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_249),
.Y(n_260)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_254),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_307),
.B(n_315),
.Y(n_255)
);

OAI21x1_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_264),
.B(n_306),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_261),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_260),
.B(n_309),
.C(n_310),
.Y(n_308)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_263),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_298),
.B(n_305),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_284),
.B(n_297),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI32xp33_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_272),
.A3(n_276),
.B1(n_278),
.B2(n_280),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_294),
.B(n_296),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_291),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_300),
.Y(n_305)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_311),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_311),
.Y(n_315)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_346),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_322),
.B(n_323),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_332),
.B2(n_333),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2x1_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_331),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);


endmodule