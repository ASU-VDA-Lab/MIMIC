module fake_jpeg_11615_n_518 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_518);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_518;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_59),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_60),
.B(n_68),
.Y(n_132)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_61),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_63),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_64),
.B(n_66),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_65),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_27),
.B(n_45),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_17),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_69),
.Y(n_179)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_71),
.Y(n_182)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_26),
.B(n_15),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_85),
.Y(n_130)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_76),
.Y(n_172)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_26),
.B(n_13),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_80),
.B(n_94),
.Y(n_136)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_32),
.C(n_49),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_82),
.B(n_28),
.C(n_51),
.Y(n_151)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_38),
.B(n_12),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_86),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_88),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_91),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_38),
.B(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_92),
.B(n_111),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_93),
.Y(n_204)
);

BUFx12f_ASAP7_75t_SL g94 ( 
.A(n_32),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

CKINVDCx9p33_ASAP7_75t_R g125 ( 
.A(n_95),
.Y(n_125)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

BUFx4f_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_41),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_101),
.A2(n_85),
.B1(n_92),
.B2(n_73),
.Y(n_203)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

BUFx4f_ASAP7_75t_SL g191 ( 
.A(n_103),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_104),
.Y(n_202)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_107),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_108),
.Y(n_149)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_110),
.Y(n_147)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_57),
.B(n_0),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_112),
.B(n_113),
.Y(n_171)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_25),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_115),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_118),
.Y(n_137)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_41),
.B(n_0),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_121),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_37),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_123),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_61),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_22),
.B1(n_21),
.B2(n_43),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_126),
.A2(n_139),
.B1(n_156),
.B2(n_175),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_69),
.B(n_52),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_134),
.B(n_143),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_59),
.A2(n_22),
.B1(n_21),
.B2(n_43),
.Y(n_139)
);

AND2x4_ASAP7_75t_L g143 ( 
.A(n_60),
.B(n_54),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_103),
.A2(n_54),
.B1(n_95),
.B2(n_96),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_145),
.A2(n_168),
.B1(n_174),
.B2(n_180),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_151),
.B(n_153),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_62),
.A2(n_50),
.B1(n_51),
.B2(n_28),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_66),
.B(n_50),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_159),
.B(n_162),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_80),
.B(n_40),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_68),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_164),
.B(n_169),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_100),
.A2(n_52),
.B1(n_40),
.B2(n_34),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_64),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_34),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_173),
.B(n_187),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_104),
.A2(n_52),
.B1(n_30),
.B2(n_44),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_65),
.A2(n_30),
.B1(n_44),
.B2(n_3),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_71),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_178),
.A2(n_194),
.B1(n_203),
.B2(n_160),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_106),
.A2(n_87),
.B1(n_93),
.B2(n_91),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_75),
.A2(n_0),
.B1(n_4),
.B2(n_7),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_184),
.A2(n_125),
.B1(n_151),
.B2(n_144),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_76),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_185),
.A2(n_190),
.B1(n_196),
.B2(n_198),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_8),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_121),
.B(n_8),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_189),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_98),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_89),
.A2(n_8),
.B1(n_9),
.B2(n_123),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_82),
.A2(n_9),
.B1(n_101),
.B2(n_87),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_111),
.A2(n_9),
.B1(n_62),
.B2(n_71),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_69),
.A2(n_33),
.B1(n_57),
.B2(n_29),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_94),
.A2(n_60),
.B(n_42),
.C(n_68),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_136),
.B(n_140),
.C(n_128),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_82),
.B(n_111),
.C(n_83),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_134),
.Y(n_235)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_207),
.Y(n_287)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_208),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_128),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_209),
.B(n_218),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_171),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_211),
.B(n_221),
.Y(n_274)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_142),
.Y(n_212)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_212),
.Y(n_316)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_213),
.Y(n_293)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_146),
.Y(n_214)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_214),
.Y(n_294)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_215),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_217),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_128),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_219),
.A2(n_227),
.B1(n_250),
.B2(n_253),
.Y(n_303)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_220),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_171),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_134),
.B(n_127),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_222),
.Y(n_297)
);

AO22x1_ASAP7_75t_SL g223 ( 
.A1(n_201),
.A2(n_143),
.B1(n_127),
.B2(n_125),
.Y(n_223)
);

OA22x2_ASAP7_75t_L g308 ( 
.A1(n_223),
.A2(n_261),
.B1(n_248),
.B2(n_266),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_171),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_224),
.B(n_229),
.Y(n_275)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_184),
.A2(n_130),
.B1(n_132),
.B2(n_202),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_147),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_150),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_244),
.Y(n_278)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_152),
.Y(n_231)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_231),
.Y(n_310)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_129),
.Y(n_233)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_233),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_178),
.A2(n_147),
.B1(n_165),
.B2(n_183),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_SL g304 ( 
.A1(n_234),
.A2(n_237),
.B(n_222),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_235),
.B(n_248),
.C(n_249),
.Y(n_291)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_152),
.Y(n_236)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_236),
.Y(n_315)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_238),
.Y(n_324)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_133),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_239),
.Y(n_314)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_141),
.Y(n_240)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_240),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_177),
.B(n_161),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_241),
.B(n_246),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_138),
.B(n_143),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_243),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_143),
.B(n_137),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_163),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_179),
.Y(n_245)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_245),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_160),
.B(n_195),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_247),
.A2(n_266),
.B1(n_243),
.B2(n_242),
.Y(n_289)
);

NAND2x1_ASAP7_75t_L g248 ( 
.A(n_147),
.B(n_141),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_181),
.A2(n_197),
.B(n_195),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_135),
.A2(n_131),
.B1(n_176),
.B2(n_183),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_135),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_254),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_155),
.B(n_181),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_252),
.B(n_265),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_135),
.A2(n_131),
.B1(n_176),
.B2(n_165),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_155),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_135),
.A2(n_192),
.B1(n_182),
.B2(n_197),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_256),
.A2(n_258),
.B1(n_264),
.B2(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_259),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_182),
.A2(n_200),
.B1(n_148),
.B2(n_193),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_154),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_158),
.B(n_167),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_260),
.B(n_271),
.Y(n_281)
);

OA22x2_ASAP7_75t_L g261 ( 
.A1(n_200),
.A2(n_148),
.B1(n_167),
.B2(n_158),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_154),
.A2(n_166),
.B1(n_149),
.B2(n_133),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_166),
.B(n_191),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_172),
.A2(n_179),
.B1(n_205),
.B2(n_157),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_172),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_267),
.Y(n_276)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_157),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_270),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_191),
.B(n_186),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_269),
.B(n_259),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_157),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_186),
.B(n_191),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_196),
.A2(n_144),
.B1(n_126),
.B2(n_164),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_260),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_277),
.B(n_286),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_271),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_289),
.A2(n_302),
.B1(n_304),
.B2(n_320),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_228),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_306),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_230),
.B(n_206),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_292),
.B(n_295),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_272),
.B(n_214),
.Y(n_295)
);

A2O1A1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_263),
.A2(n_244),
.B(n_237),
.C(n_272),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_296),
.B(n_305),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_247),
.A2(n_262),
.B1(n_224),
.B2(n_211),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_263),
.C(n_226),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_255),
.B(n_233),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_312),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_256),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_250),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_313),
.B(n_317),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_253),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_219),
.A2(n_227),
.B1(n_210),
.B2(n_263),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_318),
.A2(n_288),
.B1(n_305),
.B2(n_309),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_223),
.B(n_254),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_288),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_223),
.A2(n_232),
.B1(n_251),
.B2(n_222),
.Y(n_320)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_282),
.Y(n_326)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_326),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_295),
.B(n_222),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_328),
.B(n_322),
.C(n_287),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_320),
.A2(n_249),
.B1(n_261),
.B2(n_248),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_330),
.A2(n_331),
.B1(n_347),
.B2(n_350),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_302),
.A2(n_261),
.B1(n_231),
.B2(n_236),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_291),
.A2(n_257),
.B(n_261),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_332),
.A2(n_348),
.B(n_315),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_277),
.B(n_240),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_333),
.B(n_334),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_225),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_303),
.A2(n_215),
.B1(n_216),
.B2(n_207),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_335),
.A2(n_338),
.B1(n_353),
.B2(n_355),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_291),
.A2(n_217),
.B1(n_212),
.B2(n_267),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_336),
.A2(n_356),
.B(n_363),
.Y(n_372)
);

AO22x1_ASAP7_75t_SL g337 ( 
.A1(n_308),
.A2(n_213),
.B1(n_239),
.B2(n_268),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_337),
.B(n_349),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_303),
.A2(n_220),
.B1(n_238),
.B2(n_208),
.Y(n_338)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_285),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_352),
.Y(n_365)
);

BUFx12_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_289),
.A2(n_245),
.B1(n_312),
.B2(n_317),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_278),
.A2(n_286),
.B(n_281),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_290),
.B(n_283),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_313),
.A2(n_294),
.B1(n_308),
.B2(n_297),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_325),
.Y(n_351)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_351),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_285),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_297),
.A2(n_300),
.B1(n_294),
.B2(n_308),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_283),
.B(n_296),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_354),
.B(n_361),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_300),
.A2(n_274),
.B1(n_275),
.B2(n_311),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_357),
.A2(n_314),
.B1(n_299),
.B2(n_307),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_284),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_293),
.Y(n_387)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_325),
.Y(n_360)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_360),
.Y(n_374)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_301),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_301),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_362),
.B(n_322),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_279),
.A2(n_299),
.B1(n_323),
.B2(n_314),
.Y(n_363)
);

AND2x2_ASAP7_75t_SL g364 ( 
.A(n_350),
.B(n_310),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_364),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_373),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_388),
.C(n_389),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_279),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_358),
.B(n_276),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_375),
.B(n_384),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_287),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_376),
.B(n_355),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_346),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_377),
.Y(n_400)
);

AND2x2_ASAP7_75t_SL g381 ( 
.A(n_327),
.B(n_310),
.Y(n_381)
);

NOR2x1_ASAP7_75t_R g382 ( 
.A(n_339),
.B(n_315),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_383),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_349),
.B(n_323),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_385),
.A2(n_391),
.B1(n_363),
.B2(n_336),
.Y(n_402)
);

OA22x2_ASAP7_75t_L g386 ( 
.A1(n_330),
.A2(n_327),
.B1(n_347),
.B2(n_331),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_387),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_293),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_328),
.B(n_307),
.C(n_324),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_344),
.A2(n_316),
.B(n_321),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_390),
.A2(n_338),
.B1(n_326),
.B2(n_359),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_344),
.A2(n_280),
.B1(n_324),
.B2(n_321),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_373),
.A2(n_345),
.B1(n_332),
.B2(n_341),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_393),
.A2(n_402),
.B1(n_413),
.B2(n_384),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_357),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_412),
.C(n_389),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_395),
.B(n_376),
.Y(n_419)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_370),
.Y(n_396)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_396),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_367),
.B(n_342),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_415),
.Y(n_421)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_401),
.Y(n_422)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_374),
.Y(n_404)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_404),
.Y(n_426)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_374),
.Y(n_405)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_405),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_406),
.A2(n_390),
.B(n_364),
.Y(n_438)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_369),
.Y(n_409)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_365),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_410),
.Y(n_437)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_379),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_379),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_352),
.C(n_348),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_373),
.A2(n_343),
.B1(n_329),
.B2(n_333),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_378),
.A2(n_337),
.B1(n_335),
.B2(n_334),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_414),
.A2(n_368),
.B1(n_385),
.B2(n_386),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_367),
.B(n_340),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_375),
.B(n_360),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_417),
.B(n_397),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_416),
.A2(n_380),
.B1(n_368),
.B2(n_383),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_386),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_423),
.Y(n_456)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_420),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_382),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_429),
.C(n_392),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_425),
.B(n_430),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_377),
.Y(n_427)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_427),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_366),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_428),
.B(n_407),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_366),
.C(n_386),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_410),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_400),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_432),
.B(n_436),
.Y(n_455)
);

MAJx2_ASAP7_75t_L g433 ( 
.A(n_394),
.B(n_372),
.C(n_380),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_395),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_434),
.A2(n_438),
.B1(n_440),
.B2(n_406),
.Y(n_453)
);

NOR3xp33_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_372),
.C(n_351),
.Y(n_436)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_439),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_416),
.A2(n_378),
.B1(n_381),
.B2(n_393),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_459),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_443),
.A2(n_414),
.B(n_381),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_427),
.B(n_411),
.Y(n_446)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_446),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_437),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_447),
.A2(n_441),
.B(n_403),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_409),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_448),
.B(n_449),
.Y(n_462)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_421),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_420),
.B(n_413),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_451),
.B(n_457),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_453),
.A2(n_418),
.B1(n_416),
.B2(n_438),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_454),
.B(n_423),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_392),
.C(n_403),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_401),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_460),
.Y(n_469)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_444),
.B(n_397),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_464),
.B(n_470),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_467),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_466),
.A2(n_472),
.B1(n_440),
.B2(n_447),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_456),
.B(n_419),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_434),
.Y(n_470)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_471),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_452),
.A2(n_453),
.B1(n_443),
.B2(n_450),
.Y(n_472)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_473),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_428),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_474),
.B(n_442),
.C(n_457),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_429),
.Y(n_475)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_475),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_465),
.C(n_467),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_461),
.B(n_450),
.C(n_452),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_483),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_454),
.C(n_446),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_466),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_448),
.C(n_433),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_485),
.B(n_458),
.Y(n_497)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_462),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_486),
.B(n_451),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_469),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_487),
.B(n_445),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_480),
.A2(n_468),
.B(n_473),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_489),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_483),
.A2(n_482),
.B(n_478),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_476),
.A2(n_472),
.B(n_463),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_364),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_491),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_492),
.B(n_497),
.C(n_477),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g494 ( 
.A(n_481),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_494),
.B(n_485),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_495),
.B(n_435),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_496),
.B(n_471),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_500),
.Y(n_509)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_499),
.Y(n_508)
);

AOI322xp5_ASAP7_75t_L g500 ( 
.A1(n_496),
.A2(n_484),
.A3(n_481),
.B1(n_445),
.B2(n_476),
.C1(n_460),
.C2(n_431),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_501),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_502),
.A2(n_493),
.B1(n_431),
.B2(n_422),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_364),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_507),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_510),
.B(n_479),
.C(n_505),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_512),
.A2(n_513),
.B(n_506),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_503),
.C(n_501),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_514),
.B(n_515),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_511),
.A2(n_509),
.B(n_506),
.Y(n_515)
);

AO21x1_ASAP7_75t_SL g517 ( 
.A1(n_516),
.A2(n_502),
.B(n_426),
.Y(n_517)
);

OAI32xp33_ASAP7_75t_L g518 ( 
.A1(n_517),
.A2(n_426),
.A3(n_396),
.B1(n_404),
.B2(n_405),
.Y(n_518)
);


endmodule