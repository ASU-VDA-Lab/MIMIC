module fake_jpeg_25220_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx12f_ASAP7_75t_SL g41 ( 
.A(n_18),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_21),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_19),
.B1(n_20),
.B2(n_31),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_42),
.B1(n_18),
.B2(n_20),
.Y(n_78)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_56),
.Y(n_108)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_61),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_30),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_18),
.B1(n_20),
.B2(n_19),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_62),
.A2(n_42),
.B1(n_29),
.B2(n_48),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_29),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_78),
.A2(n_87),
.B1(n_110),
.B2(n_39),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_88),
.Y(n_121)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVxp67_ASAP7_75t_SL g138 ( 
.A(n_81),
.Y(n_138)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_42),
.B1(n_37),
.B2(n_18),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_92),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_24),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_105),
.B1(n_106),
.B2(n_115),
.Y(n_133)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_31),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_40),
.C(n_39),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_47),
.Y(n_137)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_34),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_68),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_62),
.A2(n_31),
.B1(n_32),
.B2(n_25),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_54),
.B(n_47),
.Y(n_113)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_47),
.Y(n_136)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_53),
.B(n_24),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_0),
.B(n_1),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_118),
.A2(n_122),
.B(n_129),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_0),
.B(n_1),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_81),
.A2(n_66),
.B1(n_82),
.B2(n_98),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_125),
.A2(n_140),
.B1(n_124),
.B2(n_146),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_87),
.A2(n_0),
.B(n_38),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_137),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_84),
.A2(n_53),
.B1(n_25),
.B2(n_66),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_99),
.B1(n_101),
.B2(n_88),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_87),
.B(n_40),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_108),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_38),
.B(n_37),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_85),
.B1(n_83),
.B2(n_107),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_92),
.C(n_80),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_148),
.A2(n_176),
.B(n_3),
.Y(n_209)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_151),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_150),
.A2(n_159),
.B1(n_162),
.B2(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_152),
.A2(n_17),
.B(n_33),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_86),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_153),
.B(n_154),
.Y(n_211)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_23),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_127),
.B(n_120),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_94),
.B1(n_109),
.B2(n_79),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_95),
.C(n_90),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_127),
.C(n_143),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_144),
.A2(n_90),
.B1(n_25),
.B2(n_33),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_34),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_172),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_32),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_17),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_16),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_33),
.Y(n_213)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_26),
.B1(n_22),
.B2(n_33),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_175),
.A2(n_135),
.B1(n_142),
.B2(n_22),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_132),
.B(n_143),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_179),
.B1(n_181),
.B2(n_46),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_16),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_140),
.A2(n_17),
.B1(n_26),
.B2(n_22),
.Y(n_179)
);

AO21x2_ASAP7_75t_L g180 ( 
.A1(n_117),
.A2(n_49),
.B(n_46),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_135),
.B(n_49),
.Y(n_201)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_194),
.C(n_212),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_180),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_197),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_200),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_119),
.B(n_120),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_193),
.A2(n_207),
.B(n_5),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_130),
.C(n_119),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_174),
.B1(n_177),
.B2(n_166),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_142),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_3),
.B(n_4),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_208),
.Y(n_216)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_49),
.C(n_46),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_215),
.A2(n_217),
.B1(n_220),
.B2(n_233),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_195),
.A2(n_160),
.B1(n_161),
.B2(n_170),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_170),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_231),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_185),
.A2(n_168),
.B1(n_175),
.B2(n_26),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_26),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_224),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_44),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_183),
.A2(n_17),
.B1(n_4),
.B2(n_5),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_225),
.A2(n_182),
.B1(n_197),
.B2(n_196),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_3),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_229),
.A2(n_240),
.B(n_203),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_187),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_185),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_236),
.Y(n_258)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_206),
.A2(n_15),
.B1(n_8),
.B2(n_9),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_198),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_216),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_243),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_219),
.B(n_188),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_244),
.B(n_265),
.Y(n_278)
);

OA21x2_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_201),
.B(n_207),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_246),
.A2(n_228),
.B(n_222),
.Y(n_271)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_247),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_251),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_224),
.Y(n_249)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_184),
.Y(n_252)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_252),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_229),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_253),
.B(n_257),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_231),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_233),
.Y(n_273)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_188),
.C(n_212),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_234),
.C(n_217),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_261),
.A2(n_264),
.B(n_229),
.Y(n_266)
);

AO22x1_ASAP7_75t_SL g262 ( 
.A1(n_226),
.A2(n_201),
.B1(n_190),
.B2(n_196),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_262),
.A2(n_263),
.B1(n_10),
.B2(n_11),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_222),
.A2(n_202),
.B1(n_186),
.B2(n_191),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_184),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_266),
.A2(n_259),
.B(n_247),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_272),
.C(n_274),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_244),
.B(n_240),
.CI(n_220),
.CON(n_270),
.SN(n_270)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_280),
.B(n_246),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_232),
.C(n_230),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_265),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_227),
.C(n_242),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_258),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_279),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_227),
.C(n_11),
.Y(n_279)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_10),
.C(n_11),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_245),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_287),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_284),
.A2(n_253),
.B(n_254),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_292),
.B(n_295),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_291),
.A2(n_270),
.B1(n_12),
.B2(n_14),
.Y(n_311)
);

XNOR2x1_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_261),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_275),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_297),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_273),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_278),
.B(n_263),
.Y(n_296)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_262),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_299),
.C(n_271),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_262),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_15),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_294),
.A2(n_276),
.B1(n_259),
.B2(n_272),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_311),
.B1(n_290),
.B2(n_292),
.Y(n_314)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_306),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_283),
.C(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_282),
.C(n_246),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_312),
.C(n_296),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_270),
.B1(n_269),
.B2(n_13),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_302),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_10),
.C(n_12),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_319),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_298),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_320),
.B(n_304),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_321),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_313),
.A2(n_288),
.B(n_14),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_301),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_312),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_308),
.Y(n_325)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_325),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_309),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_326),
.A2(n_318),
.B(n_315),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_327),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_328),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_329),
.B(n_324),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_333),
.B(n_334),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_330),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_331),
.B(n_323),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_332),
.B(n_315),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_310),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_310),
.Y(n_340)
);


endmodule