module real_jpeg_7624_n_16 (n_5, n_4, n_8, n_0, n_12, n_345, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_346, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_345;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_346;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_1),
.A2(n_22),
.B1(n_24),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_1),
.A2(n_34),
.B1(n_69),
.B2(n_70),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_1),
.A2(n_34),
.B1(n_48),
.B2(n_51),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_2),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_2),
.A2(n_23),
.B1(n_48),
.B2(n_51),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_2),
.A2(n_23),
.B1(n_69),
.B2(n_70),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_4),
.A2(n_22),
.B1(n_24),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_4),
.A2(n_61),
.B1(n_69),
.B2(n_70),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_4),
.A2(n_48),
.B1(n_51),
.B2(n_61),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_61),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_5),
.A2(n_69),
.B1(n_70),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_5),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_5),
.A2(n_48),
.B1(n_51),
.B2(n_96),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_96),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_5),
.A2(n_22),
.B1(n_24),
.B2(n_96),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g98 ( 
.A(n_6),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_11),
.A2(n_48),
.B1(n_51),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_11),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_11),
.A2(n_69),
.B1(n_70),
.B2(n_108),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_108),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_11),
.A2(n_22),
.B1(n_24),
.B2(n_108),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_13),
.A2(n_51),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_13),
.B(n_51),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_13),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_13),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_13),
.B(n_25),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_13),
.A2(n_27),
.B(n_29),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_13),
.A2(n_22),
.B1(n_24),
.B2(n_117),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_69),
.B1(n_70),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_14),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_14),
.A2(n_48),
.B1(n_51),
.B2(n_101),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_101),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_14),
.A2(n_22),
.B1(n_24),
.B2(n_101),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_15),
.A2(n_22),
.B1(n_24),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_15),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_15),
.A2(n_48),
.B1(n_51),
.B2(n_63),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_63),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_83),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_81),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_38),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_19),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_20),
.A2(n_36),
.B(n_242),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_25),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_21),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_22),
.A2(n_26),
.B(n_31),
.C(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_31),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_22),
.A2(n_31),
.B(n_117),
.C(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_25),
.B(n_33),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_25),
.A2(n_35),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_26),
.A2(n_36),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_26),
.A2(n_36),
.B1(n_214),
.B2(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_26),
.A2(n_36),
.B1(n_223),
.B2(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_26),
.A2(n_32),
.B(n_60),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_26)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_29),
.A2(n_45),
.B(n_46),
.C(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_46),
.Y(n_55)
);

HAxp5_ASAP7_75t_SL g147 ( 
.A(n_29),
.B(n_117),
.CON(n_147),
.SN(n_147)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_35),
.A2(n_76),
.B(n_77),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_36),
.A2(n_78),
.B(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_75),
.C(n_79),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_40),
.A2(n_41),
.B1(n_340),
.B2(n_342),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_58),
.C(n_64),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_42),
.A2(n_43),
.B1(n_64),
.B2(n_319),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_53),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_44),
.A2(n_166),
.B(n_210),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_52),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_52),
.B(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_45),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_45),
.A2(n_54),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_45),
.A2(n_54),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_46),
.B(n_51),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_48),
.A2(n_55),
.B1(n_147),
.B2(n_153),
.Y(n_152)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_66),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_52),
.A2(n_54),
.B(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_53),
.A2(n_133),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_54),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_57),
.B(n_133),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_58),
.A2(n_59),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_64),
.A2(n_316),
.B1(n_319),
.B2(n_320),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_64),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_68),
.B(n_73),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_65),
.A2(n_68),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_65),
.A2(n_68),
.B1(n_107),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_65),
.A2(n_68),
.B1(n_135),
.B2(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_65),
.A2(n_145),
.B(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_65),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_65),
.A2(n_68),
.B1(n_229),
.B2(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_65),
.A2(n_249),
.B(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_68),
.B(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_68),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_68),
.B(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_68),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_69),
.B(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_69),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_109)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_74),
.B(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_74),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_75),
.A2(n_79),
.B1(n_80),
.B2(n_341),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_75),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_337),
.B(n_343),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_309),
.A3(n_330),
.B1(n_335),
.B2(n_336),
.C(n_345),
.Y(n_84)
);

AOI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_257),
.A3(n_279),
.B1(n_302),
.B2(n_308),
.C(n_346),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_216),
.C(n_253),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_187),
.B(n_215),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_160),
.B(n_186),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_140),
.B(n_159),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_128),
.B(n_139),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_114),
.B(n_127),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_93),
.B(n_102),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_97),
.B(n_157),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_98),
.B(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_120),
.B(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_109),
.B2(n_113),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_113),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_109),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_122),
.B(n_126),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_116),
.B(n_118),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_121),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_120),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_120),
.A2(n_121),
.B1(n_172),
.B2(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_120),
.A2(n_156),
.B(n_197),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_120),
.A2(n_121),
.B(n_155),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_121),
.A2(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_129),
.B(n_130),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_131),
.B(n_141),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_134),
.CI(n_136),
.CON(n_131),
.SN(n_131)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_133),
.A2(n_166),
.B1(n_168),
.B2(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_137),
.B(n_173),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_138),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_151),
.B2(n_158),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_144),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_146),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_150),
.C(n_158),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_148),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_151),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_162),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_178),
.B2(n_179),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_181),
.C(n_184),
.Y(n_188)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_169),
.B1(n_170),
.B2(n_177),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_165),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_166),
.A2(n_317),
.B(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_171),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_174),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_175),
.C(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_180),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_181),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_182),
.B(n_230),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_188),
.B(n_189),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_201),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_191),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_191),
.B(n_200),
.C(n_201),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_196),
.Y(n_219)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_211),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_208),
.B2(n_209),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_208),
.C(n_211),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_206),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_216),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_235),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_217),
.B(n_235),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_226),
.C(n_233),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_221),
.C(n_225),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_224),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_226),
.A2(n_227),
.B1(n_233),
.B2(n_234),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_232),
.Y(n_238)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_246),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_246),
.C(n_250),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_240),
.C(n_244),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_245),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_248),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_254),
.B(n_255),
.Y(n_305)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_258),
.A2(n_303),
.B(n_307),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_259),
.B(n_260),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_278),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_271),
.B2(n_272),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_272),
.C(n_278),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_266),
.C(n_270),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_270),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_268),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_269),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_277),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_274),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_273),
.A2(n_288),
.B(n_291),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_275),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_280),
.B(n_281),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_300),
.B2(n_301),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_292),
.B1(n_293),
.B2(n_299),
.Y(n_283)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_290),
.B2(n_291),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_299),
.C(n_301),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_297),
.B(n_298),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_297),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_296),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_298),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_298),
.A2(n_311),
.B1(n_321),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_300),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_323),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_310),
.B(n_323),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_321),
.C(n_322),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_311),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_312),
.A2(n_313),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_319),
.C(n_320),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_325),
.C(n_329),
.Y(n_338)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_316),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_333),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_329),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_331),
.B(n_332),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_339),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_340),
.Y(n_342)
);


endmodule