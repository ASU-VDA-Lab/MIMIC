module real_jpeg_21934_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_334, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_334;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_176;
wire n_166;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_0),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_0),
.A2(n_26),
.B1(n_32),
.B2(n_126),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_0),
.A2(n_62),
.B1(n_63),
.B2(n_126),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_0),
.A2(n_45),
.B1(n_46),
.B2(n_126),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_1),
.A2(n_26),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_1),
.A2(n_35),
.B1(n_62),
.B2(n_63),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_1),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_2),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_128),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_128),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_2),
.A2(n_26),
.B1(n_32),
.B2(n_128),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_3),
.A2(n_50),
.B1(n_62),
.B2(n_63),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_3),
.A2(n_26),
.B1(n_32),
.B2(n_50),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_4),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_4),
.B(n_28),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_4),
.A2(n_14),
.B(n_63),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_131),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_4),
.A2(n_105),
.B1(n_110),
.B2(n_190),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_4),
.B(n_87),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_4),
.B(n_30),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_4),
.A2(n_30),
.B(n_218),
.Y(n_222)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_6),
.A2(n_26),
.B1(n_32),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_6),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_133),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_133),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_133),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_7),
.B(n_62),
.Y(n_106)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_7),
.Y(n_191)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_9),
.A2(n_26),
.B1(n_32),
.B2(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_9),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_57),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_11),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_11),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_11),
.A2(n_33),
.B1(n_62),
.B2(n_63),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_282)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_13),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_14),
.A2(n_45),
.B(n_60),
.C(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_14),
.B(n_45),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_15),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_94),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_78),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_73),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_20),
.A2(n_21),
.B1(n_70),
.B2(n_320),
.Y(n_326)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_37),
.B1(n_38),
.B2(n_69),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_23),
.A2(n_36),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_23),
.A2(n_36),
.B1(n_144),
.B2(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_23),
.A2(n_266),
.B(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_23),
.A2(n_84),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_24),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_24),
.A2(n_28),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_26),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_25),
.B(n_30),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g130 ( 
.A(n_26),
.B(n_131),
.CON(n_130),
.SN(n_130)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_27),
.A2(n_29),
.B1(n_130),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_28),
.B(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_28),
.B(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g217 ( 
.A1(n_29),
.A2(n_44),
.A3(n_45),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_42),
.B(n_43),
.C(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_43),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_31),
.A2(n_36),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_58),
.B1(n_67),
.B2(n_68),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_51),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_41),
.A2(n_52),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_49),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_42),
.A2(n_53),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_42),
.A2(n_53),
.B1(n_163),
.B2(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_42),
.A2(n_51),
.B(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_42),
.A2(n_53),
.B1(n_76),
.B2(n_282),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g219 ( 
.A(n_43),
.B(n_46),
.Y(n_219)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_46),
.A2(n_64),
.B(n_131),
.C(n_181),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_75),
.B(n_77),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_52),
.A2(n_87),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_52),
.A2(n_77),
.B(n_88),
.Y(n_268)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_68),
.C(n_69),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_58),
.A2(n_67),
.B1(n_74),
.B2(n_323),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_61),
.B(n_65),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_59),
.A2(n_65),
.B(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_59),
.A2(n_61),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_59),
.A2(n_61),
.B1(n_185),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_59),
.A2(n_61),
.B1(n_206),
.B2(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_59),
.A2(n_225),
.B(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_59),
.A2(n_61),
.B1(n_113),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_59),
.A2(n_121),
.B(n_258),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_61),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_61),
.B(n_131),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_62),
.B(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_66),
.B(n_122),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_70),
.C(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_70),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_70),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_73),
.B(n_326),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_74),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_317),
.A3(n_327),
.B1(n_330),
.B2(n_331),
.C(n_334),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_297),
.B(n_316),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_273),
.B(n_296),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_165),
.B(n_249),
.C(n_272),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_149),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_99),
.B(n_149),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_134),
.B2(n_148),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_118),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_102),
.B(n_118),
.C(n_148),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_112),
.B2(n_117),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_103),
.B(n_117),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B(n_108),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_105),
.A2(n_107),
.B1(n_110),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_105),
.A2(n_174),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_105),
.A2(n_177),
.B(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_105),
.A2(n_191),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_106),
.B(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_106),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_106),
.A2(n_109),
.B(n_210),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_110),
.A2(n_139),
.B(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_110),
.B(n_131),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_114),
.B(n_240),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_115),
.B(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_129),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_127),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_129),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_140),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_135),
.B(n_141),
.C(n_146),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_138),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_154),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_150),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.C(n_161),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_158),
.B(n_208),
.Y(n_256)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_161),
.B(n_235),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_248),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_243),
.B(n_247),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_230),
.B(n_242),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_212),
.B(n_229),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_198),
.B(n_211),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_186),
.B(n_197),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_178),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_178),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_182),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_192),
.B(n_196),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_189),
.Y(n_196)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_199),
.B(n_200),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_205),
.C(n_207),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_210),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_214),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_220),
.B1(n_227),
.B2(n_228),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_217),
.Y(n_241)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_221),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_226),
.C(n_227),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_231),
.B(n_232),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_238),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_239),
.C(n_241),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_244),
.B(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_250),
.B(n_251),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_270),
.B2(n_271),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_259),
.B2(n_260),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_260),
.C(n_271),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_257),
.Y(n_279)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_269),
.Y(n_260)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_268),
.C(n_269),
.Y(n_295)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_270),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_274),
.B(n_275),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_295),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_288),
.B2(n_289),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_289),
.C(n_295),
.Y(n_298)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_283),
.C(n_287),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_283),
.B1(n_284),
.B2(n_287),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_281),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_286),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_293),
.B2(n_294),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_290),
.A2(n_291),
.B1(n_311),
.B2(n_313),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_290),
.A2(n_307),
.B(n_311),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_293),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_293),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_298),
.B(n_299),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_314),
.B2(n_315),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_306),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_306),
.C(n_315),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B(n_305),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_304),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_319),
.C(n_324),
.Y(n_318)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_305),
.B(n_319),
.CI(n_324),
.CON(n_329),
.SN(n_329)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_311),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_314),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_325),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_325),
.Y(n_331)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_328),
.B(n_329),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_329),
.Y(n_333)
);


endmodule