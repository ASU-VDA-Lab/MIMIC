module fake_aes_12486_n_673 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_96, n_39, n_673);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_96;
input n_39;
output n_673;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx10_ASAP7_75t_L g97 ( .A(n_36), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_13), .Y(n_98) );
INVxp67_ASAP7_75t_L g99 ( .A(n_10), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_59), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_92), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_0), .Y(n_102) );
INVx3_ASAP7_75t_L g103 ( .A(n_60), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_11), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_34), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_30), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_94), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_70), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_26), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_7), .Y(n_110) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_81), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_24), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_32), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_1), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_53), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_83), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_93), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_0), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_56), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_17), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_50), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_37), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_85), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_39), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_89), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_65), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_69), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_49), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_63), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_64), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_88), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_79), .Y(n_133) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_9), .Y(n_134) );
INVx2_ASAP7_75t_SL g135 ( .A(n_51), .Y(n_135) );
AND2x2_ASAP7_75t_SL g136 ( .A(n_106), .B(n_23), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_134), .B(n_1), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_113), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_106), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_103), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_135), .B(n_2), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_103), .Y(n_142) );
AOI22xp5_ASAP7_75t_L g143 ( .A1(n_98), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_103), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_108), .Y(n_146) );
BUFx8_ASAP7_75t_L g147 ( .A(n_135), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_99), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_111), .B(n_3), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g150 ( .A1(n_102), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_116), .Y(n_151) );
OAI22x1_ASAP7_75t_SL g152 ( .A1(n_120), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_114), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_114), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_97), .Y(n_155) );
INVxp67_ASAP7_75t_SL g156 ( .A(n_149), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_140), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_140), .Y(n_158) );
NAND3xp33_ASAP7_75t_L g159 ( .A(n_139), .B(n_116), .C(n_131), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_140), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_148), .B(n_97), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_153), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_139), .B(n_117), .Y(n_163) );
INVxp67_ASAP7_75t_SL g164 ( .A(n_149), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_140), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g166 ( .A1(n_143), .A2(n_102), .B1(n_104), .B2(n_118), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_142), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_140), .Y(n_168) );
AND3x1_ASAP7_75t_L g169 ( .A(n_143), .B(n_104), .C(n_110), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_144), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_136), .A2(n_114), .B1(n_131), .B2(n_101), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_136), .A2(n_114), .B1(n_109), .B2(n_112), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_142), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_136), .A2(n_133), .B1(n_107), .B2(n_130), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
AND2x6_ASAP7_75t_L g181 ( .A(n_145), .B(n_100), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_153), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_156), .B(n_147), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_161), .B(n_137), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_164), .B(n_137), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_184), .A2(n_141), .B(n_146), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_168), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_161), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_178), .A2(n_155), .B1(n_146), .B2(n_151), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_175), .A2(n_151), .B1(n_147), .B2(n_114), .Y(n_193) );
OR2x2_ASAP7_75t_L g194 ( .A(n_166), .B(n_138), .Y(n_194) );
NOR2xp67_ASAP7_75t_SL g195 ( .A(n_184), .B(n_107), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_176), .B(n_147), .Y(n_196) );
NAND2x1_ASAP7_75t_L g197 ( .A(n_181), .B(n_115), .Y(n_197) );
INVx2_ASAP7_75t_SL g198 ( .A(n_181), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_159), .A2(n_129), .B(n_124), .C(n_122), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_168), .B(n_147), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_178), .B(n_128), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_181), .A2(n_150), .B1(n_119), .B2(n_97), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_163), .B(n_121), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_168), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_163), .B(n_121), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_181), .B(n_123), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_167), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_181), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_168), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_166), .A2(n_127), .B(n_117), .C(n_132), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_167), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_169), .A2(n_152), .B1(n_123), .B2(n_130), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_181), .B(n_125), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_159), .A2(n_132), .B(n_127), .C(n_126), .Y(n_214) );
INVxp67_ASAP7_75t_L g215 ( .A(n_169), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_181), .B(n_125), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_181), .A2(n_152), .B1(n_133), .B2(n_126), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_167), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_167), .A2(n_105), .B1(n_154), .B2(n_153), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_177), .B(n_154), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_160), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_177), .B(n_154), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_177), .Y(n_223) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_214), .A2(n_171), .B(n_157), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_223), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_186), .A2(n_171), .B(n_157), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_188), .B(n_177), .Y(n_227) );
OR2x2_ASAP7_75t_L g228 ( .A(n_194), .B(n_8), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_191), .B(n_8), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_198), .B(n_158), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_198), .B(n_158), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_208), .B(n_172), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_191), .B(n_9), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_188), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_189), .A2(n_172), .B(n_173), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_188), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_210), .A2(n_173), .B(n_160), .C(n_174), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_190), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_203), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_208), .B(n_160), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_200), .A2(n_174), .B(n_165), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_201), .B(n_10), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_200), .A2(n_174), .B(n_165), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g244 ( .A1(n_196), .A2(n_180), .B(n_179), .C(n_170), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_192), .A2(n_179), .B1(n_165), .B2(n_170), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_205), .A2(n_179), .B(n_170), .C(n_180), .Y(n_246) );
OAI21xp33_ASAP7_75t_L g247 ( .A1(n_187), .A2(n_180), .B(n_154), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_196), .A2(n_185), .B(n_183), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_190), .A2(n_204), .B(n_209), .Y(n_249) );
NOR2xp67_ASAP7_75t_L g250 ( .A(n_217), .B(n_11), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_206), .B(n_154), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_213), .B(n_12), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_204), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_216), .B(n_154), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_SL g255 ( .A1(n_214), .A2(n_183), .B(n_182), .C(n_185), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_226), .A2(n_209), .B(n_193), .Y(n_256) );
BUFx10_ASAP7_75t_L g257 ( .A(n_229), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_236), .B(n_215), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_241), .A2(n_218), .B(n_207), .Y(n_259) );
AO21x1_ASAP7_75t_L g260 ( .A1(n_252), .A2(n_220), .B(n_222), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_229), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_249), .A2(n_211), .B(n_199), .Y(n_262) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_248), .A2(n_197), .B(n_222), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_234), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_243), .A2(n_221), .B(n_223), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_234), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_242), .B(n_202), .Y(n_267) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_224), .A2(n_219), .B(n_221), .Y(n_268) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_224), .A2(n_185), .B(n_183), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_SL g270 ( .A1(n_246), .A2(n_199), .B(n_182), .C(n_212), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_228), .A2(n_223), .B1(n_195), .B2(n_153), .Y(n_271) );
AOI221xp5_ASAP7_75t_SL g272 ( .A1(n_242), .A2(n_223), .B1(n_182), .B2(n_162), .C(n_15), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_225), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_239), .A2(n_162), .B1(n_13), .B2(n_14), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_227), .A2(n_12), .B1(n_14), .B2(n_15), .Y(n_275) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_235), .A2(n_162), .B(n_55), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_233), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_269), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_264), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_269), .Y(n_280) );
OA21x2_ASAP7_75t_L g281 ( .A1(n_272), .A2(n_247), .B(n_254), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_256), .A2(n_255), .B(n_244), .Y(n_282) );
BUFx8_ASAP7_75t_L g283 ( .A(n_266), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_267), .B(n_252), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_273), .Y(n_285) );
OAI21x1_ASAP7_75t_SL g286 ( .A1(n_260), .A2(n_237), .B(n_245), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_265), .A2(n_251), .B(n_225), .Y(n_287) );
OA21x2_ASAP7_75t_L g288 ( .A1(n_276), .A2(n_253), .B(n_238), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_262), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_259), .A2(n_225), .B(n_240), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_261), .B(n_250), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_258), .B(n_225), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_270), .B(n_232), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_273), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_271), .B(n_16), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
CKINVDCx8_ASAP7_75t_R g298 ( .A(n_257), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_273), .Y(n_299) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_286), .A2(n_260), .B(n_268), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_279), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_278), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_278), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_283), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_278), .Y(n_305) );
OR2x6_ASAP7_75t_L g306 ( .A(n_286), .B(n_268), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_279), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_280), .Y(n_308) );
INVxp67_ASAP7_75t_SL g309 ( .A(n_280), .Y(n_309) );
OR2x6_ASAP7_75t_L g310 ( .A(n_299), .B(n_263), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_280), .Y(n_311) );
BUFx4f_ASAP7_75t_SL g312 ( .A(n_283), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_289), .Y(n_313) );
OR2x6_ASAP7_75t_L g314 ( .A(n_299), .B(n_263), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_283), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_289), .B(n_296), .Y(n_316) );
AOI21x1_ASAP7_75t_L g317 ( .A1(n_282), .A2(n_277), .B(n_231), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_299), .Y(n_318) );
INVx5_ASAP7_75t_L g319 ( .A(n_299), .Y(n_319) );
OR2x6_ASAP7_75t_L g320 ( .A(n_299), .B(n_257), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_283), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_299), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_297), .Y(n_323) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_295), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_297), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_297), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_288), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_296), .A2(n_257), .B1(n_274), .B2(n_270), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_298), .Y(n_329) );
AO21x2_ASAP7_75t_L g330 ( .A1(n_282), .A2(n_230), .B(n_19), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_304), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_316), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_302), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_321), .B(n_291), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_316), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_324), .B(n_291), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_316), .B(n_285), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_305), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_301), .B(n_285), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_301), .B(n_284), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_313), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_302), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_324), .B(n_295), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_305), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_305), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_307), .B(n_294), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_304), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_307), .B(n_294), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_319), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_313), .B(n_294), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_303), .B(n_292), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_304), .B(n_284), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_303), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_302), .B(n_294), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_310), .B(n_299), .Y(n_355) );
AOI211x1_ASAP7_75t_SL g356 ( .A1(n_327), .A2(n_293), .B(n_287), .C(n_290), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_312), .A2(n_298), .B1(n_292), .B2(n_281), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_315), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_308), .B(n_281), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_311), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_319), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_315), .B(n_298), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_311), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_311), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_308), .B(n_281), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_308), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_315), .B(n_285), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_309), .B(n_281), .Y(n_368) );
INVx6_ASAP7_75t_L g369 ( .A(n_319), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_321), .B(n_281), .Y(n_370) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_328), .A2(n_287), .B(n_293), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_319), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_312), .B(n_18), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_300), .B(n_288), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_300), .B(n_288), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_329), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_300), .B(n_288), .Y(n_377) );
INVxp67_ASAP7_75t_L g378 ( .A(n_329), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_300), .B(n_288), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_310), .B(n_290), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_323), .Y(n_381) );
INVx2_ASAP7_75t_SL g382 ( .A(n_329), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_320), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_341), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_341), .Y(n_385) );
NOR2x1p5_ASAP7_75t_L g386 ( .A(n_373), .B(n_327), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_332), .B(n_306), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_335), .Y(n_388) );
NAND4xp25_ASAP7_75t_L g389 ( .A(n_334), .B(n_328), .C(n_327), .D(n_325), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_336), .B(n_300), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_358), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_360), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_337), .B(n_306), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_360), .Y(n_394) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_333), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_338), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_351), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_352), .B(n_19), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_361), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_337), .B(n_306), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_381), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_354), .B(n_306), .Y(n_402) );
INVx2_ASAP7_75t_SL g403 ( .A(n_369), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_361), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_351), .B(n_306), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_338), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g407 ( .A(n_370), .B(n_306), .C(n_310), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_340), .B(n_330), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_338), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_343), .B(n_330), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_343), .B(n_326), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_339), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_354), .B(n_326), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_353), .B(n_326), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_344), .Y(n_415) );
INVx4_ASAP7_75t_L g416 ( .A(n_349), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_350), .B(n_325), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_333), .Y(n_418) );
AND3x1_ASAP7_75t_L g419 ( .A(n_331), .B(n_20), .C(n_21), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_339), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_342), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_344), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_355), .B(n_310), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_344), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_345), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_346), .Y(n_426) );
NAND2x1_ASAP7_75t_SL g427 ( .A(n_349), .B(n_322), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_350), .B(n_325), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_345), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_376), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_345), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_355), .B(n_310), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_363), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_363), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_363), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_364), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_374), .B(n_323), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_364), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_374), .B(n_323), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_364), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_375), .B(n_310), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_353), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_366), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_348), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_366), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_347), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_375), .B(n_314), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_377), .B(n_314), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_342), .Y(n_449) );
INVxp67_ASAP7_75t_SL g450 ( .A(n_368), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_368), .Y(n_451) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_361), .Y(n_452) );
NAND5xp2_ASAP7_75t_L g453 ( .A(n_362), .B(n_317), .C(n_330), .D(n_22), .E(n_21), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_377), .B(n_314), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_397), .B(n_383), .Y(n_455) );
OAI21xp33_ASAP7_75t_SL g456 ( .A1(n_386), .A2(n_372), .B(n_382), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_412), .B(n_359), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_442), .B(n_379), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_442), .B(n_379), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_384), .Y(n_460) );
OAI32xp33_ASAP7_75t_L g461 ( .A1(n_430), .A2(n_357), .A3(n_372), .B1(n_349), .B2(n_365), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_398), .A2(n_349), .B(n_382), .C(n_378), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_385), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_421), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_402), .B(n_355), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_416), .B(n_380), .Y(n_466) );
NAND2x1_ASAP7_75t_L g467 ( .A(n_416), .B(n_369), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_420), .B(n_365), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_388), .B(n_356), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_421), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_437), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_402), .B(n_355), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_445), .B(n_356), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_390), .B(n_371), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_393), .B(n_371), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_437), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_408), .B(n_371), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_419), .A2(n_367), .B(n_317), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_392), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_443), .B(n_380), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_389), .A2(n_369), .B1(n_380), .B2(n_320), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_426), .B(n_314), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_393), .B(n_380), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_394), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_416), .B(n_314), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_439), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_443), .B(n_314), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_394), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_400), .B(n_369), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_396), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_418), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_400), .B(n_322), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_444), .B(n_322), .Y(n_494) );
BUFx2_ASAP7_75t_L g495 ( .A(n_404), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_441), .B(n_322), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_401), .B(n_322), .Y(n_497) );
NOR2x1_ASAP7_75t_SL g498 ( .A(n_404), .B(n_320), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_446), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_441), .B(n_318), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_411), .B(n_318), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_410), .B(n_318), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_406), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_447), .B(n_318), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_414), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_447), .B(n_318), .Y(n_506) );
OAI22x1_ASAP7_75t_L g507 ( .A1(n_391), .A2(n_319), .B1(n_317), .B2(n_20), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_448), .B(n_319), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_448), .B(n_319), .Y(n_509) );
NAND2x1p5_ASAP7_75t_L g510 ( .A(n_399), .B(n_319), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_454), .B(n_320), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_451), .B(n_320), .Y(n_512) );
NAND2xp33_ASAP7_75t_SL g513 ( .A(n_399), .B(n_320), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_454), .B(n_22), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_413), .B(n_25), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_407), .A2(n_27), .B(n_28), .C(n_29), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_453), .B(n_31), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_411), .B(n_33), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_413), .B(n_35), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_451), .B(n_38), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_450), .B(n_40), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_414), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_449), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_431), .B(n_41), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_417), .B(n_42), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_405), .B(n_43), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_406), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_417), .B(n_44), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_387), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_428), .B(n_45), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_387), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_405), .B(n_46), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_471), .B(n_395), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_499), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_456), .A2(n_403), .B(n_427), .C(n_399), .Y(n_535) );
INVx2_ASAP7_75t_SL g536 ( .A(n_495), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_470), .Y(n_537) );
INVxp67_ASAP7_75t_L g538 ( .A(n_470), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_517), .A2(n_423), .B1(n_432), .B2(n_428), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_465), .B(n_423), .Y(n_540) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_464), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_476), .B(n_431), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_460), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_463), .Y(n_544) );
NOR2x1_ASAP7_75t_L g545 ( .A(n_462), .B(n_452), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_491), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_486), .B(n_433), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_491), .Y(n_548) );
INVx1_ASAP7_75t_SL g549 ( .A(n_513), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_472), .B(n_423), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_487), .B(n_435), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_458), .B(n_435), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_459), .B(n_436), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_459), .B(n_436), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_513), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_523), .Y(n_556) );
OAI32xp33_ASAP7_75t_L g557 ( .A1(n_464), .A2(n_438), .A3(n_440), .B1(n_429), .B2(n_434), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_467), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_483), .B(n_432), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_529), .B(n_438), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_490), .B(n_432), .Y(n_561) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_462), .B(n_452), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_479), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_505), .B(n_425), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_484), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_489), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_455), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_514), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_481), .A2(n_452), .B1(n_399), .B2(n_434), .Y(n_569) );
NOR2xp67_ASAP7_75t_L g570 ( .A(n_507), .B(n_399), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_496), .B(n_452), .Y(n_571) );
INVx2_ASAP7_75t_SL g572 ( .A(n_508), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_522), .B(n_424), .Y(n_573) );
INVxp67_ASAP7_75t_SL g574 ( .A(n_498), .Y(n_574) );
INVxp67_ASAP7_75t_SL g575 ( .A(n_492), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_500), .B(n_452), .Y(n_576) );
NAND2x2_ASAP7_75t_L g577 ( .A(n_526), .B(n_427), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_457), .B(n_440), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_504), .B(n_424), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_506), .B(n_429), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_468), .B(n_422), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_531), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_469), .B(n_422), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_492), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_L g585 ( .A1(n_517), .A2(n_415), .B(n_409), .C(n_52), .Y(n_585) );
OR2x6_ASAP7_75t_L g586 ( .A(n_485), .B(n_415), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_469), .B(n_409), .Y(n_587) );
INVx3_ASAP7_75t_L g588 ( .A(n_485), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_509), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_493), .B(n_47), .Y(n_590) );
INVxp67_ASAP7_75t_SL g591 ( .A(n_503), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_578), .B(n_502), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_584), .B(n_475), .Y(n_593) );
AOI222xp33_ASAP7_75t_L g594 ( .A1(n_574), .A2(n_478), .B1(n_474), .B2(n_473), .C1(n_477), .C2(n_502), .Y(n_594) );
AOI321xp33_ASAP7_75t_L g595 ( .A1(n_569), .A2(n_461), .A3(n_474), .B1(n_477), .B2(n_473), .C(n_480), .Y(n_595) );
NAND3x2_ASAP7_75t_L g596 ( .A(n_555), .B(n_466), .C(n_553), .Y(n_596) );
AOI322xp5_ASAP7_75t_L g597 ( .A1(n_549), .A2(n_511), .A3(n_480), .B1(n_466), .B2(n_512), .C1(n_521), .C2(n_519), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_559), .B(n_482), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_577), .A2(n_478), .B1(n_512), .B2(n_532), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_568), .A2(n_516), .B1(n_510), .B2(n_521), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_541), .A2(n_488), .B(n_516), .Y(n_601) );
OAI21xp5_ASAP7_75t_SL g602 ( .A1(n_545), .A2(n_510), .B(n_515), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_539), .A2(n_530), .B1(n_528), .B2(n_525), .Y(n_603) );
AOI322xp5_ASAP7_75t_L g604 ( .A1(n_549), .A2(n_488), .A3(n_520), .B1(n_497), .B2(n_524), .C1(n_527), .C2(n_518), .Y(n_604) );
OAI21xp33_ASAP7_75t_L g605 ( .A1(n_562), .A2(n_494), .B(n_501), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g606 ( .A1(n_535), .A2(n_520), .B1(n_524), .B2(n_162), .C(n_58), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_543), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_575), .B(n_48), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_581), .B(n_54), .Y(n_609) );
AOI222xp33_ASAP7_75t_L g610 ( .A1(n_537), .A2(n_162), .B1(n_61), .B2(n_62), .C1(n_66), .C2(n_67), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_583), .B(n_57), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_540), .B(n_550), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_561), .B(n_68), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_558), .Y(n_614) );
AOI211xp5_ASAP7_75t_SL g615 ( .A1(n_570), .A2(n_71), .B(n_72), .C(n_73), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_544), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_583), .B(n_74), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_556), .A2(n_162), .B1(n_75), .B2(n_76), .C(n_77), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_587), .B(n_582), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_587), .B(n_96), .Y(n_620) );
NOR4xp25_ASAP7_75t_L g621 ( .A(n_534), .B(n_78), .C(n_80), .D(n_82), .Y(n_621) );
AOI222xp33_ASAP7_75t_L g622 ( .A1(n_569), .A2(n_86), .B1(n_87), .B2(n_90), .C1(n_91), .C2(n_95), .Y(n_622) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_538), .B(n_585), .C(n_536), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_552), .Y(n_624) );
NAND2x1p5_ASAP7_75t_L g625 ( .A(n_558), .B(n_590), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_600), .A2(n_557), .B(n_567), .C(n_588), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_602), .A2(n_589), .B(n_572), .C(n_591), .Y(n_627) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_602), .A2(n_586), .B1(n_533), .B2(n_554), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_619), .Y(n_629) );
OAI221xp5_ASAP7_75t_SL g630 ( .A1(n_597), .A2(n_586), .B1(n_576), .B2(n_571), .C(n_542), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_594), .B(n_563), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_625), .B(n_586), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_596), .A2(n_564), .B(n_573), .Y(n_633) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_614), .A2(n_564), .B(n_573), .C(n_566), .Y(n_634) );
A2O1A1Ixp33_ASAP7_75t_L g635 ( .A1(n_605), .A2(n_547), .B(n_551), .C(n_565), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g636 ( .A1(n_601), .A2(n_560), .B(n_548), .C(n_546), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_623), .A2(n_579), .B(n_580), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_594), .B(n_624), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_599), .A2(n_606), .B1(n_614), .B2(n_616), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_621), .A2(n_615), .B(n_625), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_604), .B(n_593), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_607), .B(n_592), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_612), .B(n_598), .Y(n_643) );
AOI211xp5_ASAP7_75t_L g644 ( .A1(n_621), .A2(n_603), .B(n_613), .C(n_608), .Y(n_644) );
NOR2x1_ASAP7_75t_L g645 ( .A(n_609), .B(n_611), .Y(n_645) );
INVxp67_ASAP7_75t_L g646 ( .A(n_617), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_620), .B(n_622), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_595), .B(n_622), .C(n_610), .Y(n_648) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_618), .A2(n_600), .B(n_602), .C(n_574), .Y(n_649) );
OAI221xp5_ASAP7_75t_L g650 ( .A1(n_595), .A2(n_602), .B1(n_605), .B2(n_601), .C(n_594), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_614), .B(n_574), .Y(n_651) );
AND2x4_ASAP7_75t_L g652 ( .A(n_651), .B(n_632), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_638), .B(n_631), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_650), .A2(n_648), .B(n_630), .C(n_626), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_627), .A2(n_651), .B(n_640), .Y(n_655) );
NOR2x1p5_ASAP7_75t_L g656 ( .A(n_641), .B(n_647), .Y(n_656) );
NAND3xp33_ASAP7_75t_SL g657 ( .A(n_649), .B(n_627), .C(n_639), .Y(n_657) );
AND3x2_ASAP7_75t_L g658 ( .A(n_652), .B(n_636), .C(n_644), .Y(n_658) );
NAND4xp75_ASAP7_75t_L g659 ( .A(n_655), .B(n_645), .C(n_637), .D(n_633), .Y(n_659) );
NOR2x1_ASAP7_75t_L g660 ( .A(n_657), .B(n_628), .Y(n_660) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_654), .B(n_635), .Y(n_661) );
NAND2x1p5_ASAP7_75t_L g662 ( .A(n_661), .B(n_656), .Y(n_662) );
INVx5_ASAP7_75t_L g663 ( .A(n_658), .Y(n_663) );
NOR2x1p5_ASAP7_75t_L g664 ( .A(n_659), .B(n_653), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_662), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_664), .B(n_660), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_666), .B(n_663), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_665), .B(n_663), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_668), .B(n_643), .Y(n_669) );
NAND2xp33_ASAP7_75t_SL g670 ( .A(n_669), .B(n_667), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_670), .A2(n_639), .B(n_634), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g672 ( .A1(n_671), .A2(n_635), .B(n_646), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_672), .A2(n_642), .B(n_629), .Y(n_673) );
endmodule