module fake_jpeg_14639_n_295 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_181;
wire n_38;
wire n_26;
wire n_28;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_21),
.B1(n_31),
.B2(n_17),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_48),
.A2(n_43),
.B1(n_32),
.B2(n_20),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_68),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_21),
.B1(n_31),
.B2(n_34),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_63),
.B1(n_42),
.B2(n_43),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_21),
.B1(n_31),
.B2(n_34),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_57),
.B1(n_42),
.B2(n_45),
.Y(n_92)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx2_ASAP7_75t_SL g77 ( 
.A(n_56),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_17),
.B1(n_20),
.B2(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_17),
.B1(n_35),
.B2(n_27),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_20),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_94),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_82),
.Y(n_117)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_90),
.Y(n_118)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_97),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_93),
.B1(n_56),
.B2(n_26),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_20),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_101),
.B1(n_46),
.B2(n_66),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_100),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_58),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_37),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_104),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_48),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_37),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_1),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_108),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_39),
.C(n_30),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_109),
.B(n_112),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_39),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_39),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_132),
.B(n_26),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_121),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_73),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_126),
.B1(n_129),
.B2(n_82),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_26),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_25),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_94),
.B1(n_106),
.B2(n_86),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_25),
.Y(n_132)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_75),
.Y(n_139)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_110),
.B(n_74),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_156),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_141),
.B(n_142),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_96),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_96),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_149),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_155),
.B1(n_134),
.B2(n_125),
.Y(n_168)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_76),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_97),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_87),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_157),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_22),
.B(n_27),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_19),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_110),
.B(n_18),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_87),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_162),
.Y(n_174)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_95),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_164),
.Y(n_180)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_129),
.A2(n_77),
.B1(n_30),
.B2(n_78),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_128),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_168),
.A2(n_172),
.B1(n_176),
.B2(n_188),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_107),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_169),
.B(n_184),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_125),
.B1(n_132),
.B2(n_108),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_155),
.A2(n_123),
.B1(n_130),
.B2(n_132),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_189),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_120),
.Y(n_181)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_194),
.B1(n_158),
.B2(n_157),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_84),
.C(n_124),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_84),
.B(n_25),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_30),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_128),
.B1(n_22),
.B2(n_18),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_30),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_191),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_84),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_29),
.B(n_28),
.C(n_3),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_156),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_136),
.A2(n_29),
.B1(n_28),
.B2(n_3),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_196),
.A2(n_218),
.B(n_186),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_203),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_194),
.B(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_207),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_147),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_208),
.B(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_150),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_193),
.B(n_173),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_162),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_1),
.Y(n_234)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_188),
.B1(n_189),
.B2(n_144),
.Y(n_231)
);

AO22x1_ASAP7_75t_L g218 ( 
.A1(n_176),
.A2(n_165),
.B1(n_145),
.B2(n_144),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_183),
.B1(n_175),
.B2(n_178),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_220),
.A2(n_224),
.B1(n_204),
.B2(n_201),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_169),
.C(n_184),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_225),
.C(n_237),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_191),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_238),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_178),
.B1(n_165),
.B2(n_173),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_172),
.C(n_190),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_226),
.A2(n_232),
.B(n_202),
.Y(n_247)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

OAI22x1_ASAP7_75t_L g232 ( 
.A1(n_198),
.A2(n_192),
.B1(n_135),
.B2(n_3),
.Y(n_232)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_195),
.C(n_204),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_16),
.C(n_15),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_215),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_249),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_247),
.A2(n_220),
.B(n_229),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_227),
.B1(n_238),
.B2(n_222),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_214),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_228),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_252),
.Y(n_266)
);

NOR3xp33_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_196),
.C(n_207),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_224),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_1),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_2),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_219),
.C(n_230),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_245),
.A2(n_226),
.B(n_237),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_276)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_256),
.A2(n_264),
.B(n_248),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_262),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_266),
.C(n_259),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_13),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_239),
.B(n_223),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_253),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_4),
.B(n_5),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_258),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_240),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_274),
.Y(n_280)
);

AOI21x1_ASAP7_75t_SL g277 ( 
.A1(n_270),
.A2(n_256),
.B(n_262),
.Y(n_277)
);

NOR3xp33_ASAP7_75t_SL g272 ( 
.A(n_264),
.B(n_243),
.C(n_241),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_273),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_265),
.A2(n_241),
.B(n_240),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_276),
.B(n_269),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_268),
.B(n_272),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_279),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_260),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_13),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_281),
.A2(n_280),
.B(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_288),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_287),
.A2(n_10),
.B(n_11),
.Y(n_290)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_7),
.CI(n_8),
.CON(n_288),
.SN(n_288)
);

OA21x2_ASAP7_75t_SL g289 ( 
.A1(n_285),
.A2(n_10),
.B(n_11),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_SL g293 ( 
.A(n_289),
.B(n_10),
.C(n_284),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_288),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_293),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_291),
.Y(n_295)
);


endmodule