module fake_aes_2026_n_279 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_3, n_18, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_14, n_10, n_15, n_42, n_24, n_19, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_279);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_3;
input n_18;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_42;
input n_24;
input n_19;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_279;
wire n_117;
wire n_219;
wire n_133;
wire n_149;
wire n_220;
wire n_81;
wire n_69;
wire n_214;
wire n_267;
wire n_204;
wire n_221;
wire n_249;
wire n_185;
wire n_203;
wire n_57;
wire n_88;
wire n_244;
wire n_102;
wire n_119;
wire n_73;
wire n_141;
wire n_115;
wire n_97;
wire n_80;
wire n_167;
wire n_107;
wire n_158;
wire n_278;
wire n_60;
wire n_114;
wire n_121;
wire n_94;
wire n_65;
wire n_171;
wire n_196;
wire n_125;
wire n_192;
wire n_240;
wire n_254;
wire n_161;
wire n_262;
wire n_177;
wire n_130;
wire n_189;
wire n_103;
wire n_239;
wire n_137;
wire n_87;
wire n_180;
wire n_104;
wire n_277;
wire n_160;
wire n_98;
wire n_74;
wire n_206;
wire n_276;
wire n_154;
wire n_272;
wire n_195;
wire n_165;
wire n_146;
wire n_85;
wire n_250;
wire n_237;
wire n_181;
wire n_101;
wire n_62;
wire n_255;
wire n_215;
wire n_116;
wire n_108;
wire n_91;
wire n_155;
wire n_209;
wire n_217;
wire n_139;
wire n_229;
wire n_230;
wire n_274;
wire n_198;
wire n_169;
wire n_193;
wire n_273;
wire n_252;
wire n_152;
wire n_113;
wire n_241;
wire n_95;
wire n_124;
wire n_156;
wire n_238;
wire n_128;
wire n_120;
wire n_129;
wire n_70;
wire n_90;
wire n_71;
wire n_63;
wire n_56;
wire n_135;
wire n_188;
wire n_78;
wire n_247;
wire n_197;
wire n_201;
wire n_242;
wire n_260;
wire n_127;
wire n_170;
wire n_111;
wire n_157;
wire n_79;
wire n_202;
wire n_210;
wire n_64;
wire n_142;
wire n_184;
wire n_245;
wire n_265;
wire n_191;
wire n_264;
wire n_232;
wire n_200;
wire n_208;
wire n_211;
wire n_58;
wire n_122;
wire n_187;
wire n_138;
wire n_126;
wire n_275;
wire n_178;
wire n_118;
wire n_258;
wire n_253;
wire n_179;
wire n_84;
wire n_131;
wire n_112;
wire n_266;
wire n_205;
wire n_86;
wire n_143;
wire n_213;
wire n_235;
wire n_243;
wire n_182;
wire n_263;
wire n_166;
wire n_162;
wire n_186;
wire n_75;
wire n_163;
wire n_226;
wire n_105;
wire n_159;
wire n_174;
wire n_227;
wire n_248;
wire n_268;
wire n_231;
wire n_72;
wire n_136;
wire n_89;
wire n_76;
wire n_176;
wire n_68;
wire n_144;
wire n_183;
wire n_256;
wire n_67;
wire n_77;
wire n_216;
wire n_147;
wire n_199;
wire n_148;
wire n_123;
wire n_83;
wire n_172;
wire n_100;
wire n_212;
wire n_228;
wire n_92;
wire n_223;
wire n_251;
wire n_59;
wire n_236;
wire n_150;
wire n_218;
wire n_168;
wire n_194;
wire n_110;
wire n_261;
wire n_66;
wire n_134;
wire n_222;
wire n_234;
wire n_164;
wire n_233;
wire n_271;
wire n_82;
wire n_106;
wire n_175;
wire n_173;
wire n_190;
wire n_145;
wire n_270;
wire n_246;
wire n_153;
wire n_61;
wire n_259;
wire n_132;
wire n_99;
wire n_109;
wire n_93;
wire n_151;
wire n_140;
wire n_207;
wire n_257;
wire n_224;
wire n_96;
wire n_269;
wire n_225;
INVx2_ASAP7_75t_L g56 ( .A(n_24), .Y(n_56) );
CKINVDCx16_ASAP7_75t_R g57 ( .A(n_48), .Y(n_57) );
INVx2_ASAP7_75t_L g58 ( .A(n_52), .Y(n_58) );
INVx2_ASAP7_75t_L g59 ( .A(n_46), .Y(n_59) );
BUFx3_ASAP7_75t_L g60 ( .A(n_36), .Y(n_60) );
INVx2_ASAP7_75t_L g61 ( .A(n_41), .Y(n_61) );
INVx2_ASAP7_75t_L g62 ( .A(n_8), .Y(n_62) );
INVx1_ASAP7_75t_L g63 ( .A(n_37), .Y(n_63) );
INVx1_ASAP7_75t_L g64 ( .A(n_45), .Y(n_64) );
INVx1_ASAP7_75t_L g65 ( .A(n_40), .Y(n_65) );
INVx1_ASAP7_75t_L g66 ( .A(n_10), .Y(n_66) );
CKINVDCx5p33_ASAP7_75t_R g67 ( .A(n_30), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_15), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_7), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_9), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_18), .Y(n_71) );
CKINVDCx5p33_ASAP7_75t_R g72 ( .A(n_55), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_12), .Y(n_73) );
CKINVDCx5p33_ASAP7_75t_R g74 ( .A(n_39), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_50), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_54), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_25), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_27), .Y(n_78) );
BUFx2_ASAP7_75t_L g79 ( .A(n_38), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_6), .Y(n_80) );
INVxp33_ASAP7_75t_L g81 ( .A(n_43), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_35), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_3), .Y(n_83) );
BUFx3_ASAP7_75t_L g84 ( .A(n_23), .Y(n_84) );
BUFx3_ASAP7_75t_L g85 ( .A(n_31), .Y(n_85) );
CKINVDCx14_ASAP7_75t_R g86 ( .A(n_51), .Y(n_86) );
BUFx3_ASAP7_75t_L g87 ( .A(n_5), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_44), .Y(n_88) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_47), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_62), .Y(n_90) );
OA21x2_ASAP7_75t_L g91 ( .A1(n_56), .A2(n_26), .B(n_22), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_62), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_83), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_83), .Y(n_94) );
INVx3_ASAP7_75t_L g95 ( .A(n_87), .Y(n_95) );
AND2x4_ASAP7_75t_L g96 ( .A(n_79), .B(n_0), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_89), .Y(n_97) );
BUFx6f_ASAP7_75t_L g98 ( .A(n_89), .Y(n_98) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_89), .Y(n_99) );
HB1xp67_ASAP7_75t_L g100 ( .A(n_87), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_89), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_56), .A2(n_29), .B(n_28), .Y(n_102) );
AND2x4_ASAP7_75t_L g103 ( .A(n_58), .B(n_1), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_60), .Y(n_104) );
AND2x2_ASAP7_75t_L g105 ( .A(n_81), .B(n_2), .Y(n_105) );
AND2x4_ASAP7_75t_L g106 ( .A(n_59), .B(n_61), .Y(n_106) );
AND2x4_ASAP7_75t_L g107 ( .A(n_59), .B(n_2), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_98), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_104), .Y(n_109) );
INVx4_ASAP7_75t_SL g110 ( .A(n_103), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_104), .Y(n_111) );
AND2x6_ASAP7_75t_L g112 ( .A(n_96), .B(n_84), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_100), .B(n_57), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_103), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_103), .Y(n_115) );
INVx3_ASAP7_75t_L g116 ( .A(n_103), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_98), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_105), .B(n_86), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_107), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_107), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_105), .B(n_80), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_107), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_98), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_98), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_118), .B(n_96), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_118), .B(n_96), .Y(n_126) );
AND2x6_ASAP7_75t_L g127 ( .A(n_114), .B(n_106), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_121), .B(n_106), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_113), .B(n_95), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_114), .A2(n_106), .B1(n_95), .B2(n_92), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_110), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_116), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_115), .B(n_90), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_112), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_110), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_119), .B(n_93), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_112), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_120), .B(n_94), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_122), .B(n_67), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_122), .B(n_74), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_109), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_111), .B(n_84), .Y(n_142) );
AOI22xp5_ASAP7_75t_L g143 ( .A1(n_111), .A2(n_66), .B1(n_69), .B2(n_68), .Y(n_143) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_108), .A2(n_71), .B1(n_73), .B2(n_70), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_126), .A2(n_102), .B(n_91), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_128), .A2(n_102), .B(n_91), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_134), .B(n_85), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_125), .A2(n_102), .B(n_91), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_132), .Y(n_149) );
AND2x6_ASAP7_75t_L g150 ( .A(n_134), .B(n_88), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_132), .Y(n_151) );
AO21x1_ASAP7_75t_L g152 ( .A1(n_133), .A2(n_138), .B(n_136), .Y(n_152) );
INVx5_ASAP7_75t_L g153 ( .A(n_127), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_127), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g155 ( .A1(n_133), .A2(n_64), .B(n_65), .C(n_63), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_130), .B(n_72), .Y(n_156) );
O2A1O1Ixp5_ASAP7_75t_SL g157 ( .A1(n_141), .A2(n_75), .B(n_77), .C(n_76), .Y(n_157) );
AO21x1_ASAP7_75t_L g158 ( .A1(n_136), .A2(n_82), .B(n_78), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_131), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g161 ( .A1(n_137), .A2(n_144), .B1(n_139), .B2(n_140), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_143), .B(n_104), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_144), .B(n_4), .Y(n_163) );
AO21x1_ASAP7_75t_L g164 ( .A1(n_142), .A2(n_97), .B(n_98), .Y(n_164) );
INVx5_ASAP7_75t_L g165 ( .A(n_134), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_126), .A2(n_123), .B(n_117), .Y(n_166) );
AO21x1_ASAP7_75t_L g167 ( .A1(n_129), .A2(n_101), .B(n_99), .Y(n_167) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_145), .A2(n_101), .B(n_99), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_154), .Y(n_169) );
NOR2x1_ASAP7_75t_SL g170 ( .A(n_153), .B(n_99), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_148), .A2(n_124), .B(n_123), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_146), .A2(n_166), .B(n_161), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_151), .Y(n_175) );
AO31x2_ASAP7_75t_L g176 ( .A1(n_158), .A2(n_11), .A3(n_13), .B(n_14), .Y(n_176) );
AO31x2_ASAP7_75t_L g177 ( .A1(n_164), .A2(n_16), .A3(n_17), .B(n_19), .Y(n_177) );
AO31x2_ASAP7_75t_L g178 ( .A1(n_155), .A2(n_19), .A3(n_20), .B(n_21), .Y(n_178) );
AO31x2_ASAP7_75t_L g179 ( .A1(n_162), .A2(n_32), .A3(n_33), .B(n_34), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_163), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_165), .Y(n_181) );
INVx1_ASAP7_75t_SL g182 ( .A(n_147), .Y(n_182) );
OR2x2_ASAP7_75t_L g183 ( .A(n_156), .B(n_42), .Y(n_183) );
BUFx2_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_159), .B(n_53), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_159), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
INVx5_ASAP7_75t_L g189 ( .A(n_169), .Y(n_189) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_172), .A2(n_150), .B(n_49), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_174), .B(n_175), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_178), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_185), .A2(n_183), .B1(n_184), .B2(n_182), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_178), .Y(n_194) );
OR2x6_ASAP7_75t_L g195 ( .A(n_187), .B(n_181), .Y(n_195) );
BUFx12f_ASAP7_75t_L g196 ( .A(n_169), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_176), .B(n_181), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_186), .B(n_188), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_176), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_177), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_179), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_170), .B(n_179), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_168), .A2(n_173), .B(n_171), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_168), .A2(n_173), .B(n_171), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_168), .A2(n_173), .B(n_171), .Y(n_205) );
AO31x2_ASAP7_75t_L g206 ( .A1(n_172), .A2(n_152), .A3(n_173), .B(n_167), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_180), .B(n_172), .Y(n_207) );
AOI21x1_ASAP7_75t_L g208 ( .A1(n_171), .A2(n_173), .B(n_172), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_173), .A2(n_172), .B(n_157), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_173), .A2(n_172), .B(n_157), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_198), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_207), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_198), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_206), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_192), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_197), .B(n_202), .Y(n_216) );
BUFx2_ASAP7_75t_L g217 ( .A(n_202), .Y(n_217) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_209), .A2(n_210), .B(n_201), .Y(n_218) );
INVx6_ASAP7_75t_L g219 ( .A(n_196), .Y(n_219) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_200), .A2(n_199), .B(n_194), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_191), .Y(n_221) );
NAND2x1_ASAP7_75t_L g222 ( .A(n_190), .B(n_193), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_189), .B(n_195), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_195), .B(n_189), .Y(n_224) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_203), .A2(n_205), .B(n_204), .Y(n_225) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_203), .A2(n_205), .B(n_204), .Y(n_226) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_203), .A2(n_205), .B(n_204), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_189), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_208), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_215), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_211), .B(n_213), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_213), .B(n_212), .Y(n_232) );
INVx4_ASAP7_75t_L g233 ( .A(n_228), .Y(n_233) );
OR2x6_ASAP7_75t_L g234 ( .A(n_217), .B(n_222), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_220), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_220), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_220), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_228), .Y(n_238) );
INVx2_ASAP7_75t_SL g239 ( .A(n_228), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_216), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_229), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_221), .B(n_218), .Y(n_242) );
INVx4_ASAP7_75t_L g243 ( .A(n_223), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_242), .B(n_214), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_230), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_241), .Y(n_246) );
INVx4_ASAP7_75t_L g247 ( .A(n_233), .Y(n_247) );
INVx4_ASAP7_75t_L g248 ( .A(n_233), .Y(n_248) );
BUFx2_ASAP7_75t_L g249 ( .A(n_240), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_231), .B(n_227), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_231), .B(n_226), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_234), .B(n_226), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_232), .B(n_225), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_245), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_246), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_250), .B(n_235), .Y(n_256) );
AND2x2_ASAP7_75t_SL g257 ( .A(n_247), .B(n_243), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_251), .B(n_236), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_253), .B(n_237), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_254), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_255), .Y(n_261) );
NAND2x1p5_ASAP7_75t_L g262 ( .A(n_257), .B(n_247), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_259), .B(n_244), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_260), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_261), .Y(n_265) );
INVxp67_ASAP7_75t_SL g266 ( .A(n_262), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_266), .A2(n_248), .B1(n_243), .B2(n_263), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_265), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_264), .Y(n_269) );
NOR2xp33_ASAP7_75t_R g270 ( .A(n_269), .B(n_219), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_270), .B(n_267), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_271), .B(n_268), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_272), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_273), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_274), .Y(n_275) );
OAI222xp33_ASAP7_75t_L g276 ( .A1(n_275), .A2(n_224), .B1(n_234), .B2(n_238), .C1(n_239), .C2(n_249), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_276), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_277), .B(n_261), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_278), .A2(n_252), .B1(n_258), .B2(n_256), .Y(n_279) );
endmodule