module fake_netlist_6_4232_n_1636 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1636);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1636;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_25),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_65),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_26),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_39),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_2),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_14),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_41),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_51),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_59),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_82),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_120),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_72),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_118),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_30),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_135),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_108),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_92),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_98),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_28),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_131),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_100),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_8),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_88),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_7),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_61),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_97),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_20),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_2),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_81),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_109),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_74),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_17),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_29),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_112),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_31),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_64),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_76),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_60),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_110),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_47),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_137),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_101),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_113),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_50),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_40),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_127),
.Y(n_202)
);

BUFx8_ASAP7_75t_SL g203 ( 
.A(n_96),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_26),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_25),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_79),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_130),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_19),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_33),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_30),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_45),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_114),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_54),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_3),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_73),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_67),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_146),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_8),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_49),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_16),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_139),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_99),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_15),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_31),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_71),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_123),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_21),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_89),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_50),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_102),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_116),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_124),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_95),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_115),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_94),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_56),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_57),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_133),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_143),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_27),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_55),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_132),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_17),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_43),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_16),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_145),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_53),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_87),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_62),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_122),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_5),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_23),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_141),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_44),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_47),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_140),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_22),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_44),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_69),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_46),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_80),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_107),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_37),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_142),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_20),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_12),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_32),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_134),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_1),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_128),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_29),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_63),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_111),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_138),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_9),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_4),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_36),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_5),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_18),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_24),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_33),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_42),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_85),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_1),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_106),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_93),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_35),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_12),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_66),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_27),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_23),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_105),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_0),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_121),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_228),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_221),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_203),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_206),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_206),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_150),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_150),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_168),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_228),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_169),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_295),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_150),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_150),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_150),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_196),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_149),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_156),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_160),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_161),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_155),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_155),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_197),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_256),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_258),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_172),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_162),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_188),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_197),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_196),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_279),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_175),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_157),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_175),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_163),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_197),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_212),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_216),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_167),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_171),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_153),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_177),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_287),
.B(n_0),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_148),
.B(n_3),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_157),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_170),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_177),
.Y(n_345)
);

BUFx10_ASAP7_75t_L g346 ( 
.A(n_193),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_181),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_181),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_189),
.B(n_4),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_147),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_189),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_173),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_243),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_269),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_293),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_151),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_176),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_208),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_179),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_208),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_246),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_215),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_215),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_219),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_182),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_158),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_183),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_219),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_244),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_303),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_311),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_301),
.Y(n_372)
);

OAI21x1_ASAP7_75t_L g373 ( 
.A1(n_342),
.A2(n_165),
.B(n_148),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_301),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_312),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_305),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_302),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_310),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_346),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_300),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_302),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_324),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_326),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_313),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_316),
.B(n_191),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_297),
.B(n_202),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_336),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_158),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_314),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_316),
.B(n_192),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_319),
.B(n_165),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_325),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_327),
.B(n_190),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_307),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_308),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_308),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_346),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_328),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_346),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_R g402 ( 
.A(n_298),
.B(n_195),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_309),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_338),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_353),
.Y(n_405)
);

AND3x1_ASAP7_75t_L g406 ( 
.A(n_341),
.B(n_288),
.C(n_255),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_309),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_330),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_332),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_332),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_356),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_331),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_331),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_315),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_340),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_340),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_315),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_333),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g421 ( 
.A1(n_317),
.A2(n_174),
.B(n_164),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_337),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_354),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_316),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_355),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_R g426 ( 
.A(n_344),
.B(n_199),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_317),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_318),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_345),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_335),
.B(n_159),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_352),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_357),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_297),
.B(n_202),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_345),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_339),
.B(n_202),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_318),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_359),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_367),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_334),
.B(n_190),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_366),
.B(n_207),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_365),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_388),
.A2(n_395),
.B1(n_439),
.B2(n_393),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_306),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_430),
.B(n_350),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_339),
.Y(n_446)
);

NAND3xp33_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_299),
.C(n_296),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_393),
.B(n_198),
.Y(n_448)
);

INVx5_ASAP7_75t_L g449 ( 
.A(n_379),
.Y(n_449)
);

INVx5_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_404),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_L g452 ( 
.A(n_379),
.B(n_193),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_388),
.B(n_320),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_424),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_424),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_385),
.B(n_238),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_440),
.B(n_371),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_385),
.Y(n_458)
);

BUFx4f_ASAP7_75t_L g459 ( 
.A(n_421),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_372),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_393),
.B(n_395),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_406),
.A2(n_361),
.B1(n_220),
.B2(n_294),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_372),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_393),
.B(n_198),
.Y(n_464)
);

BUFx4f_ASAP7_75t_L g465 ( 
.A(n_421),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_408),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_412),
.B(n_420),
.C(n_388),
.Y(n_467)
);

NOR2x1p5_ASAP7_75t_L g468 ( 
.A(n_432),
.B(n_349),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_304),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_379),
.Y(n_470)
);

AND2x6_ASAP7_75t_L g471 ( 
.A(n_395),
.B(n_231),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_374),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_392),
.Y(n_473)
);

BUFx10_ASAP7_75t_L g474 ( 
.A(n_375),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_395),
.B(n_193),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_374),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_379),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_379),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_379),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_380),
.Y(n_480)
);

INVx4_ASAP7_75t_SL g481 ( 
.A(n_389),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_384),
.B(n_255),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_409),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_439),
.B(n_213),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_401),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_390),
.B(n_288),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_439),
.B(n_193),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_409),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_439),
.B(n_406),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_380),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_374),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_410),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_439),
.B(n_320),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_401),
.B(n_217),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_402),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_401),
.B(n_218),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_389),
.B(n_226),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_426),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_404),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_394),
.B(n_419),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_389),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_411),
.B(n_164),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_389),
.B(n_227),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_422),
.B(n_349),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_386),
.A2(n_187),
.B1(n_289),
.B2(n_291),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_389),
.B(n_193),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_420),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_411),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_432),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_431),
.B(n_152),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_381),
.Y(n_512)
);

BUFx8_ASAP7_75t_SL g513 ( 
.A(n_370),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_416),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_389),
.B(n_174),
.Y(n_515)
);

INVx4_ASAP7_75t_SL g516 ( 
.A(n_389),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_399),
.B(n_178),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_437),
.B(n_154),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_399),
.B(n_178),
.Y(n_519)
);

AO22x2_ASAP7_75t_L g520 ( 
.A1(n_435),
.A2(n_272),
.B1(n_244),
.B2(n_253),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_399),
.B(n_233),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_378),
.B(n_347),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_441),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_426),
.Y(n_524)
);

OR2x2_ASAP7_75t_SL g525 ( 
.A(n_435),
.B(n_253),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_416),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_391),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_399),
.B(n_234),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_438),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_L g530 ( 
.A(n_399),
.B(n_184),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_391),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_399),
.B(n_236),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_378),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_399),
.B(n_237),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_377),
.B(n_239),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_417),
.Y(n_536)
);

AND2x2_ASAP7_75t_SL g537 ( 
.A(n_421),
.B(n_184),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_432),
.B(n_202),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_421),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_396),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_396),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_417),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_386),
.B(n_433),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_421),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_429),
.Y(n_545)
);

OAI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_433),
.A2(n_229),
.B1(n_223),
.B2(n_290),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_377),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_400),
.B(n_186),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_397),
.B(n_242),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_407),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_429),
.B(n_166),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_434),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_418),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_396),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_413),
.B(n_248),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_413),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_413),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_418),
.B(n_180),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_418),
.A2(n_224),
.B1(n_292),
.B2(n_210),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_373),
.A2(n_276),
.B1(n_272),
.B2(n_270),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_373),
.B(n_186),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_398),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_414),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_414),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_414),
.B(n_249),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_373),
.A2(n_261),
.B1(n_264),
.B2(n_276),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_402),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_L g568 ( 
.A(n_398),
.B(n_194),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_403),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_403),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_403),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_418),
.B(n_185),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_415),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_415),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_427),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_427),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_427),
.B(n_194),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_428),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_428),
.B(n_251),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_436),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_458),
.B(n_200),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_442),
.B(n_254),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_485),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_480),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_457),
.B(n_257),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_494),
.B(n_347),
.Y(n_586)
);

OA21x2_ASAP7_75t_L g587 ( 
.A1(n_560),
.A2(n_235),
.B(n_290),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_563),
.Y(n_588)
);

NOR2xp67_ASAP7_75t_SL g589 ( 
.A(n_470),
.B(n_211),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_537),
.A2(n_261),
.B1(n_264),
.B2(n_270),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_468),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_563),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_445),
.B(n_260),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_538),
.B(n_262),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_485),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_470),
.Y(n_596)
);

OR2x6_ASAP7_75t_L g597 ( 
.A(n_490),
.B(n_211),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_522),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_466),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_473),
.B(n_265),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_580),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_580),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_537),
.A2(n_214),
.B1(n_250),
.B2(n_247),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_L g604 ( 
.A1(n_543),
.A2(n_232),
.B1(n_222),
.B2(n_223),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_469),
.B(n_271),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_573),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_573),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_456),
.B(n_222),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_575),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_483),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_558),
.B(n_229),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_572),
.B(n_232),
.Y(n_612)
);

O2A1O1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_489),
.A2(n_461),
.B(n_464),
.C(n_448),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_505),
.B(n_467),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_489),
.A2(n_286),
.B1(n_273),
.B2(n_274),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_488),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_492),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_446),
.B(n_201),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_513),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_508),
.Y(n_620)
);

NOR2xp67_ASAP7_75t_L g621 ( 
.A(n_567),
.B(n_275),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_470),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_496),
.B(n_284),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_461),
.B(n_235),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_496),
.B(n_240),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_493),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_509),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_444),
.B(n_454),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_514),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_499),
.B(n_240),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_455),
.B(n_247),
.Y(n_631)
);

AND2x2_ASAP7_75t_SL g632 ( 
.A(n_459),
.B(n_250),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_524),
.B(n_263),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_526),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_575),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_443),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_482),
.B(n_204),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_453),
.A2(n_263),
.B1(n_387),
.B2(n_425),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_536),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_546),
.B(n_205),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_547),
.B(n_428),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_542),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_545),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_443),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_486),
.B(n_209),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_547),
.B(n_436),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_552),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_511),
.B(n_225),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_550),
.B(n_453),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_518),
.B(n_230),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_508),
.Y(n_651)
);

AND2x6_ASAP7_75t_SL g652 ( 
.A(n_501),
.B(n_348),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_550),
.B(n_436),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_478),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_510),
.B(n_348),
.Y(n_655)
);

AND2x4_ASAP7_75t_SL g656 ( 
.A(n_474),
.B(n_423),
.Y(n_656)
);

AND2x6_ASAP7_75t_SL g657 ( 
.A(n_551),
.B(n_351),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_539),
.A2(n_285),
.B1(n_277),
.B2(n_358),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_539),
.A2(n_285),
.B1(n_277),
.B2(n_358),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_484),
.B(n_360),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_533),
.B(n_277),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_447),
.B(n_241),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_460),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_576),
.B(n_553),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_559),
.B(n_245),
.Y(n_665)
);

BUFx6f_ASAP7_75t_SL g666 ( 
.A(n_474),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_503),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_525),
.B(n_252),
.Y(n_668)
);

AOI22x1_ASAP7_75t_L g669 ( 
.A1(n_539),
.A2(n_369),
.B1(n_368),
.B2(n_364),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_503),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_478),
.B(n_362),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_503),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_479),
.B(n_363),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_479),
.B(n_363),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_479),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_479),
.B(n_502),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_574),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_502),
.B(n_364),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_462),
.A2(n_405),
.B1(n_383),
.B2(n_382),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_535),
.B(n_259),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_502),
.B(n_369),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_459),
.A2(n_283),
.B1(n_267),
.B2(n_268),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_579),
.B(n_266),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_555),
.B(n_280),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_565),
.B(n_281),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_460),
.Y(n_686)
);

CKINVDCx11_ASAP7_75t_R g687 ( 
.A(n_474),
.Y(n_687)
);

INVx8_ASAP7_75t_L g688 ( 
.A(n_471),
.Y(n_688)
);

AOI221xp5_ASAP7_75t_L g689 ( 
.A1(n_506),
.A2(n_282),
.B1(n_329),
.B2(n_323),
.C(n_322),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_529),
.B(n_277),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_471),
.B(n_544),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_448),
.B(n_321),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_529),
.B(n_285),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_544),
.A2(n_459),
.B1(n_465),
.B2(n_561),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_544),
.B(n_90),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_465),
.A2(n_376),
.B1(n_285),
.B2(n_144),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_578),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_549),
.B(n_6),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_451),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_472),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_472),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_477),
.B(n_129),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_561),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_476),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_548),
.B(n_10),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_476),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_500),
.B(n_10),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_529),
.B(n_11),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_548),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_481),
.B(n_86),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_491),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_495),
.B(n_11),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_520),
.A2(n_84),
.B1(n_78),
.B2(n_77),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_497),
.B(n_13),
.Y(n_714)
);

AND2x6_ASAP7_75t_SL g715 ( 
.A(n_513),
.B(n_13),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_556),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_520),
.Y(n_717)
);

NAND2x1_ASAP7_75t_L g718 ( 
.A(n_463),
.B(n_75),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_520),
.B(n_15),
.Y(n_719)
);

BUFx5_ASAP7_75t_L g720 ( 
.A(n_557),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_491),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_564),
.Y(n_722)
);

AND2x2_ASAP7_75t_SL g723 ( 
.A(n_566),
.B(n_58),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_481),
.B(n_18),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_601),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_596),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_588),
.Y(n_727)
);

NOR2x1p5_ASAP7_75t_L g728 ( 
.A(n_619),
.B(n_523),
.Y(n_728)
);

O2A1O1Ixp5_ASAP7_75t_L g729 ( 
.A1(n_611),
.A2(n_517),
.B(n_515),
.C(n_519),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_691),
.A2(n_450),
.B(n_449),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_614),
.B(n_481),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_603),
.B(n_590),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_596),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_590),
.B(n_649),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_614),
.B(n_532),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_723),
.A2(n_504),
.B1(n_534),
.B2(n_498),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_596),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_676),
.A2(n_449),
.B(n_450),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_723),
.B(n_475),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_694),
.B(n_487),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_618),
.B(n_521),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_618),
.A2(n_528),
.B1(n_519),
.B2(n_517),
.Y(n_742)
);

NAND2x1p5_ASAP7_75t_L g743 ( 
.A(n_596),
.B(n_654),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_654),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_654),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_613),
.A2(n_449),
.B(n_450),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_669),
.A2(n_695),
.B(n_702),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_620),
.B(n_651),
.Y(n_748)
);

OA21x2_ASAP7_75t_L g749 ( 
.A1(n_694),
.A2(n_515),
.B(n_507),
.Y(n_749)
);

O2A1O1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_717),
.A2(n_568),
.B(n_577),
.C(n_530),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_588),
.Y(n_751)
);

BUFx8_ASAP7_75t_L g752 ( 
.A(n_666),
.Y(n_752)
);

AND3x2_ASAP7_75t_L g753 ( 
.A(n_705),
.B(n_21),
.C(n_22),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_648),
.A2(n_530),
.B(n_507),
.C(n_568),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_584),
.B(n_577),
.Y(n_755)
);

AO21x1_ASAP7_75t_L g756 ( 
.A1(n_612),
.A2(n_452),
.B(n_571),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_592),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_632),
.A2(n_452),
.B1(n_562),
.B2(n_554),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_622),
.A2(n_449),
.B(n_450),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_592),
.Y(n_760)
);

BUFx12f_ASAP7_75t_L g761 ( 
.A(n_687),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_598),
.B(n_463),
.Y(n_762)
);

AO21x1_ASAP7_75t_L g763 ( 
.A1(n_712),
.A2(n_570),
.B(n_569),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_656),
.Y(n_764)
);

NAND2x1p5_ASAP7_75t_L g765 ( 
.A(n_654),
.B(n_463),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_628),
.A2(n_516),
.B(n_570),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_688),
.A2(n_516),
.B(n_569),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_675),
.Y(n_768)
);

NOR3xp33_ASAP7_75t_L g769 ( 
.A(n_648),
.B(n_527),
.C(n_554),
.Y(n_769)
);

NOR2xp67_ASAP7_75t_L g770 ( 
.A(n_709),
.B(n_527),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_602),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_661),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_606),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_650),
.B(n_637),
.Y(n_774)
);

INVx5_ASAP7_75t_L g775 ( 
.A(n_675),
.Y(n_775)
);

AO21x1_ASAP7_75t_L g776 ( 
.A1(n_712),
.A2(n_541),
.B(n_531),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_650),
.B(n_562),
.Y(n_777)
);

CKINVDCx16_ASAP7_75t_R g778 ( 
.A(n_666),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_586),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_675),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_606),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_599),
.Y(n_782)
);

CKINVDCx6p67_ASAP7_75t_R g783 ( 
.A(n_597),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_680),
.B(n_554),
.Y(n_784)
);

AOI21x1_ASAP7_75t_L g785 ( 
.A1(n_641),
.A2(n_512),
.B(n_540),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_610),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_703),
.A2(n_512),
.B1(n_34),
.B2(n_35),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_SL g788 ( 
.A(n_656),
.B(n_52),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_604),
.A2(n_28),
.B(n_34),
.C(n_36),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_646),
.A2(n_37),
.B(n_38),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_581),
.B(n_38),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_581),
.B(n_39),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_699),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_655),
.B(n_40),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_660),
.B(n_637),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_607),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_703),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_797)
);

O2A1O1Ixp5_ASAP7_75t_L g798 ( 
.A1(n_605),
.A2(n_48),
.B(n_49),
.C(n_624),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_616),
.Y(n_799)
);

O2A1O1Ixp5_ASAP7_75t_L g800 ( 
.A1(n_608),
.A2(n_48),
.B(n_585),
.C(n_685),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_655),
.Y(n_801)
);

O2A1O1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_705),
.A2(n_582),
.B(n_714),
.C(n_696),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_607),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_583),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_645),
.B(n_667),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_645),
.B(n_593),
.Y(n_806)
);

AOI33xp33_ASAP7_75t_L g807 ( 
.A1(n_658),
.A2(n_659),
.A3(n_638),
.B1(n_707),
.B2(n_719),
.B3(n_689),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_670),
.B(n_672),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_586),
.Y(n_809)
);

AOI21x1_ASAP7_75t_L g810 ( 
.A1(n_653),
.A2(n_671),
.B(n_673),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_617),
.B(n_626),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_609),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_600),
.B(n_625),
.Y(n_813)
);

AOI21x1_ASAP7_75t_L g814 ( 
.A1(n_674),
.A2(n_681),
.B(n_678),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_627),
.B(n_629),
.Y(n_815)
);

AND2x2_ASAP7_75t_SL g816 ( 
.A(n_658),
.B(n_659),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_634),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_600),
.B(n_630),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_621),
.B(n_583),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_591),
.B(n_597),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_698),
.A2(n_683),
.B1(n_684),
.B2(n_668),
.Y(n_821)
);

AOI21x1_ASAP7_75t_L g822 ( 
.A1(n_631),
.A2(n_677),
.B(n_697),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_639),
.B(n_642),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_710),
.A2(n_686),
.B(n_700),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_633),
.B(n_623),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_635),
.A2(n_686),
.B(n_721),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_595),
.B(n_710),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_597),
.Y(n_828)
);

CKINVDCx11_ASAP7_75t_R g829 ( 
.A(n_652),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_698),
.A2(n_668),
.B(n_662),
.C(n_647),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_636),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_643),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_690),
.B(n_693),
.C(n_662),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_692),
.B(n_722),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_636),
.B(n_644),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_644),
.B(n_706),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_663),
.B(n_700),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_595),
.B(n_708),
.Y(n_838)
);

NOR2xp67_ASAP7_75t_L g839 ( 
.A(n_615),
.B(n_679),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_701),
.B(n_711),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_704),
.B(n_716),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_724),
.A2(n_665),
.B(n_682),
.C(n_640),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_587),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_718),
.A2(n_594),
.B(n_587),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_657),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_720),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_720),
.B(n_713),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_720),
.B(n_589),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_720),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_715),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_694),
.A2(n_465),
.B(n_459),
.Y(n_851)
);

BUFx2_ASAP7_75t_SL g852 ( 
.A(n_666),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_603),
.A2(n_590),
.B1(n_723),
.B2(n_703),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_603),
.B(n_590),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_614),
.B(n_543),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_723),
.A2(n_603),
.B1(n_590),
.B2(n_632),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_603),
.B(n_590),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_664),
.A2(n_676),
.B(n_669),
.Y(n_858)
);

O2A1O1Ixp5_ASAP7_75t_L g859 ( 
.A1(n_611),
.A2(n_543),
.B(n_612),
.C(n_561),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_603),
.B(n_590),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_603),
.B(n_590),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_603),
.B(n_590),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_603),
.B(n_458),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_584),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_694),
.A2(n_465),
.B(n_459),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_614),
.B(n_543),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_588),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_694),
.A2(n_465),
.B(n_459),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_596),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_588),
.Y(n_870)
);

BUFx8_ASAP7_75t_L g871 ( 
.A(n_666),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_717),
.A2(n_489),
.B(n_604),
.C(n_705),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_614),
.B(n_445),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_614),
.B(n_445),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_588),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_603),
.B(n_458),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_588),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_588),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_614),
.B(n_543),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_SL g880 ( 
.A(n_584),
.B(n_474),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_603),
.B(n_458),
.Y(n_881)
);

BUFx4f_ASAP7_75t_L g882 ( 
.A(n_656),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_664),
.A2(n_477),
.B(n_470),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_873),
.B(n_874),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_748),
.B(n_864),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_774),
.B(n_795),
.Y(n_886)
);

AOI21x1_ASAP7_75t_L g887 ( 
.A1(n_746),
.A2(n_731),
.B(n_785),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_853),
.A2(n_856),
.B(n_732),
.C(n_862),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_851),
.A2(n_868),
.B(n_865),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_779),
.B(n_809),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_851),
.A2(n_868),
.B(n_865),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_855),
.B(n_866),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_853),
.A2(n_854),
.B(n_857),
.C(n_732),
.Y(n_893)
);

AOI21xp33_ASAP7_75t_L g894 ( 
.A1(n_806),
.A2(n_802),
.B(n_879),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_735),
.B(n_741),
.Y(n_895)
);

OAI21x1_ASAP7_75t_L g896 ( 
.A1(n_824),
.A2(n_858),
.B(n_826),
.Y(n_896)
);

AOI21x1_ASAP7_75t_L g897 ( 
.A1(n_822),
.A2(n_844),
.B(n_784),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_859),
.A2(n_740),
.B(n_739),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_793),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_883),
.A2(n_775),
.B(n_777),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_755),
.Y(n_901)
);

NAND2x1p5_ASAP7_75t_L g902 ( 
.A(n_775),
.B(n_726),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_726),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_804),
.Y(n_904)
);

O2A1O1Ixp5_ASAP7_75t_L g905 ( 
.A1(n_763),
.A2(n_776),
.B(n_756),
.C(n_792),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_821),
.B(n_805),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_773),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_772),
.B(n_779),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_863),
.B(n_876),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_881),
.B(n_854),
.Y(n_910)
);

CKINVDCx8_ASAP7_75t_R g911 ( 
.A(n_852),
.Y(n_911)
);

AO31x2_ASAP7_75t_L g912 ( 
.A1(n_787),
.A2(n_830),
.A3(n_754),
.B(n_797),
.Y(n_912)
);

AOI21x1_ASAP7_75t_SL g913 ( 
.A1(n_847),
.A2(n_848),
.B(n_734),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_857),
.B(n_860),
.Y(n_914)
);

OA21x2_ASAP7_75t_L g915 ( 
.A1(n_747),
.A2(n_843),
.B(n_847),
.Y(n_915)
);

OAI21x1_ASAP7_75t_L g916 ( 
.A1(n_810),
.A2(n_814),
.B(n_766),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_726),
.Y(n_917)
);

INVx6_ASAP7_75t_L g918 ( 
.A(n_804),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_729),
.A2(n_742),
.B(n_734),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_804),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_860),
.B(n_861),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_839),
.A2(n_813),
.B1(n_818),
.B2(n_825),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_SL g923 ( 
.A1(n_833),
.A2(n_797),
.B(n_753),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_733),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_SL g925 ( 
.A1(n_787),
.A2(n_862),
.B(n_861),
.Y(n_925)
);

AOI211x1_ASAP7_75t_L g926 ( 
.A1(n_791),
.A2(n_815),
.B(n_811),
.C(n_823),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_738),
.A2(n_730),
.B(n_767),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_SL g928 ( 
.A1(n_789),
.A2(n_842),
.B(n_794),
.C(n_872),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_733),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_809),
.B(n_762),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_816),
.A2(n_827),
.B1(n_736),
.B2(n_834),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_781),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_782),
.B(n_786),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_828),
.Y(n_934)
);

OAI21x1_ASAP7_75t_L g935 ( 
.A1(n_835),
.A2(n_840),
.B(n_836),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_838),
.B(n_880),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_835),
.A2(n_836),
.B(n_837),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_807),
.A2(n_750),
.B(n_798),
.C(n_800),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_733),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_799),
.A2(n_817),
.B(n_832),
.C(n_790),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_841),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_846),
.A2(n_849),
.B(n_759),
.Y(n_942)
);

AND3x2_ASAP7_75t_L g943 ( 
.A(n_788),
.B(n_850),
.C(n_801),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_764),
.Y(n_944)
);

NAND2xp33_ASAP7_75t_SL g945 ( 
.A(n_737),
.B(n_869),
.Y(n_945)
);

AND3x4_ASAP7_75t_L g946 ( 
.A(n_770),
.B(n_829),
.C(n_769),
.Y(n_946)
);

OAI21xp33_ASAP7_75t_L g947 ( 
.A1(n_808),
.A2(n_845),
.B(n_838),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_838),
.B(n_820),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_SL g949 ( 
.A1(n_749),
.A2(n_827),
.B(n_768),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_820),
.B(n_882),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_820),
.B(n_882),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_758),
.A2(n_771),
.B(n_727),
.C(n_877),
.Y(n_952)
);

AO31x2_ASAP7_75t_L g953 ( 
.A1(n_796),
.A2(n_812),
.A3(n_803),
.B(n_831),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_783),
.B(n_728),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_765),
.A2(n_743),
.B(n_725),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_751),
.B(n_878),
.Y(n_956)
);

AOI21x1_ASAP7_75t_SL g957 ( 
.A1(n_749),
.A2(n_819),
.B(n_744),
.Y(n_957)
);

AO31x2_ASAP7_75t_L g958 ( 
.A1(n_757),
.A2(n_875),
.A3(n_870),
.B(n_867),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_760),
.B(n_737),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_737),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_745),
.A2(n_768),
.B(n_780),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_745),
.A2(n_768),
.B(n_780),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_745),
.A2(n_780),
.B(n_869),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_778),
.B(n_869),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_752),
.B(n_871),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_871),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_752),
.Y(n_967)
);

NAND2x1_ASAP7_75t_SL g968 ( 
.A(n_761),
.B(n_543),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_873),
.B(n_874),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_824),
.A2(n_858),
.B(n_785),
.Y(n_970)
);

OAI21x1_ASAP7_75t_L g971 ( 
.A1(n_858),
.A2(n_785),
.B(n_746),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_773),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_804),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_774),
.A2(n_859),
.B(n_740),
.Y(n_974)
);

O2A1O1Ixp5_ASAP7_75t_L g975 ( 
.A1(n_774),
.A2(n_741),
.B(n_776),
.C(n_763),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_873),
.B(n_874),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_841),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_873),
.B(n_874),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_824),
.A2(n_858),
.B(n_785),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_804),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_873),
.B(n_874),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_774),
.A2(n_874),
.B1(n_873),
.B2(n_853),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_824),
.A2(n_858),
.B(n_785),
.Y(n_983)
);

AO31x2_ASAP7_75t_L g984 ( 
.A1(n_763),
.A2(n_776),
.A3(n_756),
.B(n_853),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_841),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_873),
.B(n_874),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_856),
.A2(n_774),
.B1(n_853),
.B2(n_732),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_774),
.B(n_873),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_774),
.A2(n_874),
.B1(n_873),
.B2(n_853),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_774),
.A2(n_873),
.B(n_874),
.C(n_853),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_856),
.A2(n_774),
.B1(n_853),
.B2(n_732),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_873),
.B(n_874),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_824),
.A2(n_858),
.B(n_785),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_774),
.B(n_873),
.Y(n_994)
);

CKINVDCx20_ASAP7_75t_R g995 ( 
.A(n_778),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_873),
.B(n_874),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_824),
.A2(n_858),
.B(n_785),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_856),
.B(n_853),
.Y(n_998)
);

AO31x2_ASAP7_75t_L g999 ( 
.A1(n_763),
.A2(n_776),
.A3(n_756),
.B(n_853),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_841),
.Y(n_1000)
);

AO21x1_ASAP7_75t_L g1001 ( 
.A1(n_853),
.A2(n_774),
.B(n_802),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_774),
.B(n_873),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_774),
.B(n_873),
.Y(n_1003)
);

OAI21xp33_ASAP7_75t_L g1004 ( 
.A1(n_873),
.A2(n_874),
.B(n_774),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_774),
.B(n_873),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_774),
.A2(n_859),
.B(n_740),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_804),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_824),
.A2(n_858),
.B(n_785),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_774),
.A2(n_859),
.B(n_740),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_856),
.B(n_853),
.Y(n_1010)
);

OAI22x1_ASAP7_75t_L g1011 ( 
.A1(n_873),
.A2(n_874),
.B1(n_543),
.B2(n_774),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_SL g1012 ( 
.A(n_864),
.B(n_584),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_774),
.B(n_873),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_873),
.B(n_874),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_726),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_824),
.A2(n_858),
.B(n_785),
.Y(n_1016)
);

AO31x2_ASAP7_75t_L g1017 ( 
.A1(n_763),
.A2(n_776),
.A3(n_756),
.B(n_853),
.Y(n_1017)
);

O2A1O1Ixp5_ASAP7_75t_L g1018 ( 
.A1(n_774),
.A2(n_741),
.B(n_776),
.C(n_763),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_885),
.Y(n_1019)
);

INVx5_ASAP7_75t_L g1020 ( 
.A(n_903),
.Y(n_1020)
);

OR2x2_ASAP7_75t_SL g1021 ( 
.A(n_988),
.B(n_994),
.Y(n_1021)
);

AO31x2_ASAP7_75t_L g1022 ( 
.A1(n_1001),
.A2(n_987),
.A3(n_991),
.B(n_889),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_964),
.Y(n_1023)
);

AO32x1_ASAP7_75t_L g1024 ( 
.A1(n_931),
.A2(n_913),
.A3(n_941),
.B1(n_977),
.B2(n_1000),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_895),
.B(n_886),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_990),
.A2(n_989),
.B(n_982),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_976),
.B(n_978),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_990),
.A2(n_1004),
.B(n_1014),
.C(n_969),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_884),
.B(n_969),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_884),
.B(n_1014),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_981),
.B(n_986),
.Y(n_1031)
);

O2A1O1Ixp5_ASAP7_75t_L g1032 ( 
.A1(n_998),
.A2(n_1010),
.B(n_975),
.C(n_1018),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_995),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_992),
.B(n_996),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_907),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_953),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_904),
.B(n_920),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1002),
.B(n_1003),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_1005),
.B(n_1013),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_904),
.B(n_920),
.Y(n_1040)
);

CKINVDCx8_ASAP7_75t_R g1041 ( 
.A(n_934),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_892),
.B(n_901),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_901),
.B(n_1011),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_985),
.B(n_906),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_907),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_973),
.B(n_980),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_890),
.Y(n_1047)
);

OA21x2_ASAP7_75t_L g1048 ( 
.A1(n_896),
.A2(n_891),
.B(n_919),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_932),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_930),
.B(n_922),
.Y(n_1050)
);

INVx5_ASAP7_75t_L g1051 ( 
.A(n_903),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_L g1052 ( 
.A(n_888),
.B(n_940),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_995),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_944),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_SL g1055 ( 
.A1(n_974),
.A2(n_1006),
.B(n_1009),
.C(n_898),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_972),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_925),
.B(n_909),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_894),
.A2(n_928),
.B(n_1010),
.C(n_998),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_903),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1012),
.A2(n_923),
.B1(n_946),
.B2(n_947),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_908),
.B(n_936),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_944),
.Y(n_1062)
);

NAND2x1p5_ASAP7_75t_L g1063 ( 
.A(n_973),
.B(n_980),
.Y(n_1063)
);

INVx6_ASAP7_75t_L g1064 ( 
.A(n_918),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_958),
.Y(n_1065)
);

OA21x2_ASAP7_75t_L g1066 ( 
.A1(n_905),
.A2(n_971),
.B(n_1016),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_888),
.B(n_910),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_899),
.Y(n_1068)
);

NAND2x1p5_ASAP7_75t_L g1069 ( 
.A(n_1007),
.B(n_903),
.Y(n_1069)
);

INVxp67_ASAP7_75t_SL g1070 ( 
.A(n_902),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_971),
.A2(n_970),
.B(n_979),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_890),
.B(n_911),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_946),
.A2(n_950),
.B1(n_951),
.B2(n_890),
.Y(n_1073)
);

OR2x6_ASAP7_75t_L g1074 ( 
.A(n_948),
.B(n_967),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_SL g1075 ( 
.A(n_943),
.B(n_954),
.Y(n_1075)
);

OR2x6_ASAP7_75t_L g1076 ( 
.A(n_967),
.B(n_902),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_1007),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_943),
.B(n_960),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_960),
.B(n_939),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_893),
.A2(n_921),
.B1(n_914),
.B2(n_926),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_893),
.B(n_912),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_918),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_956),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_924),
.B(n_939),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_949),
.A2(n_900),
.B(n_928),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_940),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_959),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_968),
.B(n_938),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_966),
.Y(n_1089)
);

BUFx12f_ASAP7_75t_L g1090 ( 
.A(n_917),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_938),
.B(n_929),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_952),
.Y(n_1092)
);

O2A1O1Ixp5_ASAP7_75t_L g1093 ( 
.A1(n_975),
.A2(n_1018),
.B(n_905),
.C(n_887),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_924),
.A2(n_1015),
.B1(n_929),
.B2(n_945),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_935),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1015),
.B(n_912),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_952),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_965),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_942),
.A2(n_961),
.B(n_915),
.C(n_912),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_R g1100 ( 
.A(n_945),
.B(n_917),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_912),
.B(n_937),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_984),
.B(n_1017),
.Y(n_1102)
);

NAND3xp33_ASAP7_75t_L g1103 ( 
.A(n_915),
.B(n_917),
.C(n_913),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_962),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_963),
.Y(n_1105)
);

OR2x6_ASAP7_75t_L g1106 ( 
.A(n_955),
.B(n_916),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_915),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_984),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_984),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_983),
.A2(n_993),
.B1(n_1008),
.B2(n_997),
.Y(n_1110)
);

INVxp67_ASAP7_75t_L g1111 ( 
.A(n_897),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_984),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_927),
.B(n_957),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1017),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_999),
.B(n_1017),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_957),
.A2(n_999),
.B(n_1017),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_SL g1117 ( 
.A1(n_999),
.A2(n_853),
.B(n_1001),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_999),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_933),
.Y(n_1119)
);

INVx3_ASAP7_75t_SL g1120 ( 
.A(n_995),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_895),
.B(n_886),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_976),
.B(n_978),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_884),
.A2(n_774),
.B1(n_874),
.B2(n_873),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_895),
.A2(n_856),
.B1(n_853),
.B2(n_982),
.Y(n_1124)
);

INVx6_ASAP7_75t_L g1125 ( 
.A(n_918),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_995),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_976),
.B(n_978),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_903),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_895),
.B(n_886),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_976),
.B(n_978),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_922),
.B(n_774),
.Y(n_1131)
);

BUFx10_ASAP7_75t_L g1132 ( 
.A(n_943),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_895),
.B(n_886),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_933),
.Y(n_1134)
);

NOR2xp67_ASAP7_75t_L g1135 ( 
.A(n_922),
.B(n_793),
.Y(n_1135)
);

OR2x6_ASAP7_75t_L g1136 ( 
.A(n_964),
.B(n_853),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_904),
.B(n_920),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_903),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_895),
.B(n_886),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_895),
.A2(n_873),
.B(n_874),
.C(n_774),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_944),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_976),
.B(n_978),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_976),
.B(n_978),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_976),
.B(n_978),
.Y(n_1144)
);

INVx3_ASAP7_75t_SL g1145 ( 
.A(n_995),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_990),
.A2(n_774),
.B(n_874),
.C(n_873),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_990),
.A2(n_774),
.B(n_982),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_995),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_SL g1149 ( 
.A1(n_990),
.A2(n_853),
.B(n_851),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_885),
.Y(n_1150)
);

AO21x1_ASAP7_75t_L g1151 ( 
.A1(n_1124),
.A2(n_1131),
.B(n_1147),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1123),
.B(n_1038),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_1033),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1105),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1060),
.A2(n_1075),
.B1(n_1135),
.B2(n_1124),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1147),
.A2(n_1026),
.B1(n_1029),
.B2(n_1030),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_SL g1157 ( 
.A(n_1054),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1034),
.B(n_1031),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1045),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1027),
.B(n_1122),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1062),
.Y(n_1161)
);

CKINVDCx11_ASAP7_75t_R g1162 ( 
.A(n_1120),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1026),
.A2(n_1030),
.B1(n_1029),
.B2(n_1052),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_SL g1164 ( 
.A1(n_1075),
.A2(n_1088),
.B1(n_1132),
.B2(n_1038),
.Y(n_1164)
);

AO21x1_ASAP7_75t_L g1165 ( 
.A1(n_1140),
.A2(n_1058),
.B(n_1057),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_1053),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_SL g1167 ( 
.A1(n_1132),
.A2(n_1139),
.B1(n_1025),
.B2(n_1129),
.Y(n_1167)
);

BUFx8_ASAP7_75t_L g1168 ( 
.A(n_1150),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1140),
.B(n_1039),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_1068),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1141),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1020),
.Y(n_1172)
);

INVx8_ASAP7_75t_L g1173 ( 
.A(n_1051),
.Y(n_1173)
);

AO21x1_ASAP7_75t_L g1174 ( 
.A1(n_1058),
.A2(n_1057),
.B(n_1080),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1025),
.B(n_1121),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1049),
.Y(n_1176)
);

BUFx4_ASAP7_75t_R g1177 ( 
.A(n_1108),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1136),
.A2(n_1050),
.B1(n_1121),
.B2(n_1133),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_SL g1179 ( 
.A1(n_1129),
.A2(n_1133),
.B1(n_1139),
.B2(n_1061),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1056),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1136),
.A2(n_1117),
.B1(n_1043),
.B2(n_1119),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1019),
.Y(n_1182)
);

OAI22x1_ASAP7_75t_L g1183 ( 
.A1(n_1073),
.A2(n_1114),
.B1(n_1086),
.B2(n_1109),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_1042),
.Y(n_1184)
);

AO21x1_ASAP7_75t_SL g1185 ( 
.A1(n_1102),
.A2(n_1081),
.B(n_1067),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1134),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1136),
.A2(n_1044),
.B1(n_1142),
.B2(n_1144),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1127),
.B(n_1130),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1083),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1143),
.B(n_1023),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1110),
.A2(n_1099),
.B(n_1095),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1037),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1145),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1105),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_1077),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1051),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1044),
.A2(n_1118),
.B1(n_1092),
.B2(n_1097),
.Y(n_1197)
);

AO21x2_ASAP7_75t_L g1198 ( 
.A1(n_1103),
.A2(n_1055),
.B(n_1113),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1087),
.Y(n_1199)
);

BUFx4f_ASAP7_75t_SL g1200 ( 
.A(n_1090),
.Y(n_1200)
);

NAND2x1_ASAP7_75t_L g1201 ( 
.A(n_1104),
.B(n_1047),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1078),
.A2(n_1126),
.B1(n_1148),
.B2(n_1081),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1087),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1091),
.A2(n_1146),
.B1(n_1028),
.B2(n_1096),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1065),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1099),
.A2(n_1116),
.B(n_1093),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1074),
.A2(n_1078),
.B1(n_1149),
.B2(n_1072),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1047),
.Y(n_1208)
);

AOI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1106),
.A2(n_1101),
.B(n_1107),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1101),
.Y(n_1210)
);

CKINVDCx6p67_ASAP7_75t_R g1211 ( 
.A(n_1082),
.Y(n_1211)
);

INVx6_ASAP7_75t_L g1212 ( 
.A(n_1040),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_SL g1213 ( 
.A1(n_1098),
.A2(n_1100),
.B1(n_1074),
.B2(n_1021),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1074),
.A2(n_1048),
.B1(n_1115),
.B2(n_1112),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1079),
.Y(n_1215)
);

INVx4_ASAP7_75t_L g1216 ( 
.A(n_1040),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1069),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_SL g1218 ( 
.A1(n_1089),
.A2(n_1076),
.B1(n_1070),
.B2(n_1137),
.Y(n_1218)
);

INVx8_ASAP7_75t_L g1219 ( 
.A(n_1046),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1084),
.Y(n_1220)
);

OAI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1041),
.A2(n_1076),
.B1(n_1063),
.B2(n_1070),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1137),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1076),
.A2(n_1022),
.B1(n_1048),
.B2(n_1125),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1084),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1093),
.A2(n_1066),
.B(n_1032),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_SL g1226 ( 
.A1(n_1094),
.A2(n_1102),
.B(n_1111),
.Y(n_1226)
);

INVx6_ASAP7_75t_L g1227 ( 
.A(n_1064),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1138),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1138),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1059),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1066),
.A2(n_1032),
.B(n_1106),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1111),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1022),
.A2(n_1064),
.B1(n_1125),
.B2(n_1059),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1128),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1064),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1128),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1106),
.B(n_1125),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1024),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1024),
.B(n_1047),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1035),
.Y(n_1240)
);

OR2x6_ASAP7_75t_L g1241 ( 
.A(n_1149),
.B(n_1085),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1123),
.A2(n_988),
.B1(n_1002),
.B2(n_994),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1123),
.B(n_884),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1123),
.B(n_884),
.Y(n_1244)
);

BUFx12f_ASAP7_75t_L g1245 ( 
.A(n_1033),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1029),
.B(n_884),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1071),
.A2(n_971),
.B(n_970),
.Y(n_1247)
);

CKINVDCx9p33_ASAP7_75t_R g1248 ( 
.A(n_1021),
.Y(n_1248)
);

NAND2x1p5_ASAP7_75t_L g1249 ( 
.A(n_1020),
.B(n_1051),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1105),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1124),
.A2(n_774),
.B1(n_874),
.B2(n_873),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1036),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1124),
.A2(n_774),
.B1(n_874),
.B2(n_873),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_SL g1254 ( 
.A1(n_1124),
.A2(n_774),
.B1(n_874),
.B2(n_873),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1182),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1210),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1185),
.B(n_1197),
.Y(n_1257)
);

AND2x6_ASAP7_75t_L g1258 ( 
.A(n_1177),
.B(n_1172),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1205),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1195),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1237),
.B(n_1154),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1197),
.B(n_1156),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1232),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1232),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1156),
.B(n_1204),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1241),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1237),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1204),
.B(n_1214),
.Y(n_1268)
);

INVxp67_ASAP7_75t_R g1269 ( 
.A(n_1158),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1237),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1206),
.A2(n_1225),
.B(n_1238),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_1153),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1214),
.B(n_1163),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1163),
.B(n_1178),
.Y(n_1274)
);

OR2x6_ASAP7_75t_L g1275 ( 
.A(n_1241),
.B(n_1183),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1178),
.B(n_1181),
.Y(n_1276)
);

INVx4_ASAP7_75t_L g1277 ( 
.A(n_1177),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1181),
.B(n_1151),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1165),
.B(n_1187),
.Y(n_1279)
);

AO21x2_ASAP7_75t_L g1280 ( 
.A1(n_1191),
.A2(n_1209),
.B(n_1231),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1184),
.Y(n_1281)
);

INVxp67_ASAP7_75t_L g1282 ( 
.A(n_1199),
.Y(n_1282)
);

BUFx4f_ASAP7_75t_SL g1283 ( 
.A(n_1245),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1251),
.B(n_1253),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1187),
.B(n_1174),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1252),
.B(n_1239),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1247),
.A2(n_1241),
.B(n_1169),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1203),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1159),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1247),
.A2(n_1194),
.B(n_1250),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1176),
.Y(n_1291)
);

BUFx10_ASAP7_75t_L g1292 ( 
.A(n_1157),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1198),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1246),
.B(n_1175),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1183),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1180),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1239),
.B(n_1223),
.Y(n_1297)
);

INVx5_ASAP7_75t_SL g1298 ( 
.A(n_1248),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1179),
.B(n_1240),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1246),
.B(n_1152),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1254),
.B(n_1242),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1189),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1186),
.Y(n_1303)
);

INVxp33_ASAP7_75t_L g1304 ( 
.A(n_1160),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1201),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1233),
.A2(n_1207),
.B(n_1208),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1226),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1188),
.B(n_1155),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1243),
.B(n_1244),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1208),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1208),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1215),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1168),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1217),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1248),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1164),
.A2(n_1167),
.B1(n_1213),
.B2(n_1202),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1190),
.B(n_1224),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1301),
.A2(n_1265),
.B1(n_1262),
.B2(n_1268),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1284),
.A2(n_1221),
.B1(n_1170),
.B2(n_1193),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1259),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1286),
.B(n_1222),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1260),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1300),
.B(n_1218),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1292),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1304),
.B(n_1153),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1292),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1300),
.B(n_1309),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1295),
.B(n_1192),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1297),
.B(n_1230),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1301),
.A2(n_1162),
.B1(n_1168),
.B2(n_1245),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1297),
.B(n_1229),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1271),
.B(n_1236),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1271),
.B(n_1228),
.Y(n_1333)
);

OAI31xp33_ASAP7_75t_L g1334 ( 
.A1(n_1265),
.A2(n_1220),
.A3(n_1161),
.B(n_1171),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1290),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1275),
.B(n_1216),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1307),
.A2(n_1162),
.B1(n_1168),
.B2(n_1157),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1309),
.B(n_1234),
.Y(n_1338)
);

NOR2x1_ASAP7_75t_SL g1339 ( 
.A(n_1275),
.B(n_1172),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_1288),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1256),
.Y(n_1341)
);

AOI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1262),
.A2(n_1157),
.B1(n_1166),
.B2(n_1212),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1295),
.B(n_1235),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1263),
.Y(n_1344)
);

NAND2xp33_ASAP7_75t_R g1345 ( 
.A(n_1313),
.B(n_1200),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1293),
.B(n_1257),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1293),
.B(n_1161),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1266),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1293),
.B(n_1171),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1257),
.B(n_1196),
.Y(n_1350)
);

NOR2x1_ASAP7_75t_SL g1351 ( 
.A(n_1275),
.B(n_1172),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1263),
.Y(n_1352)
);

NOR3xp33_ASAP7_75t_L g1353 ( 
.A(n_1323),
.B(n_1307),
.C(n_1315),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1319),
.A2(n_1316),
.B1(n_1277),
.B2(n_1298),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1346),
.B(n_1278),
.Y(n_1355)
);

OAI221xp5_ASAP7_75t_L g1356 ( 
.A1(n_1319),
.A2(n_1315),
.B1(n_1294),
.B2(n_1281),
.C(n_1277),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1346),
.B(n_1273),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_L g1358 ( 
.A(n_1334),
.B(n_1279),
.C(n_1299),
.Y(n_1358)
);

OAI221xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1318),
.A2(n_1279),
.B1(n_1285),
.B2(n_1268),
.C(n_1276),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1327),
.B(n_1255),
.Y(n_1360)
);

OAI221xp5_ASAP7_75t_L g1361 ( 
.A1(n_1342),
.A2(n_1294),
.B1(n_1277),
.B2(n_1282),
.C(n_1299),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1329),
.B(n_1273),
.Y(n_1362)
);

OAI221xp5_ASAP7_75t_L g1363 ( 
.A1(n_1342),
.A2(n_1277),
.B1(n_1282),
.B2(n_1313),
.C(n_1308),
.Y(n_1363)
);

AND2x2_ASAP7_75t_SL g1364 ( 
.A(n_1336),
.B(n_1285),
.Y(n_1364)
);

OA211x2_ASAP7_75t_L g1365 ( 
.A1(n_1334),
.A2(n_1298),
.B(n_1258),
.C(n_1292),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_L g1366 ( 
.A(n_1318),
.B(n_1274),
.C(n_1276),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1327),
.B(n_1298),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1330),
.A2(n_1298),
.B1(n_1269),
.B2(n_1274),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_L g1369 ( 
.A(n_1323),
.B(n_1312),
.C(n_1308),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1322),
.B(n_1302),
.Y(n_1370)
);

OAI221xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1337),
.A2(n_1317),
.B1(n_1303),
.B2(n_1302),
.C(n_1312),
.Y(n_1371)
);

NAND3xp33_ASAP7_75t_L g1372 ( 
.A(n_1343),
.B(n_1305),
.C(n_1303),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1322),
.B(n_1340),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1329),
.B(n_1287),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1338),
.B(n_1264),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1329),
.B(n_1287),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1320),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1338),
.B(n_1264),
.Y(n_1378)
);

OAI21xp33_ASAP7_75t_L g1379 ( 
.A1(n_1325),
.A2(n_1317),
.B(n_1289),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1331),
.B(n_1280),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1347),
.A2(n_1306),
.B(n_1314),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1320),
.Y(n_1382)
);

NAND2xp33_ASAP7_75t_R g1383 ( 
.A(n_1350),
.B(n_1261),
.Y(n_1383)
);

NAND3xp33_ASAP7_75t_L g1384 ( 
.A(n_1347),
.B(n_1311),
.C(n_1310),
.Y(n_1384)
);

OA211x2_ASAP7_75t_L g1385 ( 
.A1(n_1339),
.A2(n_1298),
.B(n_1258),
.C(n_1292),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1331),
.B(n_1280),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1344),
.B(n_1291),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1344),
.B(n_1291),
.Y(n_1388)
);

NAND3xp33_ASAP7_75t_L g1389 ( 
.A(n_1349),
.B(n_1311),
.C(n_1310),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1352),
.B(n_1296),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1345),
.A2(n_1269),
.B1(n_1267),
.B2(n_1270),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1349),
.A2(n_1306),
.B(n_1314),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1377),
.Y(n_1393)
);

INVxp67_ASAP7_75t_SL g1394 ( 
.A(n_1372),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1377),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1382),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1382),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1387),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1357),
.B(n_1341),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1388),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1390),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1380),
.B(n_1352),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1364),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1380),
.B(n_1332),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1370),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1386),
.B(n_1332),
.Y(n_1406)
);

INVx2_ASAP7_75t_SL g1407 ( 
.A(n_1364),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1374),
.Y(n_1408)
);

INVxp67_ASAP7_75t_SL g1409 ( 
.A(n_1384),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1374),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1376),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1376),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1373),
.B(n_1332),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1389),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1355),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1362),
.B(n_1381),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1362),
.B(n_1333),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1375),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1392),
.B(n_1333),
.Y(n_1419)
);

NOR2xp67_ASAP7_75t_L g1420 ( 
.A(n_1369),
.B(n_1335),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1418),
.B(n_1353),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1397),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1418),
.B(n_1405),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1393),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1403),
.B(n_1339),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1418),
.B(n_1360),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1405),
.B(n_1398),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1398),
.B(n_1379),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1403),
.B(n_1351),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1404),
.B(n_1406),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1393),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1397),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1393),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1420),
.B(n_1391),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1397),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1397),
.Y(n_1436)
);

AND2x6_ASAP7_75t_SL g1437 ( 
.A(n_1399),
.B(n_1283),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1403),
.B(n_1351),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1395),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1414),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1404),
.B(n_1406),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1395),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1393),
.Y(n_1443)
);

INVx2_ASAP7_75t_SL g1444 ( 
.A(n_1393),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1407),
.B(n_1367),
.Y(n_1445)
);

CKINVDCx16_ASAP7_75t_R g1446 ( 
.A(n_1407),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_L g1447 ( 
.A(n_1394),
.B(n_1358),
.C(n_1366),
.Y(n_1447)
);

OAI21xp33_ASAP7_75t_L g1448 ( 
.A1(n_1414),
.A2(n_1359),
.B(n_1379),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1400),
.B(n_1378),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1396),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1396),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1407),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1415),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1400),
.B(n_1367),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1404),
.B(n_1321),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1406),
.B(n_1321),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1415),
.Y(n_1457)
);

NOR2x1p5_ASAP7_75t_SL g1458 ( 
.A(n_1411),
.B(n_1328),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1440),
.Y(n_1459)
);

INVxp67_ASAP7_75t_SL g1460 ( 
.A(n_1421),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1423),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1424),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1439),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1448),
.B(n_1414),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1455),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1437),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1439),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1447),
.B(n_1414),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1442),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1428),
.B(n_1394),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1442),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1446),
.B(n_1445),
.Y(n_1472)
);

NAND2x1_ASAP7_75t_SL g1473 ( 
.A(n_1445),
.B(n_1420),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1452),
.B(n_1408),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1450),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1424),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1452),
.B(n_1408),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1430),
.B(n_1409),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1430),
.B(n_1441),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1454),
.B(n_1409),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1455),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1434),
.B(n_1416),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1426),
.B(n_1416),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1425),
.B(n_1408),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1425),
.B(n_1416),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1450),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1451),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1429),
.B(n_1410),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1458),
.B(n_1411),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1449),
.B(n_1419),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1427),
.B(n_1419),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1429),
.B(n_1438),
.Y(n_1492)
);

INVxp33_ASAP7_75t_L g1493 ( 
.A(n_1438),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1456),
.A2(n_1354),
.B1(n_1365),
.B2(n_1361),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1441),
.B(n_1411),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1451),
.Y(n_1496)
);

NOR2xp67_ASAP7_75t_SL g1497 ( 
.A(n_1456),
.B(n_1356),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1453),
.B(n_1410),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1422),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1422),
.Y(n_1500)
);

NAND2x1_ASAP7_75t_L g1501 ( 
.A(n_1444),
.B(n_1419),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_SL g1502 ( 
.A(n_1466),
.B(n_1258),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1492),
.B(n_1458),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1463),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1463),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1489),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1460),
.B(n_1411),
.Y(n_1507)
);

OAI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1464),
.A2(n_1363),
.B1(n_1368),
.B2(n_1371),
.C(n_1401),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1467),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1472),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1472),
.B(n_1412),
.Y(n_1511)
);

AND2x6_ASAP7_75t_L g1512 ( 
.A(n_1474),
.B(n_1324),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1478),
.B(n_1453),
.Y(n_1513)
);

AND3x2_ASAP7_75t_L g1514 ( 
.A(n_1459),
.B(n_1457),
.C(n_1348),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1467),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1469),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1470),
.B(n_1412),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1489),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1489),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1473),
.A2(n_1433),
.B(n_1431),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1469),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1473),
.A2(n_1433),
.B(n_1431),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1492),
.B(n_1412),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1485),
.B(n_1412),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1471),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1468),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1495),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1482),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1495),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1497),
.Y(n_1530)
);

AOI22x1_ASAP7_75t_L g1531 ( 
.A1(n_1461),
.A2(n_1249),
.B1(n_1444),
.B2(n_1272),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1480),
.B(n_1401),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1484),
.B(n_1474),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1485),
.B(n_1417),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1477),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1484),
.B(n_1417),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1471),
.Y(n_1537)
);

OAI321xp33_ASAP7_75t_L g1538 ( 
.A1(n_1530),
.A2(n_1528),
.A3(n_1535),
.B1(n_1508),
.B2(n_1518),
.C(n_1506),
.Y(n_1538)
);

OAI21xp33_ASAP7_75t_L g1539 ( 
.A1(n_1526),
.A2(n_1494),
.B(n_1497),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1504),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1510),
.B(n_1493),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1510),
.B(n_1533),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1504),
.Y(n_1543)
);

AOI221xp5_ASAP7_75t_L g1544 ( 
.A1(n_1526),
.A2(n_1508),
.B1(n_1510),
.B2(n_1532),
.C(n_1535),
.Y(n_1544)
);

OAI221xp5_ASAP7_75t_L g1545 ( 
.A1(n_1510),
.A2(n_1478),
.B1(n_1501),
.B2(n_1481),
.C(n_1465),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1505),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1531),
.A2(n_1501),
.B1(n_1479),
.B2(n_1483),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1502),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1532),
.B(n_1479),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1533),
.B(n_1490),
.Y(n_1550)
);

OAI22x1_ASAP7_75t_L g1551 ( 
.A1(n_1531),
.A2(n_1477),
.B1(n_1488),
.B2(n_1486),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1505),
.Y(n_1552)
);

AOI21xp33_ASAP7_75t_L g1553 ( 
.A1(n_1506),
.A2(n_1486),
.B(n_1475),
.Y(n_1553)
);

AOI222xp33_ASAP7_75t_L g1554 ( 
.A1(n_1507),
.A2(n_1491),
.B1(n_1488),
.B2(n_1498),
.C1(n_1496),
.C2(n_1487),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1535),
.B(n_1475),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1509),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1533),
.B(n_1487),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_L g1558 ( 
.A(n_1514),
.B(n_1496),
.C(n_1499),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1507),
.B(n_1413),
.Y(n_1559)
);

O2A1O1Ixp33_ASAP7_75t_L g1560 ( 
.A1(n_1506),
.A2(n_1500),
.B(n_1499),
.C(n_1476),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1509),
.Y(n_1561)
);

OAI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1502),
.A2(n_1383),
.B1(n_1413),
.B2(n_1402),
.Y(n_1562)
);

NAND2x1_ASAP7_75t_L g1563 ( 
.A(n_1558),
.B(n_1533),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1542),
.B(n_1518),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1544),
.B(n_1518),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1539),
.A2(n_1512),
.B1(n_1511),
.B2(n_1503),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1540),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1541),
.B(n_1557),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1557),
.B(n_1519),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1543),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1548),
.B(n_1519),
.Y(n_1571)
);

OAI222xp33_ASAP7_75t_L g1572 ( 
.A1(n_1547),
.A2(n_1519),
.B1(n_1503),
.B2(n_1517),
.C1(n_1511),
.C2(n_1529),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1539),
.B(n_1554),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1550),
.B(n_1536),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1546),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1552),
.B(n_1556),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1549),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1561),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1555),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1560),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1538),
.B(n_1166),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1563),
.A2(n_1558),
.B(n_1551),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1563),
.A2(n_1545),
.B(n_1553),
.C(n_1562),
.Y(n_1583)
);

OAI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1573),
.A2(n_1559),
.B1(n_1517),
.B2(n_1503),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1581),
.A2(n_1529),
.B(n_1527),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1565),
.A2(n_1529),
.B(n_1527),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1572),
.A2(n_1522),
.B(n_1520),
.Y(n_1587)
);

AOI211xp5_ASAP7_75t_L g1588 ( 
.A1(n_1580),
.A2(n_1577),
.B(n_1568),
.C(n_1571),
.Y(n_1588)
);

AOI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1580),
.A2(n_1527),
.B1(n_1521),
.B2(n_1516),
.C(n_1537),
.Y(n_1589)
);

NAND4xp75_ASAP7_75t_L g1590 ( 
.A(n_1571),
.B(n_1537),
.C(n_1515),
.D(n_1521),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1579),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1569),
.A2(n_1516),
.B(n_1515),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1588),
.B(n_1564),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1591),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_L g1595 ( 
.A(n_1582),
.B(n_1566),
.C(n_1564),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1583),
.A2(n_1576),
.B(n_1579),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_L g1597 ( 
.A(n_1589),
.B(n_1586),
.C(n_1587),
.Y(n_1597)
);

NOR2x1_ASAP7_75t_L g1598 ( 
.A(n_1590),
.B(n_1567),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1592),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1585),
.Y(n_1600)
);

NOR2x1_ASAP7_75t_L g1601 ( 
.A(n_1584),
.B(n_1567),
.Y(n_1601)
);

AO22x1_ASAP7_75t_L g1602 ( 
.A1(n_1587),
.A2(n_1578),
.B1(n_1575),
.B2(n_1570),
.Y(n_1602)
);

NAND3xp33_ASAP7_75t_L g1603 ( 
.A(n_1597),
.B(n_1601),
.C(n_1598),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1594),
.B(n_1503),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1602),
.A2(n_1574),
.B(n_1525),
.Y(n_1605)
);

OAI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1596),
.A2(n_1522),
.B(n_1520),
.Y(n_1606)
);

OAI221xp5_ASAP7_75t_L g1607 ( 
.A1(n_1595),
.A2(n_1525),
.B1(n_1513),
.B2(n_1524),
.C(n_1534),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1600),
.B(n_1513),
.Y(n_1608)
);

OAI211xp5_ASAP7_75t_SL g1609 ( 
.A1(n_1593),
.A2(n_1500),
.B(n_1476),
.C(n_1462),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1604),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1603),
.A2(n_1599),
.B1(n_1512),
.B2(n_1536),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1608),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1607),
.B(n_1534),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1605),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1606),
.A2(n_1609),
.B1(n_1512),
.B2(n_1523),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_L g1616 ( 
.A(n_1603),
.B(n_1462),
.Y(n_1616)
);

OR2x6_ASAP7_75t_L g1617 ( 
.A(n_1610),
.B(n_1227),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1611),
.A2(n_1512),
.B1(n_1524),
.B2(n_1523),
.Y(n_1618)
);

NAND4xp75_ASAP7_75t_L g1619 ( 
.A(n_1616),
.B(n_1365),
.C(n_1385),
.D(n_1498),
.Y(n_1619)
);

INVxp33_ASAP7_75t_SL g1620 ( 
.A(n_1612),
.Y(n_1620)
);

NOR2x1_ASAP7_75t_L g1621 ( 
.A(n_1614),
.B(n_1443),
.Y(n_1621)
);

NOR2xp67_ASAP7_75t_L g1622 ( 
.A(n_1618),
.B(n_1615),
.Y(n_1622)
);

AO22x2_ASAP7_75t_L g1623 ( 
.A1(n_1619),
.A2(n_1613),
.B1(n_1443),
.B2(n_1432),
.Y(n_1623)
);

NOR3xp33_ASAP7_75t_L g1624 ( 
.A(n_1620),
.B(n_1326),
.C(n_1324),
.Y(n_1624)
);

OAI22x1_ASAP7_75t_L g1625 ( 
.A1(n_1622),
.A2(n_1621),
.B1(n_1617),
.B2(n_1512),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1625),
.B(n_1624),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1626),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1626),
.B(n_1623),
.Y(n_1628)
);

NAND2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1627),
.B(n_1211),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1628),
.B(n_1512),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1630),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1629),
.A2(n_1211),
.B1(n_1457),
.B2(n_1227),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1631),
.A2(n_1512),
.B(n_1435),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1633),
.A2(n_1632),
.B1(n_1512),
.B2(n_1227),
.Y(n_1634)
);

OAI221xp5_ASAP7_75t_R g1635 ( 
.A1(n_1634),
.A2(n_1173),
.B1(n_1219),
.B2(n_1385),
.C(n_1436),
.Y(n_1635)
);

AOI211xp5_ASAP7_75t_L g1636 ( 
.A1(n_1635),
.A2(n_1324),
.B(n_1326),
.C(n_1436),
.Y(n_1636)
);


endmodule