module fake_jpeg_22337_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_34),
.Y(n_49)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_16),
.Y(n_56)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_43),
.Y(n_68)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_28),
.B1(n_29),
.B2(n_22),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_51),
.B1(n_28),
.B2(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_52),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_28),
.B1(n_23),
.B2(n_30),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_54),
.Y(n_76)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_57),
.B(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_63),
.B(n_69),
.Y(n_104)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_66),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_71),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_73),
.Y(n_90)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

BUFx16f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_51),
.C(n_34),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_39),
.C(n_34),
.Y(n_110)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_44),
.B(n_32),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_87),
.B(n_79),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_86),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_45),
.B(n_35),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_54),
.B1(n_55),
.B2(n_25),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_41),
.B1(n_33),
.B2(n_37),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_30),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_66),
.B(n_40),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_35),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_100),
.Y(n_134)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_86),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_64),
.C(n_25),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_39),
.B1(n_30),
.B2(n_41),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_115),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_107),
.B1(n_98),
.B2(n_103),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_76),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_1),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_121),
.A2(n_96),
.B(n_20),
.Y(n_141)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_105),
.B1(n_109),
.B2(n_85),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_33),
.B1(n_37),
.B2(n_58),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_40),
.B1(n_65),
.B2(n_97),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_128),
.C(n_131),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_129),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_78),
.C(n_64),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_134),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_38),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_111),
.A2(n_37),
.B1(n_50),
.B2(n_45),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_137),
.B1(n_75),
.B2(n_77),
.Y(n_147)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_37),
.B1(n_40),
.B2(n_82),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_146),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_137),
.B(n_132),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_96),
.Y(n_152)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_101),
.C(n_102),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_155),
.C(n_159),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_83),
.B(n_25),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_20),
.B1(n_16),
.B2(n_24),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_158),
.A2(n_122),
.B1(n_118),
.B2(n_120),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_113),
.A2(n_136),
.B(n_128),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_90),
.C(n_80),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_163),
.C(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_118),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_121),
.A2(n_90),
.B(n_91),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_72),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_177),
.B1(n_178),
.B2(n_182),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_169),
.B(n_170),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_172),
.B(n_174),
.Y(n_197)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_72),
.Y(n_175)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_135),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_116),
.B1(n_20),
.B2(n_24),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_186),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_116),
.B1(n_24),
.B2(n_16),
.Y(n_182)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_2),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_184),
.B(n_189),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_18),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_17),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_11),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_27),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_71),
.C(n_27),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_140),
.C(n_163),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_191),
.A2(n_202),
.B(n_205),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_194),
.C(n_211),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_153),
.C(n_159),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_203),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_171),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_213),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_147),
.B(n_146),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_139),
.B1(n_144),
.B2(n_161),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_190),
.B1(n_177),
.B2(n_189),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_148),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_209),
.A2(n_181),
.B(n_179),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_148),
.Y(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_71),
.C(n_17),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_12),
.Y(n_228)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_209),
.B(n_183),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_230),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_226),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_173),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_208),
.B(n_171),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_228),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_166),
.B1(n_21),
.B2(n_19),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_232),
.B1(n_234),
.B2(n_198),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_209),
.B(n_21),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_202),
.B(n_12),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_233),
.Y(n_239)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_194),
.C(n_192),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_246),
.C(n_248),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_220),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_238),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_191),
.B1(n_203),
.B2(n_204),
.Y(n_240)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_240),
.Y(n_270)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_192),
.C(n_193),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_207),
.C(n_200),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_226),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_251),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_220),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_250),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_211),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_216),
.A2(n_200),
.B1(n_208),
.B2(n_213),
.Y(n_252)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_212),
.C(n_18),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_225),
.C(n_21),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_218),
.Y(n_255)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_241),
.A2(n_215),
.B(n_218),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_8),
.B(n_3),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_242),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_260),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_215),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_224),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_269),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_254),
.C(n_244),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_2),
.C(n_21),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_255),
.C(n_248),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_19),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_19),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_236),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_274),
.B(n_284),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_243),
.B1(n_251),
.B2(n_19),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_258),
.B1(n_265),
.B2(n_267),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_243),
.C(n_3),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_281),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_283),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_15),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_15),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_15),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_10),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_8),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_264),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_288),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_273),
.A2(n_268),
.B(n_256),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_266),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_292),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_295),
.Y(n_301)
);

NOR3xp33_ASAP7_75t_SL g297 ( 
.A(n_296),
.B(n_283),
.C(n_277),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_299),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_272),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_291),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_279),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_8),
.B(n_4),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g309 ( 
.A1(n_302),
.A2(n_303),
.A3(n_5),
.B1(n_6),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_4),
.B(n_5),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_5),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_290),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_308),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_309),
.A2(n_311),
.B(n_301),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_6),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_310),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_13),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_307),
.B(n_301),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_314),
.C(n_313),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_13),
.C(n_14),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_14),
.C(n_2),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_2),
.Y(n_320)
);


endmodule