module fake_jpeg_999_n_142 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_142);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_49),
.Y(n_68)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_62),
.B1(n_69),
.B2(n_58),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_42),
.B1(n_49),
.B2(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_70),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_44),
.B1(n_41),
.B2(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_51),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_58),
.B1(n_55),
.B2(n_57),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_40),
.B1(n_20),
.B2(n_21),
.Y(n_92)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_76),
.Y(n_95)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_77),
.B(n_82),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_50),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_80),
.Y(n_97)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_83),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_45),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_55),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_40),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_84),
.A2(n_67),
.B1(n_53),
.B2(n_45),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_87),
.B1(n_94),
.B2(n_14),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_53),
.B1(n_43),
.B2(n_40),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_30),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_73),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_18),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_96),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_15),
.B1(n_37),
.B2(n_36),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_1),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_105),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_79),
.B1(n_72),
.B2(n_23),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_104),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_88),
.B1(n_89),
.B2(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_108),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_1),
.B(n_2),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_112),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_2),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_10),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_3),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_9),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_27),
.B(n_35),
.C(n_34),
.D(n_32),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_24),
.B(n_31),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

OAI31xp33_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_125),
.A3(n_112),
.B(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_8),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_111),
.C(n_115),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_129),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_116),
.B1(n_117),
.B2(n_130),
.Y(n_135)
);

NOR2xp67_ASAP7_75t_SL g137 ( 
.A(n_135),
.B(n_117),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_133),
.B(n_130),
.C(n_124),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_123),
.B(n_118),
.C(n_136),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_121),
.B(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_25),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_29),
.Y(n_142)
);


endmodule