module fake_jpeg_1398_n_439 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_439);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_439;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_54),
.Y(n_100)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_49),
.Y(n_126)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_50),
.Y(n_140)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_52),
.Y(n_141)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_6),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_58),
.B(n_62),
.Y(n_151)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_15),
.B(n_6),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_18),
.B(n_24),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_64),
.B(n_66),
.Y(n_152)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_18),
.B(n_6),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_7),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_69),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_16),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_78),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_31),
.B(n_7),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_83),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_37),
.B(n_7),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_86),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_92),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_31),
.B(n_14),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_91),
.B(n_98),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_17),
.B(n_5),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_25),
.Y(n_125)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_95),
.Y(n_127)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_97),
.Y(n_142)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_105),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_68),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_74),
.A2(n_44),
.B1(n_32),
.B2(n_28),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_110),
.A2(n_113),
.B1(n_114),
.B2(n_134),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_49),
.A2(n_28),
.B1(n_27),
.B2(n_20),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_112),
.A2(n_118),
.B1(n_139),
.B2(n_27),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_44),
.B1(n_32),
.B2(n_36),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_67),
.A2(n_44),
.B1(n_19),
.B2(n_40),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_50),
.A2(n_27),
.B1(n_43),
.B2(n_38),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_44),
.B1(n_17),
.B2(n_19),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_119),
.A2(n_131),
.B1(n_34),
.B2(n_27),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_55),
.B(n_45),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_0),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_25),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_87),
.A2(n_40),
.B1(n_26),
.B2(n_88),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_92),
.A2(n_83),
.B1(n_95),
.B2(n_26),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_43),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_51),
.A2(n_27),
.B1(n_38),
.B2(n_36),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_96),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_143),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_61),
.B(n_77),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_144),
.B(n_149),
.Y(n_191)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_63),
.B(n_45),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_159),
.Y(n_234)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_104),
.A2(n_98),
.B1(n_94),
.B2(n_65),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_166),
.A2(n_183),
.B1(n_188),
.B2(n_203),
.Y(n_209)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_167),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_168),
.A2(n_153),
.B1(n_145),
.B2(n_117),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_104),
.A2(n_150),
.B1(n_151),
.B2(n_100),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_170),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_220)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_113),
.A2(n_34),
.B1(n_90),
.B2(n_60),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_120),
.A2(n_56),
.B1(n_53),
.B2(n_81),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_179),
.B(n_182),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_101),
.A2(n_34),
.B1(n_30),
.B2(n_9),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_104),
.A2(n_34),
.B1(n_30),
.B2(n_2),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_178),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_R g179 ( 
.A(n_124),
.B(n_30),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_180),
.B(n_196),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_181),
.A2(n_185),
.B1(n_186),
.B2(n_190),
.Y(n_228)
);

NAND2x1_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_108),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_109),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_192),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_111),
.A2(n_5),
.B1(n_11),
.B2(n_10),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_110),
.A2(n_4),
.B1(n_13),
.B2(n_3),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_109),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_108),
.B(n_0),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_193),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_127),
.A2(n_4),
.B1(n_13),
.B2(n_1),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g192 ( 
.A(n_140),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_120),
.B(n_4),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_123),
.A2(n_13),
.B1(n_141),
.B2(n_126),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_194),
.A2(n_187),
.B1(n_161),
.B2(n_202),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_152),
.B(n_141),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_198),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_108),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_123),
.B(n_146),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_199),
.B(n_201),
.Y(n_231)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_109),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_127),
.A2(n_157),
.B1(n_107),
.B2(n_156),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_107),
.A2(n_158),
.B1(n_157),
.B2(n_156),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_103),
.B1(n_155),
.B2(n_133),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_127),
.B(n_99),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_136),
.B(n_147),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_140),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_132),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_158),
.B1(n_153),
.B2(n_145),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_207),
.A2(n_216),
.B1(n_218),
.B2(n_233),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_211),
.A2(n_204),
.B1(n_181),
.B2(n_192),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_155),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_226),
.C(n_235),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_117),
.B1(n_99),
.B2(n_128),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_189),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_223),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_103),
.B(n_132),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_221),
.A2(n_243),
.B(n_175),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_148),
.B(n_147),
.C(n_136),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_222),
.B(n_175),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_193),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_116),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_229),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_170),
.B(n_116),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_133),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_237),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_177),
.A2(n_137),
.B1(n_154),
.B2(n_135),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_232),
.A2(n_192),
.B1(n_205),
.B2(n_200),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_164),
.A2(n_137),
.B1(n_130),
.B2(n_154),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_184),
.A2(n_121),
.B1(n_135),
.B2(n_197),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_241),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_206),
.A2(n_121),
.B(n_182),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_160),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_244),
.B(n_251),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_210),
.A2(n_191),
.B1(n_182),
.B2(n_199),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_260),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_214),
.Y(n_285)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_247),
.Y(n_297)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_250),
.A2(n_265),
.B1(n_207),
.B2(n_216),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_171),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_252),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_229),
.B(n_166),
.CI(n_191),
.CON(n_253),
.SN(n_253)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_253),
.B(n_257),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_215),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_258),
.Y(n_284)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_256),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_213),
.B(n_187),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_213),
.B(n_169),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_210),
.A2(n_161),
.B1(n_205),
.B2(n_175),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_225),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_266),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_159),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_269),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_224),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_267),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_268),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_201),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_273),
.A2(n_268),
.B1(n_248),
.B2(n_271),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_271),
.A2(n_210),
.B1(n_209),
.B2(n_242),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_277),
.A2(n_278),
.B1(n_296),
.B2(n_260),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_271),
.A2(n_209),
.B1(n_211),
.B2(n_221),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_214),
.C(n_219),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_285),
.C(n_295),
.Y(n_317)
);

AOI32xp33_ASAP7_75t_L g281 ( 
.A1(n_270),
.A2(n_239),
.A3(n_221),
.B1(n_237),
.B2(n_243),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_243),
.B(n_222),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_222),
.B(n_241),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_294),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_272),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_291),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_254),
.B(n_231),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_246),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_248),
.A2(n_209),
.B1(n_220),
.B2(n_232),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_297),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_301),
.Y(n_344)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_300),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_287),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_255),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_303),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_266),
.Y(n_304)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_305),
.A2(n_320),
.B1(n_277),
.B2(n_278),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_245),
.Y(n_306)
);

XNOR2x1_ASAP7_75t_L g335 ( 
.A(n_306),
.B(n_314),
.Y(n_335)
);

A2O1A1O1Ixp25_ASAP7_75t_L g307 ( 
.A1(n_276),
.A2(n_251),
.B(n_262),
.C(n_223),
.D(n_212),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_307),
.A2(n_284),
.B(n_294),
.Y(n_327)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_308),
.Y(n_345)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_309),
.Y(n_330)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_318),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_244),
.B1(n_256),
.B2(n_259),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_313),
.A2(n_290),
.B1(n_286),
.B2(n_298),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_258),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_257),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_315),
.B(n_316),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_223),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_297),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_319),
.A2(n_274),
.B1(n_283),
.B2(n_279),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_273),
.A2(n_271),
.B1(n_248),
.B2(n_262),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_219),
.C(n_239),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_321),
.B(n_298),
.Y(n_346)
);

OAI21xp33_ASAP7_75t_SL g323 ( 
.A1(n_302),
.A2(n_289),
.B(n_276),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_327),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_324),
.A2(n_328),
.B1(n_340),
.B2(n_343),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_284),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_325),
.A2(n_329),
.B1(n_331),
.B2(n_332),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_302),
.A2(n_279),
.B(n_274),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_326),
.A2(n_334),
.B(n_341),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_322),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_300),
.B(n_286),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_312),
.A2(n_279),
.B(n_281),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_304),
.B(n_290),
.Y(n_337)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_337),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_319),
.A2(n_292),
.B1(n_263),
.B2(n_291),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_310),
.A2(n_292),
.B(n_293),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_305),
.A2(n_207),
.B1(n_265),
.B2(n_216),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g358 ( 
.A(n_346),
.B(n_307),
.C(n_282),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_317),
.C(n_316),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_348),
.C(n_353),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_317),
.C(n_306),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_327),
.B(n_314),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_349),
.B(n_358),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_332),
.A2(n_310),
.B1(n_309),
.B2(n_311),
.Y(n_352)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_352),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_346),
.B(n_321),
.C(n_303),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_320),
.C(n_212),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_355),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_261),
.C(n_226),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_345),
.Y(n_356)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_356),
.Y(n_371)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_330),
.Y(n_357)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_357),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_269),
.C(n_238),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_359),
.B(n_365),
.Y(n_368)
);

XNOR2x2_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_253),
.Y(n_363)
);

AO21x1_ASAP7_75t_L g378 ( 
.A1(n_363),
.A2(n_326),
.B(n_341),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_328),
.A2(n_253),
.B1(n_297),
.B2(n_231),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_336),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_238),
.C(n_252),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_249),
.C(n_227),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_366),
.B(n_367),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_227),
.C(n_264),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_360),
.A2(n_340),
.B1(n_324),
.B2(n_337),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_373),
.A2(n_375),
.B1(n_377),
.B2(n_382),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_350),
.A2(n_361),
.B1(n_362),
.B2(n_351),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_365),
.A2(n_336),
.B1(n_343),
.B2(n_325),
.Y(n_377)
);

OAI221xp5_ASAP7_75t_L g384 ( 
.A1(n_378),
.A2(n_363),
.B1(n_358),
.B2(n_349),
.C(n_329),
.Y(n_384)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_357),
.Y(n_379)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_367),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_331),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_344),
.Y(n_383)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_383),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_384),
.A2(n_382),
.B1(n_390),
.B2(n_378),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_347),
.C(n_353),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_385),
.B(n_388),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_383),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_386),
.B(n_387),
.Y(n_400)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_348),
.C(n_354),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_381),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_391),
.B(n_392),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_359),
.C(n_355),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_370),
.A2(n_330),
.B1(n_333),
.B2(n_345),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_393),
.A2(n_373),
.B(n_374),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_394),
.A2(n_396),
.B(n_397),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_333),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_371),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_330),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_372),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_402),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_370),
.C(n_377),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_405),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_376),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_404),
.B(n_408),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_379),
.C(n_376),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_407),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_387),
.A2(n_371),
.B(n_272),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_409),
.A2(n_232),
.B(n_167),
.Y(n_417)
);

AOI322xp5_ASAP7_75t_L g410 ( 
.A1(n_400),
.A2(n_389),
.A3(n_388),
.B1(n_272),
.B2(n_253),
.C1(n_217),
.C2(n_247),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_410),
.A2(n_419),
.B(n_162),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_247),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_414),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_407),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_401),
.A2(n_250),
.B1(n_220),
.B2(n_228),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_416),
.A2(n_218),
.B1(n_228),
.B2(n_178),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_417),
.B(n_250),
.Y(n_420)
);

AOI322xp5_ASAP7_75t_L g419 ( 
.A1(n_398),
.A2(n_408),
.A3(n_402),
.B1(n_405),
.B2(n_399),
.C1(n_217),
.C2(n_167),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_422),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_233),
.C(n_172),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_418),
.A2(n_162),
.B(n_233),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_423),
.A2(n_426),
.B(n_162),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_424),
.A2(n_425),
.B1(n_427),
.B2(n_203),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_415),
.B(n_165),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_178),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_418),
.C(n_411),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_429),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_427),
.B(n_411),
.C(n_416),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_430),
.A2(n_420),
.B(n_218),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_431),
.B(n_175),
.C(n_188),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_433),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_434),
.A2(n_432),
.B(n_183),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_435),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_438),
.B(n_436),
.Y(n_439)
);


endmodule