module real_jpeg_30453_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_0),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_0),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_0),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_1),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_2),
.A2(n_118),
.B1(n_122),
.B2(n_125),
.Y(n_117)
);

INVx2_ASAP7_75t_R g125 ( 
.A(n_2),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_2),
.A2(n_125),
.B1(n_293),
.B2(n_296),
.Y(n_292)
);

AO22x1_ASAP7_75t_L g357 ( 
.A1(n_2),
.A2(n_125),
.B1(n_358),
.B2(n_361),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_3),
.A2(n_85),
.B1(n_87),
.B2(n_92),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_3),
.A2(n_92),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_3),
.A2(n_92),
.B1(n_272),
.B2(n_274),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_3),
.A2(n_92),
.B1(n_326),
.B2(n_331),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_4),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_5),
.Y(n_100)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_5),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_6),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_7),
.A2(n_62),
.B1(n_63),
.B2(n_67),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_8),
.Y(n_109)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_8),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_8),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_8),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_9),
.A2(n_221),
.B1(n_223),
.B2(n_225),
.Y(n_220)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_9),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_9),
.A2(n_225),
.B1(n_233),
.B2(n_236),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_9),
.A2(n_225),
.B1(n_317),
.B2(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_11),
.A2(n_200),
.B1(n_205),
.B2(n_209),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_11),
.A2(n_209),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_12),
.Y(n_182)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_12),
.Y(n_192)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_12),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_13),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_14),
.A2(n_131),
.B1(n_136),
.B2(n_137),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_14),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_14),
.A2(n_136),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_15),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_15),
.A2(n_48),
.B(n_156),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_L g239 ( 
.A1(n_15),
.A2(n_101),
.A3(n_240),
.B1(n_242),
.B2(n_247),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_15),
.A2(n_54),
.B1(n_271),
.B2(n_277),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_15),
.B(n_127),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_15),
.A2(n_143),
.B1(n_377),
.B2(n_379),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_263),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_261),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_226),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_19),
.B(n_226),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_152),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_52),
.B1(n_80),
.B2(n_81),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.A3(n_32),
.B1(n_39),
.B2(n_47),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_25),
.A2(n_146),
.B1(n_148),
.B2(n_151),
.Y(n_145)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_26),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_26),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_26),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_31),
.Y(n_151)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_36),
.Y(n_158)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_36),
.Y(n_162)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_46),
.Y(n_150)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_61),
.B1(n_68),
.B2(n_71),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_53),
.A2(n_61),
.B1(n_130),
.B2(n_140),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g251 ( 
.A1(n_53),
.A2(n_130),
.B1(n_252),
.B2(n_255),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_53),
.A2(n_285),
.B1(n_341),
.B2(n_344),
.Y(n_340)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_54),
.A2(n_271),
.B1(n_292),
.B2(n_298),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_54),
.A2(n_342),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_57),
.Y(n_254)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

BUFx2_ASAP7_75t_SL g289 ( 
.A(n_59),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_60),
.Y(n_276)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_65),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_65),
.Y(n_295)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_66),
.Y(n_307)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_66),
.Y(n_320)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_76),
.Y(n_194)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

BUFx2_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_128),
.C(n_142),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_83),
.B(n_229),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_93),
.B1(n_117),
.B2(n_126),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_84),
.A2(n_93),
.B1(n_126),
.B2(n_376),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_93),
.A2(n_117),
.B1(n_126),
.B2(n_220),
.Y(n_219)
);

AO21x2_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_101),
.B(n_107),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_103),
.Y(n_224)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_103),
.Y(n_378)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B1(n_112),
.B2(n_114),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_108),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_109),
.Y(n_330)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_109),
.Y(n_360)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_124),
.Y(n_222)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2x1_ASAP7_75t_L g229 ( 
.A(n_129),
.B(n_142),
.Y(n_229)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_139),
.Y(n_257)
);

BUFx4f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp67_ASAP7_75t_R g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_143),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_143),
.B(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_143),
.B(n_210),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_143),
.B(n_314),
.Y(n_313)
);

OAI21xp33_ASAP7_75t_SL g335 ( 
.A1(n_143),
.A2(n_313),
.B(n_336),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_155),
.B1(n_159),
.B2(n_170),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_176),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_167),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_219),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_199),
.B1(n_210),
.B2(n_211),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_178),
.A2(n_199),
.B1(n_210),
.B2(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_178),
.Y(n_338)
);

AO21x2_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_185),
.B(n_193),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_194),
.B1(n_195),
.B2(n_197),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_184),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_185),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_190),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g273 ( 
.A(n_196),
.Y(n_273)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_204),
.Y(n_334)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_207),
.Y(n_361)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_210),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.C(n_237),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_227),
.A2(n_228),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_230),
.A2(n_237),
.B1(n_238),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_230),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

AOI22x1_ASAP7_75t_L g373 ( 
.A1(n_232),
.A2(n_324),
.B1(n_338),
.B2(n_357),
.Y(n_373)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_235),
.Y(n_315)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_251),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_239),
.B(n_251),
.Y(n_370)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_SL g380 ( 
.A(n_244),
.Y(n_380)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_255),
.Y(n_353)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_382),
.B(n_389),
.Y(n_264)
);

AOI21x1_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_364),
.B(n_381),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_348),
.Y(n_266)
);

AOI21x1_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_302),
.B(n_345),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_290),
.B(n_301),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_282),
.Y(n_269)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_300),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_300),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_292),
.Y(n_344)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_296),
.Y(n_343)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_340),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_322),
.B1(n_323),
.B2(n_339),
.Y(n_303)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_SL g346 ( 
.A(n_304),
.B(n_322),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_312),
.B1(n_316),
.B2(n_321),
.Y(n_304)
);

NAND2xp33_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_322),
.B(n_339),
.Y(n_349)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_339),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_335),
.B2(n_338),
.Y(n_323)
);

NAND2x1_ASAP7_75t_SL g356 ( 
.A(n_324),
.B(n_357),
.Y(n_356)
);

NAND2x1_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_338),
.Y(n_355)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_SL g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_340),
.A2(n_346),
.B(n_347),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_349),
.A2(n_365),
.B(n_366),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_350),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

MAJx2_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_362),
.C(n_368),
.Y(n_367)
);

A2O1A1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B(n_362),
.C(n_363),
.Y(n_354)
);

NAND3xp33_ASAP7_75t_L g363 ( 
.A(n_355),
.B(n_356),
.C(n_362),
.Y(n_363)
);

NAND2xp33_ASAP7_75t_R g368 ( 
.A(n_355),
.B(n_356),
.Y(n_368)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NOR2x1_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_369),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_370),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_373),
.B1(n_374),
.B2(n_375),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_374),
.C(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_387),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_383),
.B(n_387),
.Y(n_389)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);


endmodule