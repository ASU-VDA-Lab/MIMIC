module fake_jpeg_6680_n_165 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_42),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_3),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_3),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_18),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_58),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_24),
.B1(n_27),
.B2(n_20),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_52),
.B1(n_28),
.B2(n_21),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_51),
.B(n_64),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_24),
.B1(n_27),
.B2(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_45),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_63),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_19),
.C(n_26),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_72),
.B(n_14),
.Y(n_80)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_18),
.B(n_27),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_62),
.C(n_6),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_33),
.A2(n_18),
.B1(n_24),
.B2(n_29),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_20),
.B1(n_19),
.B2(n_25),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_66),
.B1(n_67),
.B2(n_29),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_30),
.C(n_26),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_29),
.B(n_14),
.C(n_13),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_33),
.A2(n_25),
.B1(n_28),
.B2(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_71),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_13),
.B(n_14),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_37),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_83),
.Y(n_100)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_59),
.B(n_62),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_37),
.B1(n_10),
.B2(n_11),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_96),
.B1(n_65),
.B2(n_57),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_6),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_96),
.Y(n_109)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_81),
.B1(n_78),
.B2(n_79),
.Y(n_112)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_95),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_65),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_97),
.Y(n_102)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_104),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_110),
.B(n_94),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_87),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_85),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_49),
.A3(n_53),
.B1(n_48),
.B2(n_66),
.C1(n_58),
.C2(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_48),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_101),
.B1(n_107),
.B2(n_86),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_69),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_121),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_126),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_89),
.C(n_83),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_78),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_129),
.B(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_128),
.A2(n_107),
.B1(n_101),
.B2(n_121),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_134),
.B(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_132),
.B(n_138),
.Y(n_144)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_112),
.B1(n_98),
.B2(n_95),
.Y(n_133)
);

AO221x1_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_74),
.B1(n_68),
.B2(n_73),
.C(n_118),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_128),
.A2(n_99),
.B1(n_98),
.B2(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_122),
.B(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_102),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_135),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_SL g142 ( 
.A(n_133),
.B(n_117),
.C(n_105),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_148),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_145),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_125),
.C(n_120),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_92),
.B(n_90),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_133),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_153),
.B(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_152),
.B(n_154),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_141),
.A2(n_136),
.B(n_134),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_149),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_9),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_157),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_147),
.A3(n_143),
.B1(n_145),
.B2(n_130),
.C1(n_91),
.C2(n_102),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_150),
.C(n_68),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_9),
.C(n_73),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_159),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_162),
.Y(n_165)
);


endmodule