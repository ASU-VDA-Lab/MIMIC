module fake_netlist_6_2242_n_2140 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2140);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2140;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_134),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_34),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_152),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_164),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_81),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_100),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_79),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_85),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_47),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_114),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_118),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_105),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_38),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_1),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_179),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_78),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_0),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_5),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_50),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_90),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_38),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_23),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_154),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_65),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_50),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_94),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_166),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_104),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_1),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_170),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_198),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_191),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_80),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_136),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_71),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_65),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_12),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_64),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_147),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_184),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_71),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_4),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_84),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_197),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_145),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_36),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_101),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_128),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_15),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_45),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_95),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_121),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_47),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_68),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_89),
.Y(n_273)
);

INVx4_ASAP7_75t_R g274 ( 
.A(n_57),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_88),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_49),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_160),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_211),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_83),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_87),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_139),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_172),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_23),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_35),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_210),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_115),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_149),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_108),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_148),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_60),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_177),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_82),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_131),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_135),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_167),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_42),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_123),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_6),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_98),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_59),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_39),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_202),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_157),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_17),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_181),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_103),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_21),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_76),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_168),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_150),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_207),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_14),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_195),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_56),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_0),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_75),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_6),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_127),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_158),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_205),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_67),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_36),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_122),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_22),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_35),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_16),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_11),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_162),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_143),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_26),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_59),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_175),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_29),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_33),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_97),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_48),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_138),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_5),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_20),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_37),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_132),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_74),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_190),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_49),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_24),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_111),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_91),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_70),
.Y(n_348)
);

BUFx10_ASAP7_75t_L g349 ( 
.A(n_129),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_199),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_60),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_174),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_28),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_144),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_142),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_62),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_34),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_182),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_193),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_189),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_183),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_42),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_63),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_4),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_64),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_37),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_102),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_10),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_86),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_33),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_169),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_187),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_156),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_77),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_69),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_56),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_141),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_24),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_52),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_43),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_163),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_73),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_107),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_57),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_130),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_153),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_62),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_41),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_67),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_72),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_66),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_44),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_52),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_133),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_16),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_54),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_196),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_176),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_46),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_3),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_72),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_45),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_13),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_119),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_161),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_28),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_55),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_58),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_178),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_3),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_17),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_171),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_70),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_20),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_12),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_200),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_93),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_165),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_206),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_29),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_31),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_15),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_354),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_278),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_214),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_345),
.Y(n_426)
);

INVxp33_ASAP7_75t_SL g427 ( 
.A(n_260),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_218),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_219),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_389),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_220),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_345),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_354),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_345),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_345),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_345),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_224),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_279),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_345),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_280),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_226),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_370),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_370),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_370),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_215),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_370),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_370),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_370),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_228),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_314),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_222),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_314),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_246),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_293),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_305),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_246),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_256),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_232),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_234),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_217),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_221),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_237),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_240),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_245),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_311),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_249),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_352),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_247),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_355),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_246),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_421),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_360),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_252),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_243),
.B(n_2),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_421),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_217),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_230),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_304),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_257),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_258),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_262),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_304),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_304),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_340),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_302),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_229),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_263),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_221),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_340),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_266),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_247),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_340),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_356),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_356),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_269),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_356),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_247),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_273),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_281),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_287),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_294),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_243),
.B(n_2),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_270),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_270),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_365),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_295),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_297),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_365),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_229),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_365),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_299),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_303),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_308),
.Y(n_513)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_270),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_309),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_313),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_319),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_393),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_393),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_393),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_235),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_328),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_329),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_332),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_235),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_264),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_341),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_320),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_264),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_271),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_271),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_426),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_468),
.B(n_320),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_432),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_432),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_434),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_434),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_435),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_491),
.B(n_244),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_435),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_436),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_497),
.B(n_244),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_445),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_503),
.B(n_342),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_430),
.A2(n_476),
.B1(n_433),
.B2(n_423),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_425),
.B(n_231),
.Y(n_547)
);

BUFx8_ASAP7_75t_L g548 ( 
.A(n_504),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_436),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_439),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_439),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_442),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_514),
.B(n_320),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_451),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_442),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_528),
.B(n_310),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_443),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_443),
.B(n_216),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_428),
.B(n_248),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_444),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_444),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_446),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_446),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_447),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_447),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_448),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_478),
.B(n_380),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_448),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_453),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_521),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_457),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_521),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_453),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_456),
.A2(n_310),
.B(n_227),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_456),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_470),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_478),
.B(n_310),
.Y(n_577)
);

NOR2x1_ASAP7_75t_L g578 ( 
.A(n_474),
.B(n_223),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_470),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_461),
.B(n_223),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_471),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_482),
.B(n_225),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_471),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_475),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_475),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_488),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_502),
.B(n_343),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_531),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_477),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_525),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_525),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_526),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_526),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_504),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_529),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_529),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_485),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_530),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_530),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_531),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_482),
.B(n_347),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_483),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_483),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_484),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_484),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_489),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_489),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_492),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_492),
.B(n_350),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_429),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_493),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_493),
.B(n_494),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_494),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_496),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_431),
.B(n_292),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_496),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_505),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_437),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_571),
.B(n_460),
.Y(n_619)
);

INVx6_ASAP7_75t_L g620 ( 
.A(n_548),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_532),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_602),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_556),
.B(n_505),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_532),
.Y(n_624)
);

INVxp67_ASAP7_75t_SL g625 ( 
.A(n_594),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_535),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_535),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_547),
.B(n_441),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_535),
.Y(n_629)
);

INVxp33_ASAP7_75t_L g630 ( 
.A(n_589),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_536),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_571),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_618),
.B(n_380),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_602),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_618),
.B(n_357),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_536),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_587),
.A2(n_495),
.B1(n_513),
.B2(n_490),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_604),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_604),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_559),
.B(n_449),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_603),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_603),
.Y(n_642)
);

BUFx4f_ASAP7_75t_L g643 ( 
.A(n_574),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_615),
.B(n_458),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_604),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_532),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_545),
.B(n_459),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_556),
.B(n_508),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_536),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_605),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_544),
.B(n_462),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_605),
.Y(n_652)
);

NAND3xp33_ASAP7_75t_L g653 ( 
.A(n_578),
.B(n_452),
.C(n_450),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_607),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_545),
.B(n_463),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_607),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_587),
.B(n_464),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_608),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_608),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_594),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_544),
.B(n_466),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_611),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_611),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_557),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_557),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_613),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_613),
.Y(n_667)
);

AND2x2_ASAP7_75t_SL g668 ( 
.A(n_556),
.B(n_251),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_604),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_557),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_578),
.A2(n_427),
.B1(n_324),
.B2(n_339),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_561),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_614),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_532),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_614),
.Y(n_675)
);

INVx4_ASAP7_75t_SL g676 ( 
.A(n_558),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_561),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_594),
.Y(n_678)
);

AND2x6_ASAP7_75t_L g679 ( 
.A(n_533),
.B(n_216),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_554),
.B(n_473),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_617),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_532),
.Y(n_682)
);

CKINVDCx6p67_ASAP7_75t_R g683 ( 
.A(n_597),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_561),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_533),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_617),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_533),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_554),
.B(n_479),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_568),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_604),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_540),
.A2(n_524),
.B1(n_517),
.B2(n_480),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_553),
.A2(n_324),
.B1(n_339),
.B2(n_317),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_568),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_568),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_604),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_553),
.B(n_481),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_548),
.B(n_487),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_604),
.Y(n_698)
);

BUFx8_ASAP7_75t_SL g699 ( 
.A(n_597),
.Y(n_699)
);

INVxp33_ASAP7_75t_SL g700 ( 
.A(n_610),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_532),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_586),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_574),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_574),
.Y(n_704)
);

INVx4_ASAP7_75t_SL g705 ( 
.A(n_558),
.Y(n_705)
);

AND3x2_ASAP7_75t_L g706 ( 
.A(n_553),
.B(n_413),
.C(n_277),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_546),
.A2(n_498),
.B1(n_500),
.B2(n_499),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_569),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_569),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_548),
.B(n_501),
.Y(n_710)
);

AND3x2_ASAP7_75t_L g711 ( 
.A(n_582),
.B(n_277),
.C(n_251),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_601),
.B(n_506),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_574),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_574),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_569),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_548),
.B(n_507),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_586),
.Y(n_717)
);

AND3x2_ASAP7_75t_L g718 ( 
.A(n_582),
.B(n_318),
.C(n_291),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_612),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_612),
.Y(n_720)
);

CKINVDCx11_ASAP7_75t_R g721 ( 
.A(n_546),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_540),
.A2(n_543),
.B1(n_580),
.B2(n_582),
.Y(n_722)
);

CKINVDCx11_ASAP7_75t_R g723 ( 
.A(n_580),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_612),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_586),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_543),
.B(n_511),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_601),
.B(n_512),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_537),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_569),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_609),
.B(n_515),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_609),
.B(n_516),
.Y(n_731)
);

NOR2x1p5_ASAP7_75t_L g732 ( 
.A(n_570),
.B(n_322),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_567),
.B(n_523),
.C(n_522),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_569),
.Y(n_734)
);

INVxp67_ASAP7_75t_SL g735 ( 
.A(n_586),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_SL g736 ( 
.A(n_570),
.B(n_424),
.Y(n_736)
);

INVx5_ASAP7_75t_L g737 ( 
.A(n_558),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_569),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_532),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_537),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_541),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_569),
.Y(n_742)
);

OR2x6_ASAP7_75t_L g743 ( 
.A(n_567),
.B(n_317),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_586),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_541),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_580),
.B(n_527),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_542),
.B(n_508),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_L g748 ( 
.A1(n_572),
.A2(n_238),
.B1(n_241),
.B2(n_233),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_586),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_573),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_573),
.Y(n_751)
);

INVx4_ASAP7_75t_L g752 ( 
.A(n_586),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_573),
.Y(n_753)
);

INVxp33_ASAP7_75t_L g754 ( 
.A(n_577),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_572),
.B(n_486),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_580),
.B(n_509),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_573),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_573),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_573),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_577),
.A2(n_455),
.B1(n_472),
.B2(n_469),
.Y(n_760)
);

BUFx4f_ASAP7_75t_L g761 ( 
.A(n_588),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_592),
.B(n_510),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_573),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_542),
.B(n_510),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_606),
.B(n_520),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_579),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_579),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_577),
.B(n_519),
.C(n_518),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_579),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_606),
.B(n_520),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_549),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_668),
.B(n_588),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_668),
.B(n_588),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_685),
.B(n_216),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_657),
.B(n_588),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_728),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_719),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_660),
.B(n_606),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_647),
.B(n_588),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_L g780 ( 
.A(n_703),
.B(n_216),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_632),
.B(n_254),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_685),
.B(n_588),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_687),
.B(n_588),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_687),
.A2(n_595),
.B(n_596),
.C(n_592),
.Y(n_784)
);

OR2x6_ASAP7_75t_L g785 ( 
.A(n_620),
.B(n_225),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_719),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_728),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_712),
.B(n_590),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_722),
.B(n_590),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_655),
.B(n_590),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_733),
.B(n_616),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_754),
.B(n_590),
.Y(n_792)
);

OAI22xp33_ASAP7_75t_L g793 ( 
.A1(n_696),
.A2(n_227),
.B1(n_261),
.B2(n_250),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_643),
.B(n_216),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_632),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_720),
.A2(n_318),
.B1(n_335),
.B2(n_291),
.Y(n_796)
);

O2A1O1Ixp5_ASAP7_75t_L g797 ( 
.A1(n_643),
.A2(n_616),
.B(n_335),
.C(n_551),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_644),
.B(n_590),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_727),
.B(n_590),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_623),
.B(n_438),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_740),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_720),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_623),
.B(n_590),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_724),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_740),
.Y(n_805)
);

BUFx8_ASAP7_75t_L g806 ( 
.A(n_678),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_699),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_648),
.B(n_591),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_648),
.B(n_591),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_724),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_622),
.B(n_591),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_688),
.B(n_440),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_643),
.B(n_216),
.Y(n_813)
);

OAI221xp5_ASAP7_75t_L g814 ( 
.A1(n_692),
.A2(n_411),
.B1(n_336),
.B2(n_396),
.C(n_348),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_741),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_770),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_741),
.Y(n_817)
);

INVxp67_ASAP7_75t_SL g818 ( 
.A(n_703),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_745),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_622),
.B(n_591),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_704),
.Y(n_821)
);

INVx6_ASAP7_75t_L g822 ( 
.A(n_620),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_745),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_755),
.B(n_454),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_634),
.B(n_591),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_770),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_771),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_704),
.B(n_369),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_660),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_634),
.B(n_591),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_625),
.B(n_616),
.Y(n_831)
);

NAND2x1_ASAP7_75t_L g832 ( 
.A(n_713),
.B(n_558),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_713),
.B(n_714),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_732),
.A2(n_671),
.B1(n_731),
.B2(n_730),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_765),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_714),
.B(n_369),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_771),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_626),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_630),
.B(n_465),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_641),
.B(n_591),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_732),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_641),
.B(n_549),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_642),
.B(n_551),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_707),
.B(n_369),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_736),
.A2(n_467),
.B1(n_359),
.B2(n_361),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_678),
.B(n_518),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_706),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_633),
.Y(n_848)
);

NAND3xp33_ASAP7_75t_L g849 ( 
.A(n_653),
.B(n_239),
.C(n_236),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_626),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_642),
.B(n_552),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_627),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_650),
.B(n_552),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_628),
.B(n_326),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_726),
.A2(n_386),
.B1(n_358),
.B2(n_367),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_627),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_640),
.B(n_382),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_669),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_L g859 ( 
.A(n_679),
.B(n_369),
.Y(n_859)
);

NOR2xp67_ASAP7_75t_L g860 ( 
.A(n_637),
.B(n_595),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_629),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_765),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_743),
.A2(n_412),
.B1(n_323),
.B2(n_374),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_650),
.B(n_555),
.Y(n_864)
);

AND2x6_ASAP7_75t_L g865 ( 
.A(n_690),
.B(n_250),
.Y(n_865)
);

NAND3xp33_ASAP7_75t_SL g866 ( 
.A(n_619),
.B(n_283),
.C(n_259),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_768),
.B(n_596),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_743),
.Y(n_868)
);

INVxp33_ASAP7_75t_L g869 ( 
.A(n_760),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_652),
.B(n_555),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_652),
.B(n_563),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_735),
.A2(n_564),
.B(n_563),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_629),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_654),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_620),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_654),
.B(n_369),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_743),
.Y(n_877)
);

NAND2xp33_ASAP7_75t_L g878 ( 
.A(n_679),
.B(n_369),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_620),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_669),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_656),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_743),
.A2(n_394),
.B1(n_275),
.B2(n_282),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_656),
.B(n_371),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_658),
.B(n_564),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_683),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_635),
.B(n_422),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_658),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_659),
.B(n_372),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_659),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_679),
.A2(n_306),
.B1(n_261),
.B2(n_275),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_662),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_662),
.B(n_565),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_691),
.B(n_242),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_663),
.B(n_666),
.Y(n_894)
);

NAND2x1p5_ASAP7_75t_L g895 ( 
.A(n_737),
.B(n_282),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_663),
.B(n_565),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_666),
.B(n_566),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_667),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_631),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_631),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_667),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_673),
.B(n_566),
.Y(n_902)
);

NOR3xp33_ASAP7_75t_L g903 ( 
.A(n_721),
.B(n_519),
.C(n_255),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_673),
.B(n_575),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_679),
.A2(n_377),
.B1(n_316),
.B2(n_404),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_633),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_635),
.B(n_599),
.Y(n_907)
);

OR2x6_ASAP7_75t_L g908 ( 
.A(n_633),
.B(n_697),
.Y(n_908)
);

AOI221xp5_ASAP7_75t_L g909 ( 
.A1(n_748),
.A2(n_307),
.B1(n_315),
.B2(n_333),
.C(n_391),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_761),
.A2(n_286),
.B(n_285),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_711),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_675),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_651),
.B(n_253),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_L g914 ( 
.A(n_679),
.B(n_558),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_669),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_636),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_675),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_681),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_636),
.Y(n_919)
);

BUFx6f_ASAP7_75t_SL g920 ( 
.A(n_635),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_681),
.B(n_575),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_718),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_635),
.B(n_599),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_762),
.A2(n_362),
.B(n_364),
.C(n_348),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_686),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_633),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_686),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_649),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_737),
.B(n_381),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_649),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_737),
.B(n_385),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_679),
.B(n_575),
.Y(n_932)
);

OAI22xp33_ASAP7_75t_L g933 ( 
.A1(n_747),
.A2(n_285),
.B1(n_286),
.B2(n_288),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_661),
.B(n_267),
.Y(n_934)
);

O2A1O1Ixp5_ASAP7_75t_L g935 ( 
.A1(n_761),
.A2(n_746),
.B(n_690),
.C(n_709),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_737),
.B(n_397),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_621),
.B(n_575),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_756),
.B(n_268),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_764),
.Y(n_939)
);

NOR2xp67_ASAP7_75t_L g940 ( 
.A(n_710),
.B(n_593),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_680),
.A2(n_419),
.B1(n_398),
.B2(n_405),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_737),
.B(n_416),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_702),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_664),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_854),
.A2(n_716),
.B(n_289),
.C(n_306),
.Y(n_945)
);

NOR2xp67_ASAP7_75t_L g946 ( 
.A(n_795),
.B(n_708),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_844),
.A2(n_288),
.B(n_316),
.C(n_289),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_829),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_822),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_776),
.Y(n_950)
);

AOI21xp33_ASAP7_75t_L g951 ( 
.A1(n_857),
.A2(n_700),
.B(n_337),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_772),
.A2(n_700),
.B1(n_761),
.B2(n_337),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_773),
.A2(n_639),
.B(n_638),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_807),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_SL g955 ( 
.A(n_885),
.B(n_683),
.Y(n_955)
);

NOR2x1_ASAP7_75t_L g956 ( 
.A(n_875),
.B(n_366),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_939),
.B(n_621),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_939),
.B(n_621),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_795),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_925),
.B(n_624),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_788),
.A2(n_639),
.B(n_638),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_925),
.B(n_624),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_776),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_818),
.B(n_624),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_872),
.A2(n_639),
.B(n_638),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_869),
.B(n_723),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_869),
.B(n_645),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_794),
.A2(n_769),
.B(n_709),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_800),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_777),
.B(n_646),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_786),
.B(n_646),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_844),
.A2(n_412),
.B(n_323),
.C(n_346),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_787),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_943),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_839),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_781),
.B(n_593),
.Y(n_976)
);

NOR2xp67_ASAP7_75t_L g977 ( 
.A(n_841),
.B(n_845),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_834),
.B(n_645),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_943),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_779),
.A2(n_698),
.B(n_645),
.Y(n_980)
);

AOI21xp33_ASAP7_75t_L g981 ( 
.A1(n_893),
.A2(n_374),
.B(n_346),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_829),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_841),
.B(n_676),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_822),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_787),
.Y(n_985)
);

NOR3xp33_ASAP7_75t_L g986 ( 
.A(n_866),
.B(n_383),
.C(n_377),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_775),
.A2(n_698),
.B(n_749),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_913),
.A2(n_383),
.B(n_394),
.C(n_404),
.Y(n_988)
);

BUFx4f_ASAP7_75t_L g989 ( 
.A(n_908),
.Y(n_989)
);

NAND2x2_ASAP7_75t_L g990 ( 
.A(n_847),
.B(n_922),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_790),
.A2(n_698),
.B(n_749),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_846),
.B(n_229),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_943),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_799),
.A2(n_780),
.B(n_798),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_891),
.B(n_676),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_780),
.A2(n_789),
.B(n_794),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_813),
.A2(n_752),
.B(n_749),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_802),
.B(n_646),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_813),
.A2(n_752),
.B(n_695),
.Y(n_999)
);

BUFx12f_ASAP7_75t_L g1000 ( 
.A(n_806),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_828),
.A2(n_715),
.B(n_708),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_804),
.B(n_674),
.Y(n_1002)
);

AOI21x1_ASAP7_75t_L g1003 ( 
.A1(n_828),
.A2(n_729),
.B(n_715),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_803),
.A2(n_752),
.B(n_695),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_810),
.B(n_674),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_808),
.A2(n_695),
.B(n_669),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_891),
.B(n_676),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_816),
.B(n_674),
.Y(n_1008)
);

O2A1O1Ixp5_ASAP7_75t_L g1009 ( 
.A1(n_797),
.A2(n_689),
.B(n_664),
.C(n_665),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_836),
.A2(n_734),
.B(n_729),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_809),
.A2(n_695),
.B(n_669),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_801),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_836),
.A2(n_409),
.B(n_598),
.C(n_593),
.Y(n_1013)
);

AOI21x1_ASAP7_75t_L g1014 ( 
.A1(n_832),
.A2(n_738),
.B(n_734),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_801),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_833),
.A2(n_769),
.B(n_742),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_SL g1017 ( 
.A(n_885),
.B(n_807),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_833),
.A2(n_742),
.B(n_738),
.Y(n_1018)
);

NOR2x1p5_ASAP7_75t_L g1019 ( 
.A(n_886),
.B(n_272),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_935),
.A2(n_767),
.B(n_751),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_805),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_805),
.Y(n_1022)
);

NAND2x1p5_ASAP7_75t_L g1023 ( 
.A(n_875),
.B(n_702),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_815),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_934),
.A2(n_860),
.B(n_784),
.C(n_867),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_792),
.A2(n_695),
.B(n_702),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_824),
.B(n_229),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_826),
.B(n_682),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_782),
.A2(n_717),
.B(n_702),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_783),
.A2(n_717),
.B(n_702),
.Y(n_1030)
);

NOR3xp33_ASAP7_75t_L g1031 ( 
.A(n_812),
.B(n_409),
.C(n_284),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_774),
.A2(n_751),
.B(n_750),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_910),
.A2(n_725),
.B(n_717),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_874),
.B(n_682),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_907),
.Y(n_1035)
);

BUFx4f_ASAP7_75t_L g1036 ( 
.A(n_908),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_835),
.B(n_276),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_829),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_923),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_868),
.Y(n_1040)
);

BUFx4f_ASAP7_75t_L g1041 ( 
.A(n_908),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_938),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_SL g1043 ( 
.A(n_924),
.B(n_298),
.C(n_290),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_881),
.B(n_682),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_831),
.A2(n_725),
.B(n_717),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_774),
.A2(n_767),
.B(n_753),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_868),
.B(n_676),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_848),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_877),
.B(n_705),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_817),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_831),
.A2(n_725),
.B(n_717),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_877),
.B(n_705),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_887),
.B(n_701),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_889),
.B(n_898),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_901),
.B(n_701),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_831),
.A2(n_744),
.B(n_725),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_912),
.B(n_701),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_817),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_917),
.B(n_739),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_791),
.A2(n_766),
.B1(n_763),
.B2(n_759),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_819),
.Y(n_1061)
);

O2A1O1Ixp5_ASAP7_75t_L g1062 ( 
.A1(n_894),
.A2(n_670),
.B(n_672),
.C(n_677),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_814),
.A2(n_396),
.B1(n_392),
.B2(n_364),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_819),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_862),
.B(n_300),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_823),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_943),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_918),
.B(n_301),
.Y(n_1068)
);

AOI21x1_ASAP7_75t_L g1069 ( 
.A1(n_811),
.A2(n_753),
.B(n_750),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_927),
.B(n_739),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_806),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_821),
.A2(n_766),
.B1(n_763),
.B2(n_759),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_778),
.A2(n_744),
.B(n_725),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_849),
.B(n_312),
.Y(n_1074)
);

AO21x1_ASAP7_75t_L g1075 ( 
.A1(n_883),
.A2(n_758),
.B(n_757),
.Y(n_1075)
);

CKINVDCx6p67_ASAP7_75t_R g1076 ( 
.A(n_920),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_867),
.B(n_296),
.Y(n_1077)
);

BUFx12f_ASAP7_75t_L g1078 ( 
.A(n_847),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_778),
.A2(n_744),
.B(n_757),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_821),
.B(n_867),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_778),
.A2(n_744),
.B(n_758),
.Y(n_1081)
);

INVx4_ASAP7_75t_L g1082 ( 
.A(n_822),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_821),
.A2(n_744),
.B(n_739),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_823),
.B(n_665),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_937),
.A2(n_672),
.B(n_670),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_859),
.A2(n_684),
.B(n_694),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_906),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_827),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_827),
.A2(n_417),
.B1(n_418),
.B2(n_693),
.Y(n_1089)
);

AOI21x1_ASAP7_75t_L g1090 ( 
.A1(n_820),
.A2(n_684),
.B(n_694),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_859),
.A2(n_693),
.B(n_689),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_837),
.B(n_677),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_793),
.A2(n_600),
.B(n_598),
.C(n_362),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_829),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_878),
.A2(n_600),
.B(n_598),
.Y(n_1095)
);

OAI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_909),
.A2(n_387),
.B(n_384),
.Y(n_1096)
);

CKINVDCx6p67_ASAP7_75t_R g1097 ( 
.A(n_920),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_904),
.A2(n_558),
.B(n_600),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_879),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_837),
.B(n_584),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_878),
.A2(n_576),
.B(n_560),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_926),
.B(n_321),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_825),
.A2(n_576),
.B(n_560),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_842),
.B(n_584),
.Y(n_1104)
);

BUFx12f_ASAP7_75t_L g1105 ( 
.A(n_911),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_903),
.B(n_296),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_940),
.B(n_921),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_830),
.A2(n_576),
.B(n_560),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_843),
.B(n_584),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_933),
.A2(n_415),
.B(n_410),
.C(n_392),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_851),
.B(n_584),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_911),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_840),
.A2(n_560),
.B(n_550),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_863),
.A2(n_399),
.B1(n_330),
.B2(n_331),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_883),
.A2(n_410),
.B(n_415),
.C(n_585),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_838),
.Y(n_1116)
);

AOI21xp33_ASAP7_75t_L g1117 ( 
.A1(n_888),
.A2(n_325),
.B(n_327),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_888),
.B(n_334),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_853),
.A2(n_581),
.B(n_585),
.C(n_583),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_838),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_864),
.A2(n_892),
.B(n_870),
.C(n_871),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_796),
.A2(n_401),
.B1(n_344),
.B2(n_351),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_884),
.B(n_584),
.Y(n_1123)
);

NAND2xp33_ASAP7_75t_L g1124 ( 
.A(n_865),
.B(n_932),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_858),
.A2(n_562),
.B(n_538),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_850),
.Y(n_1126)
);

INVx5_ASAP7_75t_L g1127 ( 
.A(n_865),
.Y(n_1127)
);

BUFx4f_ASAP7_75t_L g1128 ( 
.A(n_908),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_896),
.B(n_338),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_882),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_858),
.A2(n_562),
.B(n_538),
.Y(n_1131)
);

AND2x2_ASAP7_75t_SL g1132 ( 
.A(n_890),
.B(n_584),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_897),
.B(n_584),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_929),
.A2(n_931),
.B1(n_942),
.B2(n_936),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_850),
.A2(n_856),
.B(n_852),
.Y(n_1135)
);

NOR2x1_ASAP7_75t_L g1136 ( 
.A(n_879),
.B(n_581),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1035),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1129),
.B(n_902),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_969),
.Y(n_1139)
);

OR2x4_ASAP7_75t_L g1140 ( 
.A(n_966),
.B(n_920),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_973),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_981),
.A2(n_865),
.B1(n_905),
.B2(n_931),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_965),
.A2(n_914),
.B(n_858),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1129),
.B(n_852),
.Y(n_1144)
);

BUFx12f_ASAP7_75t_L g1145 ( 
.A(n_1000),
.Y(n_1145)
);

OAI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_951),
.A2(n_941),
.B(n_855),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1042),
.B(n_1039),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_959),
.B(n_880),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_985),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_978),
.A2(n_944),
.B(n_861),
.C(n_856),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_975),
.B(n_1035),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_994),
.A2(n_914),
.B(n_880),
.Y(n_1152)
);

NOR2x1p5_ASAP7_75t_L g1153 ( 
.A(n_1076),
.B(n_353),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_996),
.A2(n_880),
.B(n_915),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_978),
.A2(n_916),
.B(n_861),
.C(n_930),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_997),
.A2(n_915),
.B(n_936),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_976),
.B(n_873),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_974),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_953),
.A2(n_915),
.B(n_942),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_967),
.B(n_873),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1105),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_950),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1087),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1012),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_963),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1025),
.A2(n_930),
.B(n_899),
.C(n_928),
.Y(n_1166)
);

NOR2xp67_ASAP7_75t_L g1167 ( 
.A(n_966),
.B(n_876),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_992),
.B(n_296),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1118),
.A2(n_928),
.B(n_919),
.C(n_916),
.Y(n_1169)
);

INVx5_ASAP7_75t_L g1170 ( 
.A(n_974),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1080),
.A2(n_785),
.B1(n_919),
.B2(n_900),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_974),
.Y(n_1172)
);

CKINVDCx6p67_ASAP7_75t_R g1173 ( 
.A(n_954),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_1097),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1031),
.A2(n_929),
.B1(n_785),
.B2(n_865),
.Y(n_1175)
);

INVx3_ASAP7_75t_SL g1176 ( 
.A(n_1048),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_967),
.B(n_1054),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1027),
.B(n_296),
.Y(n_1178)
);

NOR2xp67_ASAP7_75t_L g1179 ( 
.A(n_1078),
.B(n_876),
.Y(n_1179)
);

OA21x2_ASAP7_75t_L g1180 ( 
.A1(n_1020),
.A2(n_900),
.B(n_899),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_977),
.B(n_705),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1015),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_SL g1183 ( 
.A(n_989),
.B(n_785),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_987),
.A2(n_785),
.B(n_895),
.Y(n_1184)
);

AO22x1_ASAP7_75t_L g1185 ( 
.A1(n_1031),
.A2(n_865),
.B1(n_400),
.B2(n_402),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1118),
.A2(n_865),
.B1(n_895),
.B2(n_265),
.Y(n_1186)
);

INVx5_ASAP7_75t_L g1187 ( 
.A(n_974),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1021),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_990),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1112),
.B(n_363),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1040),
.B(n_705),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1022),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_949),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1112),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1096),
.B(n_368),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1071),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_961),
.A2(n_980),
.B(n_991),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1121),
.B(n_581),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1064),
.B(n_583),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1074),
.A2(n_265),
.B1(n_349),
.B2(n_373),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1019),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1130),
.A2(n_406),
.B(n_403),
.C(n_375),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1024),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_R g1204 ( 
.A(n_1017),
.B(n_376),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_R g1205 ( 
.A(n_955),
.B(n_378),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1045),
.A2(n_534),
.B(n_538),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1077),
.B(n_1130),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1051),
.A2(n_534),
.B(n_538),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1050),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1058),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1132),
.A2(n_420),
.B1(n_379),
.B2(n_388),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_989),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1068),
.B(n_583),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_990),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1036),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_988),
.A2(n_585),
.B(n_274),
.C(n_265),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1040),
.B(n_390),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_949),
.B(n_92),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1102),
.B(n_395),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1102),
.B(n_407),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_979),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1056),
.A2(n_550),
.B(n_562),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1061),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1074),
.A2(n_408),
.B(n_414),
.C(n_349),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1036),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1066),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1004),
.A2(n_550),
.B(n_562),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1037),
.B(n_265),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_979),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_956),
.Y(n_1230)
);

HAxp5_ASAP7_75t_L g1231 ( 
.A(n_1106),
.B(n_274),
.CON(n_1231),
.SN(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1003),
.A2(n_539),
.B(n_562),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_984),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1088),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1037),
.B(n_1065),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1041),
.B(n_349),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1132),
.A2(n_579),
.B1(n_562),
.B2(n_560),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1068),
.B(n_579),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_979),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_957),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_999),
.A2(n_550),
.B(n_562),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1116),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_945),
.A2(n_349),
.B(n_373),
.C(n_579),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1065),
.B(n_373),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1033),
.A2(n_560),
.B(n_550),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1041),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1124),
.A2(n_560),
.B(n_550),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1052),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1128),
.A2(n_579),
.B1(n_550),
.B2(n_539),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_979),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1073),
.A2(n_539),
.B(n_538),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_946),
.B(n_534),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1128),
.A2(n_373),
.B(n_538),
.C(n_534),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_958),
.Y(n_1254)
);

INVx4_ASAP7_75t_L g1255 ( 
.A(n_984),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1043),
.A2(n_986),
.B1(n_1117),
.B2(n_952),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_993),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_986),
.A2(n_558),
.B1(n_539),
.B2(n_538),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1120),
.B(n_534),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1126),
.B(n_534),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_948),
.B(n_534),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1009),
.A2(n_558),
.B(n_539),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1006),
.A2(n_539),
.B(n_558),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1009),
.A2(n_539),
.B(n_213),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1114),
.B(n_7),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1063),
.A2(n_1127),
.B1(n_1134),
.B2(n_964),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1008),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1011),
.A2(n_208),
.B(n_204),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_947),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_993),
.Y(n_1270)
);

NOR3xp33_ASAP7_75t_L g1271 ( 
.A(n_1043),
.B(n_8),
.C(n_9),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1063),
.B(n_10),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_1082),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1026),
.A2(n_201),
.B(n_192),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_993),
.Y(n_1275)
);

AO32x1_ASAP7_75t_L g1276 ( 
.A1(n_1072),
.A2(n_11),
.A3(n_13),
.B1(n_14),
.B2(n_18),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1082),
.B(n_125),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1104),
.A2(n_188),
.B(n_186),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1127),
.B(n_185),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_947),
.A2(n_18),
.B(n_19),
.C(n_21),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1084),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1127),
.A2(n_19),
.B1(n_22),
.B2(n_25),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_993),
.Y(n_1283)
);

INVx4_ASAP7_75t_L g1284 ( 
.A(n_1067),
.Y(n_1284)
);

NAND2xp33_ASAP7_75t_SL g1285 ( 
.A(n_1099),
.B(n_25),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1115),
.A2(n_26),
.B(n_27),
.C(n_30),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1109),
.A2(n_173),
.B(n_159),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1052),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1092),
.Y(n_1289)
);

AO32x1_ASAP7_75t_L g1290 ( 
.A1(n_1089),
.A2(n_27),
.A3(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_1290)
);

INVx4_ASAP7_75t_L g1291 ( 
.A(n_1067),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1127),
.B(n_155),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1099),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1028),
.A2(n_32),
.B1(n_39),
.B2(n_40),
.Y(n_1294)
);

NOR2x1_ASAP7_75t_SL g1295 ( 
.A(n_1067),
.B(n_151),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1122),
.B(n_970),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1067),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1111),
.A2(n_146),
.B(n_140),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_948),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_982),
.B(n_137),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_982),
.B(n_126),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1235),
.A2(n_1038),
.B1(n_1094),
.B2(n_1023),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1158),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1150),
.A2(n_1075),
.A3(n_1119),
.B(n_1030),
.Y(n_1304)
);

NOR2xp67_ASAP7_75t_L g1305 ( 
.A(n_1207),
.B(n_1038),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1168),
.B(n_1178),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1266),
.A2(n_1029),
.A3(n_1133),
.B(n_1123),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1228),
.B(n_1107),
.Y(n_1308)
);

NOR2xp67_ASAP7_75t_SL g1309 ( 
.A(n_1145),
.B(n_1094),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1191),
.Y(n_1310)
);

BUFx8_ASAP7_75t_L g1311 ( 
.A(n_1163),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1244),
.A2(n_1107),
.B1(n_983),
.B2(n_998),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1137),
.B(n_1151),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1266),
.A2(n_1086),
.A3(n_1091),
.B(n_1081),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1197),
.A2(n_1079),
.B(n_968),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1264),
.A2(n_1062),
.B(n_1069),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1146),
.A2(n_972),
.B(n_1013),
.C(n_1110),
.Y(n_1317)
);

AOI31xp67_ASAP7_75t_L g1318 ( 
.A1(n_1198),
.A2(n_1060),
.A3(n_1100),
.B(n_1002),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1232),
.A2(n_1090),
.B(n_1010),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1154),
.A2(n_1062),
.B(n_1085),
.Y(n_1320)
);

AND2x4_ASAP7_75t_SL g1321 ( 
.A(n_1273),
.B(n_1023),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1138),
.A2(n_1083),
.B(n_962),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1143),
.A2(n_1001),
.B(n_1014),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_SL g1324 ( 
.A1(n_1300),
.A2(n_1047),
.B(n_1049),
.C(n_1007),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1166),
.A2(n_1095),
.A3(n_1103),
.B(n_1108),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1176),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1219),
.B(n_1110),
.Y(n_1327)
);

BUFx10_ASAP7_75t_L g1328 ( 
.A(n_1140),
.Y(n_1328)
);

AOI31xp67_ASAP7_75t_L g1329 ( 
.A1(n_1160),
.A2(n_1005),
.A3(n_971),
.B(n_1053),
.Y(n_1329)
);

NOR2xp67_ASAP7_75t_SL g1330 ( 
.A(n_1161),
.B(n_995),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1173),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1177),
.A2(n_960),
.B(n_1135),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1156),
.A2(n_1016),
.B(n_1018),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1264),
.A2(n_1046),
.B(n_1032),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1141),
.Y(n_1335)
);

AO31x2_ASAP7_75t_L g1336 ( 
.A1(n_1171),
.A2(n_1113),
.A3(n_1101),
.B(n_1034),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1256),
.A2(n_1254),
.B1(n_1240),
.B2(n_1157),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1296),
.A2(n_1059),
.B(n_1044),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1220),
.A2(n_972),
.B(n_1093),
.C(n_1013),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1265),
.A2(n_1271),
.B1(n_1272),
.B2(n_1195),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1293),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1201),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1144),
.A2(n_1055),
.B(n_1057),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1240),
.B(n_1070),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1147),
.B(n_1136),
.Y(n_1345)
);

AO32x2_ASAP7_75t_L g1346 ( 
.A1(n_1282),
.A2(n_1093),
.A3(n_1098),
.B1(n_43),
.B2(n_44),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1139),
.B(n_1131),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1254),
.B(n_1125),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1169),
.A2(n_124),
.B(n_120),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1167),
.A2(n_40),
.B(n_41),
.C(n_46),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1171),
.A2(n_117),
.B(n_116),
.Y(n_1351)
);

OAI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1200),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1159),
.A2(n_113),
.B(n_112),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1184),
.A2(n_110),
.B(n_109),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1281),
.B(n_51),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1174),
.Y(n_1356)
);

AO32x2_ASAP7_75t_L g1357 ( 
.A1(n_1282),
.A2(n_53),
.A3(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1238),
.A2(n_106),
.B(n_99),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1175),
.A2(n_61),
.B(n_63),
.C(n_66),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1213),
.A2(n_96),
.B(n_68),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1224),
.A2(n_61),
.B(n_69),
.C(n_73),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1140),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1194),
.B(n_1230),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1194),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1152),
.A2(n_1155),
.B(n_1183),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1246),
.Y(n_1366)
);

AO31x2_ASAP7_75t_L g1367 ( 
.A1(n_1237),
.A2(n_1243),
.A3(n_1253),
.B(n_1247),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1196),
.Y(n_1368)
);

AOI22x1_ASAP7_75t_L g1369 ( 
.A1(n_1267),
.A2(n_1289),
.B1(n_1278),
.B2(n_1298),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_SL g1370 ( 
.A1(n_1301),
.A2(n_1181),
.B(n_1292),
.C(n_1279),
.Y(n_1370)
);

AO32x2_ASAP7_75t_L g1371 ( 
.A1(n_1211),
.A2(n_1237),
.A3(n_1249),
.B1(n_1290),
.B2(n_1276),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1183),
.A2(n_1142),
.B(n_1252),
.Y(n_1372)
);

AO31x2_ASAP7_75t_L g1373 ( 
.A1(n_1245),
.A2(n_1249),
.A3(n_1280),
.B(n_1269),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1149),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1227),
.A2(n_1187),
.B(n_1170),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1202),
.A2(n_1236),
.B(n_1231),
.C(n_1211),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1164),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1170),
.A2(n_1187),
.B(n_1180),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1158),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1170),
.A2(n_1187),
.B(n_1180),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1190),
.B(n_1217),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1268),
.A2(n_1241),
.B(n_1274),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1199),
.A2(n_1259),
.B(n_1260),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1285),
.A2(n_1294),
.B1(n_1215),
.B2(n_1212),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1248),
.A2(n_1288),
.B1(n_1225),
.B2(n_1186),
.Y(n_1385)
);

NAND2x1p5_ASAP7_75t_L g1386 ( 
.A(n_1193),
.B(n_1233),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1204),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1248),
.B(n_1223),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1210),
.B(n_1234),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1162),
.Y(n_1390)
);

NAND3x1_ASAP7_75t_L g1391 ( 
.A(n_1153),
.B(n_1287),
.C(n_1205),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1179),
.B(n_1277),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1165),
.Y(n_1393)
);

AOI221xp5_ASAP7_75t_SL g1394 ( 
.A1(n_1286),
.A2(n_1216),
.B1(n_1199),
.B2(n_1148),
.C(n_1182),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1188),
.A2(n_1203),
.B(n_1226),
.C(n_1209),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1192),
.B(n_1299),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1218),
.B(n_1277),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1189),
.A2(n_1214),
.B(n_1297),
.C(n_1218),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1275),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1261),
.A2(n_1222),
.B(n_1208),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1193),
.B(n_1255),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1158),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1172),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1185),
.B(n_1191),
.Y(n_1404)
);

AO32x2_ASAP7_75t_L g1405 ( 
.A1(n_1290),
.A2(n_1276),
.A3(n_1291),
.B1(n_1284),
.B2(n_1233),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1206),
.A2(n_1251),
.B(n_1262),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1257),
.B(n_1255),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1257),
.B(n_1295),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1172),
.Y(n_1409)
);

AND2x2_ASAP7_75t_SL g1410 ( 
.A(n_1284),
.B(n_1291),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1172),
.B(n_1221),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1262),
.A2(n_1263),
.B(n_1229),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1221),
.A2(n_1229),
.B(n_1239),
.Y(n_1413)
);

O2A1O1Ixp33_ASAP7_75t_SL g1414 ( 
.A1(n_1258),
.A2(n_1276),
.B(n_1290),
.C(n_1250),
.Y(n_1414)
);

AOI221xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1270),
.A2(n_1283),
.B1(n_981),
.B2(n_1265),
.C(n_1272),
.Y(n_1415)
);

NOR3xp33_ASAP7_75t_L g1416 ( 
.A(n_1270),
.B(n_1244),
.C(n_1228),
.Y(n_1416)
);

AO31x2_ASAP7_75t_L g1417 ( 
.A1(n_1270),
.A2(n_1075),
.A3(n_978),
.B(n_1150),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1283),
.B(n_1235),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1283),
.B(n_1246),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1137),
.Y(n_1420)
);

INVx5_ASAP7_75t_L g1421 ( 
.A(n_1158),
.Y(n_1421)
);

AOI221x1_ASAP7_75t_L g1422 ( 
.A1(n_1228),
.A2(n_1031),
.B1(n_981),
.B2(n_1244),
.C(n_1271),
.Y(n_1422)
);

O2A1O1Ixp33_ASAP7_75t_SL g1423 ( 
.A1(n_1300),
.A2(n_981),
.B(n_1025),
.C(n_844),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1235),
.B(n_632),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1242),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1235),
.B(n_632),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1138),
.A2(n_1177),
.B(n_978),
.Y(n_1427)
);

NAND3xp33_ASAP7_75t_L g1428 ( 
.A(n_1228),
.B(n_1244),
.C(n_1235),
.Y(n_1428)
);

OAI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1228),
.A2(n_632),
.B1(n_619),
.B2(n_869),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1232),
.A2(n_1154),
.B(n_1143),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1235),
.A2(n_1177),
.B1(n_1138),
.B2(n_1228),
.Y(n_1431)
);

AOI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1235),
.A2(n_951),
.B1(n_893),
.B2(n_981),
.C(n_1228),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1235),
.B(n_424),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1235),
.B(n_1177),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1232),
.A2(n_1154),
.B(n_1143),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1137),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1197),
.A2(n_994),
.B(n_996),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1197),
.A2(n_994),
.B(n_996),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1235),
.B(n_1177),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1242),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1191),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1235),
.B(n_424),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1246),
.B(n_1035),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1242),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1197),
.A2(n_994),
.B(n_996),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1264),
.A2(n_1150),
.B(n_1197),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1242),
.Y(n_1447)
);

OR2x2_ASAP7_75t_SL g1448 ( 
.A(n_1207),
.B(n_866),
.Y(n_1448)
);

BUFx4f_ASAP7_75t_L g1449 ( 
.A(n_1173),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1176),
.Y(n_1450)
);

AOI221xp5_ASAP7_75t_L g1451 ( 
.A1(n_1235),
.A2(n_951),
.B1(n_893),
.B2(n_981),
.C(n_1228),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1138),
.A2(n_1177),
.B(n_978),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1235),
.B(n_632),
.Y(n_1453)
);

BUFx10_ASAP7_75t_L g1454 ( 
.A(n_1140),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1228),
.A2(n_951),
.B(n_1244),
.C(n_1235),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1235),
.A2(n_1177),
.B1(n_1138),
.B2(n_1228),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1158),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1138),
.A2(n_1177),
.B(n_978),
.Y(n_1458)
);

AOI221x1_ASAP7_75t_L g1459 ( 
.A1(n_1228),
.A2(n_1031),
.B1(n_981),
.B2(n_1244),
.C(n_1271),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_SL g1460 ( 
.A1(n_1300),
.A2(n_981),
.B(n_1025),
.C(n_844),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1232),
.A2(n_1154),
.B(n_1143),
.Y(n_1461)
);

AO32x2_ASAP7_75t_L g1462 ( 
.A1(n_1266),
.A2(n_1282),
.A3(n_1171),
.B1(n_1211),
.B2(n_834),
.Y(n_1462)
);

AOI221xp5_ASAP7_75t_SL g1463 ( 
.A1(n_1265),
.A2(n_981),
.B1(n_1272),
.B2(n_1146),
.C(n_793),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1207),
.B(n_632),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1228),
.A2(n_1244),
.B(n_1146),
.C(n_1235),
.Y(n_1465)
);

OAI22x1_ASAP7_75t_L g1466 ( 
.A1(n_1228),
.A2(n_1244),
.B1(n_1235),
.B2(n_1200),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1197),
.A2(n_994),
.B(n_996),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_SL g1468 ( 
.A1(n_1300),
.A2(n_981),
.B(n_1025),
.C(n_844),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1197),
.A2(n_994),
.B(n_996),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1432),
.A2(n_1451),
.B1(n_1340),
.B2(n_1428),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1424),
.B(n_1426),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1340),
.A2(n_1381),
.B1(n_1327),
.B2(n_1442),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1434),
.A2(n_1439),
.B1(n_1422),
.B2(n_1459),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_SL g1474 ( 
.A1(n_1455),
.A2(n_1429),
.B(n_1428),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1465),
.A2(n_1308),
.B(n_1431),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1466),
.A2(n_1456),
.B1(n_1352),
.B2(n_1452),
.Y(n_1476)
);

BUFx2_ASAP7_75t_SL g1477 ( 
.A(n_1326),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1351),
.A2(n_1458),
.B1(n_1427),
.B2(n_1349),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_SL g1479 ( 
.A1(n_1433),
.A2(n_1387),
.B1(n_1337),
.B2(n_1453),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1364),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1384),
.A2(n_1464),
.B1(n_1448),
.B2(n_1366),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1417),
.Y(n_1482)
);

BUFx12f_ASAP7_75t_L g1483 ( 
.A(n_1311),
.Y(n_1483)
);

BUFx4f_ASAP7_75t_SL g1484 ( 
.A(n_1311),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1421),
.B(n_1408),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1416),
.A2(n_1306),
.B1(n_1384),
.B2(n_1355),
.Y(n_1486)
);

BUFx12f_ASAP7_75t_L g1487 ( 
.A(n_1356),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1366),
.A2(n_1345),
.B1(n_1363),
.B2(n_1418),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1421),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1342),
.Y(n_1490)
);

CKINVDCx11_ASAP7_75t_R g1491 ( 
.A(n_1331),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1421),
.Y(n_1492)
);

BUFx12f_ASAP7_75t_L g1493 ( 
.A(n_1328),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1313),
.B(n_1344),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1360),
.A2(n_1347),
.B1(n_1397),
.B2(n_1392),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1357),
.A2(n_1346),
.B1(n_1463),
.B2(n_1449),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1449),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1310),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1372),
.A2(n_1335),
.B1(n_1440),
.B2(n_1444),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1326),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1450),
.Y(n_1501)
);

BUFx10_ASAP7_75t_L g1502 ( 
.A(n_1368),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1443),
.Y(n_1503)
);

INVx8_ASAP7_75t_L g1504 ( 
.A(n_1303),
.Y(n_1504)
);

INVx6_ASAP7_75t_L g1505 ( 
.A(n_1419),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1341),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1377),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1425),
.A2(n_1447),
.B1(n_1348),
.B2(n_1450),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1463),
.A2(n_1312),
.B(n_1339),
.Y(n_1509)
);

OAI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1389),
.A2(n_1312),
.B1(n_1420),
.B2(n_1436),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1310),
.Y(n_1511)
);

CKINVDCx11_ASAP7_75t_R g1512 ( 
.A(n_1328),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1454),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1390),
.A2(n_1393),
.B1(n_1305),
.B2(n_1443),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1305),
.A2(n_1362),
.B1(n_1369),
.B2(n_1385),
.Y(n_1515)
);

BUFx2_ASAP7_75t_SL g1516 ( 
.A(n_1419),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1338),
.A2(n_1396),
.B1(n_1446),
.B2(n_1404),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1388),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1399),
.B(n_1411),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_SL g1520 ( 
.A1(n_1357),
.A2(n_1346),
.B1(n_1462),
.B2(n_1446),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1391),
.A2(n_1415),
.B1(n_1330),
.B2(n_1309),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1343),
.A2(n_1365),
.B1(n_1354),
.B2(n_1358),
.Y(n_1522)
);

BUFx12f_ASAP7_75t_L g1523 ( 
.A(n_1454),
.Y(n_1523)
);

BUFx12f_ASAP7_75t_L g1524 ( 
.A(n_1303),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1357),
.A2(n_1346),
.B1(n_1462),
.B2(n_1334),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1334),
.A2(n_1332),
.B1(n_1302),
.B2(n_1462),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1359),
.A2(n_1321),
.B1(n_1322),
.B2(n_1441),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1395),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1407),
.A2(n_1415),
.B1(n_1350),
.B2(n_1412),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1370),
.A2(n_1361),
.B1(n_1468),
.B2(n_1460),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1403),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1423),
.A2(n_1394),
.B1(n_1401),
.B2(n_1410),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1406),
.A2(n_1376),
.B1(n_1382),
.B2(n_1316),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_SL g1534 ( 
.A1(n_1371),
.A2(n_1405),
.B1(n_1316),
.B2(n_1353),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1409),
.Y(n_1535)
);

OAI21xp33_ASAP7_75t_L g1536 ( 
.A1(n_1317),
.A2(n_1398),
.B(n_1386),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1315),
.A2(n_1469),
.B1(n_1438),
.B2(n_1467),
.Y(n_1537)
);

CKINVDCx6p67_ASAP7_75t_R g1538 ( 
.A(n_1402),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1371),
.A2(n_1405),
.B1(n_1333),
.B2(n_1414),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1379),
.B(n_1457),
.Y(n_1540)
);

BUFx2_ASAP7_75t_SL g1541 ( 
.A(n_1379),
.Y(n_1541)
);

CKINVDCx11_ASAP7_75t_R g1542 ( 
.A(n_1379),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1371),
.A2(n_1405),
.B1(n_1445),
.B2(n_1437),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1375),
.A2(n_1380),
.B(n_1378),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1457),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1394),
.B(n_1413),
.Y(n_1546)
);

NAND2x1p5_ASAP7_75t_L g1547 ( 
.A(n_1323),
.B(n_1461),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1417),
.Y(n_1548)
);

BUFx4f_ASAP7_75t_SL g1549 ( 
.A(n_1324),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1400),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1430),
.Y(n_1551)
);

INVxp67_ASAP7_75t_SL g1552 ( 
.A(n_1383),
.Y(n_1552)
);

OAI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1373),
.A2(n_1329),
.B1(n_1367),
.B2(n_1318),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1373),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1307),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1367),
.A2(n_1320),
.B1(n_1435),
.B2(n_1319),
.Y(n_1556)
);

NAND2x1p5_ASAP7_75t_L g1557 ( 
.A(n_1314),
.B(n_1367),
.Y(n_1557)
);

INVxp67_ASAP7_75t_SL g1558 ( 
.A(n_1314),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1307),
.A2(n_1314),
.B1(n_1304),
.B2(n_1336),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1304),
.Y(n_1560)
);

INVx4_ASAP7_75t_L g1561 ( 
.A(n_1304),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1336),
.A2(n_1432),
.B1(n_1451),
.B2(n_1340),
.Y(n_1562)
);

OAI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1325),
.A2(n_1340),
.B1(n_1381),
.B2(n_1432),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1325),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1325),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1437),
.A2(n_1445),
.B(n_1438),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1424),
.B(n_1426),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_1331),
.Y(n_1568)
);

INVx2_ASAP7_75t_R g1569 ( 
.A(n_1421),
.Y(n_1569)
);

INVxp67_ASAP7_75t_SL g1570 ( 
.A(n_1427),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1432),
.A2(n_1451),
.B1(n_1340),
.B2(n_1428),
.Y(n_1571)
);

BUFx12f_ASAP7_75t_L g1572 ( 
.A(n_1311),
.Y(n_1572)
);

INVx6_ASAP7_75t_L g1573 ( 
.A(n_1311),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1313),
.Y(n_1574)
);

BUFx8_ASAP7_75t_L g1575 ( 
.A(n_1341),
.Y(n_1575)
);

INVxp67_ASAP7_75t_SL g1576 ( 
.A(n_1427),
.Y(n_1576)
);

INVx2_ASAP7_75t_SL g1577 ( 
.A(n_1311),
.Y(n_1577)
);

BUFx8_ASAP7_75t_SL g1578 ( 
.A(n_1449),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1327),
.A2(n_1235),
.B1(n_1244),
.B2(n_1228),
.Y(n_1579)
);

BUFx10_ASAP7_75t_L g1580 ( 
.A(n_1356),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1432),
.A2(n_1451),
.B1(n_1244),
.B2(n_1228),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1311),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1310),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1374),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1434),
.B(n_1439),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1374),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1311),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1455),
.A2(n_1465),
.B(n_1451),
.Y(n_1588)
);

INVx4_ASAP7_75t_L g1589 ( 
.A(n_1421),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1434),
.B(n_1439),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1432),
.A2(n_1451),
.B1(n_1340),
.B2(n_1428),
.Y(n_1591)
);

CKINVDCx11_ASAP7_75t_R g1592 ( 
.A(n_1331),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1374),
.Y(n_1593)
);

CKINVDCx11_ASAP7_75t_R g1594 ( 
.A(n_1331),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1327),
.A2(n_1235),
.B1(n_1244),
.B2(n_1228),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1432),
.A2(n_1451),
.B1(n_1327),
.B2(n_1235),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1432),
.A2(n_1451),
.B1(n_1340),
.B2(n_1428),
.Y(n_1597)
);

OAI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1340),
.A2(n_1381),
.B1(n_1451),
.B2(n_1432),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1432),
.A2(n_1451),
.B1(n_1327),
.B2(n_1235),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1432),
.A2(n_1451),
.B1(n_1327),
.B2(n_1235),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1432),
.A2(n_1451),
.B1(n_1327),
.B2(n_1235),
.Y(n_1601)
);

INVx8_ASAP7_75t_L g1602 ( 
.A(n_1421),
.Y(n_1602)
);

BUFx10_ASAP7_75t_L g1603 ( 
.A(n_1356),
.Y(n_1603)
);

BUFx4f_ASAP7_75t_SL g1604 ( 
.A(n_1311),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_SL g1605 ( 
.A1(n_1327),
.A2(n_1235),
.B1(n_1244),
.B2(n_1228),
.Y(n_1605)
);

CKINVDCx11_ASAP7_75t_R g1606 ( 
.A(n_1331),
.Y(n_1606)
);

INVx8_ASAP7_75t_L g1607 ( 
.A(n_1421),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1311),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1311),
.Y(n_1609)
);

BUFx12f_ASAP7_75t_L g1610 ( 
.A(n_1311),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1374),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1313),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1432),
.A2(n_1451),
.B1(n_1327),
.B2(n_1235),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1432),
.A2(n_1451),
.B1(n_1340),
.B2(n_1428),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_SL g1615 ( 
.A(n_1311),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1421),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1311),
.Y(n_1617)
);

NAND2x1p5_ASAP7_75t_L g1618 ( 
.A(n_1421),
.B(n_1170),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1313),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_SL g1620 ( 
.A1(n_1327),
.A2(n_1235),
.B1(n_1244),
.B2(n_1228),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1554),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1560),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_L g1623 ( 
.A(n_1581),
.B(n_1571),
.C(n_1470),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1482),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1570),
.B(n_1576),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1564),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1565),
.B(n_1562),
.Y(n_1627)
);

BUFx12f_ASAP7_75t_L g1628 ( 
.A(n_1491),
.Y(n_1628)
);

OAI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1579),
.A2(n_1620),
.B1(n_1595),
.B2(n_1605),
.C(n_1596),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1482),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1548),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1585),
.B(n_1590),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1566),
.A2(n_1547),
.B(n_1537),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1509),
.B(n_1520),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1558),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1557),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1547),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1558),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1557),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1537),
.A2(n_1533),
.B(n_1555),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1555),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1561),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1552),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1552),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1550),
.B(n_1507),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1551),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1546),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1499),
.B(n_1498),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1559),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1602),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1533),
.A2(n_1588),
.B(n_1526),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1528),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1480),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1549),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1494),
.B(n_1598),
.Y(n_1655)
);

INVx3_ASAP7_75t_L g1656 ( 
.A(n_1549),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1520),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1525),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1525),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1496),
.B(n_1475),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1553),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1553),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1539),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1591),
.A2(n_1597),
.B1(n_1614),
.B2(n_1481),
.Y(n_1664)
);

BUFx2_ASAP7_75t_SL g1665 ( 
.A(n_1489),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1598),
.A2(n_1599),
.B1(n_1596),
.B2(n_1600),
.C(n_1601),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1480),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1593),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1539),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_SL g1670 ( 
.A1(n_1477),
.A2(n_1620),
.B1(n_1579),
.B2(n_1595),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1522),
.A2(n_1544),
.B(n_1526),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_R g1672 ( 
.A(n_1483),
.B(n_1572),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1543),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1543),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1611),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1488),
.Y(n_1676)
);

OAI21x1_ASAP7_75t_L g1677 ( 
.A1(n_1522),
.A2(n_1530),
.B(n_1499),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1485),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1472),
.B(n_1471),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_1489),
.Y(n_1680)
);

OAI21xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1476),
.A2(n_1532),
.B(n_1599),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1600),
.B(n_1601),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1510),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1534),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1534),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1574),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1515),
.A2(n_1527),
.B(n_1517),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1556),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1515),
.A2(n_1527),
.B(n_1517),
.Y(n_1689)
);

BUFx12f_ASAP7_75t_L g1690 ( 
.A(n_1592),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1556),
.Y(n_1691)
);

OA21x2_ASAP7_75t_L g1692 ( 
.A1(n_1474),
.A2(n_1476),
.B(n_1536),
.Y(n_1692)
);

BUFx3_ASAP7_75t_L g1693 ( 
.A(n_1575),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1584),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1586),
.Y(n_1695)
);

NOR2x1_ASAP7_75t_SL g1696 ( 
.A(n_1489),
.B(n_1492),
.Y(n_1696)
);

INVxp33_ASAP7_75t_L g1697 ( 
.A(n_1567),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1495),
.A2(n_1514),
.B(n_1521),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1605),
.A2(n_1613),
.B1(n_1478),
.B2(n_1479),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1518),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1612),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1508),
.Y(n_1702)
);

OAI21x1_ASAP7_75t_L g1703 ( 
.A1(n_1495),
.A2(n_1514),
.B(n_1531),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1508),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_L g1705 ( 
.A1(n_1535),
.A2(n_1511),
.B(n_1583),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1563),
.B(n_1619),
.Y(n_1706)
);

INVx2_ASAP7_75t_SL g1707 ( 
.A(n_1602),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1563),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1510),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1529),
.Y(n_1710)
);

OR2x6_ASAP7_75t_L g1711 ( 
.A(n_1602),
.B(n_1607),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1529),
.Y(n_1712)
);

INVx4_ASAP7_75t_L g1713 ( 
.A(n_1607),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1607),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1545),
.Y(n_1715)
);

OR2x6_ASAP7_75t_L g1716 ( 
.A(n_1516),
.B(n_1513),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1473),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1540),
.B(n_1503),
.Y(n_1718)
);

NAND2x1p5_ASAP7_75t_L g1719 ( 
.A(n_1589),
.B(n_1616),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1473),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1519),
.B(n_1616),
.Y(n_1721)
);

BUFx2_ASAP7_75t_L g1722 ( 
.A(n_1505),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1478),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1613),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1505),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1505),
.Y(n_1726)
);

INVx5_ASAP7_75t_L g1727 ( 
.A(n_1492),
.Y(n_1727)
);

OAI21x1_ASAP7_75t_L g1728 ( 
.A1(n_1618),
.A2(n_1486),
.B(n_1569),
.Y(n_1728)
);

OAI21x1_ASAP7_75t_L g1729 ( 
.A1(n_1618),
.A2(n_1486),
.B(n_1541),
.Y(n_1729)
);

OR2x6_ASAP7_75t_L g1730 ( 
.A(n_1493),
.B(n_1523),
.Y(n_1730)
);

OAI21x1_ASAP7_75t_L g1731 ( 
.A1(n_1479),
.A2(n_1504),
.B(n_1524),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1500),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1501),
.B(n_1506),
.Y(n_1733)
);

OAI21x1_ASAP7_75t_L g1734 ( 
.A1(n_1504),
.A2(n_1542),
.B(n_1512),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1502),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1502),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1538),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1575),
.Y(n_1738)
);

AND2x2_ASAP7_75t_SL g1739 ( 
.A(n_1660),
.B(n_1608),
.Y(n_1739)
);

AOI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1623),
.A2(n_1664),
.B1(n_1666),
.B2(n_1681),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1718),
.B(n_1603),
.Y(n_1741)
);

OAI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1681),
.A2(n_1577),
.B(n_1609),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1625),
.B(n_1603),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1715),
.Y(n_1744)
);

O2A1O1Ixp33_ASAP7_75t_SL g1745 ( 
.A1(n_1654),
.A2(n_1568),
.B(n_1615),
.C(n_1484),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1632),
.B(n_1490),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1718),
.B(n_1580),
.Y(n_1747)
);

OR2x6_ASAP7_75t_L g1748 ( 
.A(n_1671),
.B(n_1573),
.Y(n_1748)
);

OR2x2_ASAP7_75t_SL g1749 ( 
.A(n_1692),
.B(n_1573),
.Y(n_1749)
);

OA21x2_ASAP7_75t_L g1750 ( 
.A1(n_1671),
.A2(n_1497),
.B(n_1573),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1715),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1718),
.B(n_1587),
.Y(n_1752)
);

CKINVDCx16_ASAP7_75t_R g1753 ( 
.A(n_1628),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_SL g1754 ( 
.A1(n_1670),
.A2(n_1604),
.B1(n_1610),
.B2(n_1582),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1655),
.B(n_1487),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1721),
.B(n_1617),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_SL g1757 ( 
.A1(n_1629),
.A2(n_1578),
.B1(n_1606),
.B2(n_1594),
.Y(n_1757)
);

AOI221xp5_ASAP7_75t_L g1758 ( 
.A1(n_1699),
.A2(n_1723),
.B1(n_1660),
.B2(n_1720),
.C(n_1717),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1721),
.B(n_1697),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1627),
.B(n_1706),
.Y(n_1760)
);

BUFx3_ASAP7_75t_L g1761 ( 
.A(n_1693),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_SL g1762 ( 
.A(n_1693),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1645),
.Y(n_1763)
);

AO32x2_ASAP7_75t_L g1764 ( 
.A1(n_1663),
.A2(n_1669),
.A3(n_1685),
.B1(n_1684),
.B2(n_1659),
.Y(n_1764)
);

BUFx3_ASAP7_75t_L g1765 ( 
.A(n_1693),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1682),
.A2(n_1724),
.B1(n_1692),
.B2(n_1679),
.Y(n_1766)
);

AND2x6_ASAP7_75t_L g1767 ( 
.A(n_1648),
.B(n_1710),
.Y(n_1767)
);

AND2x4_ASAP7_75t_SL g1768 ( 
.A(n_1732),
.B(n_1686),
.Y(n_1768)
);

CKINVDCx8_ASAP7_75t_R g1769 ( 
.A(n_1665),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1622),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1628),
.Y(n_1771)
);

AOI221xp5_ASAP7_75t_L g1772 ( 
.A1(n_1723),
.A2(n_1724),
.B1(n_1720),
.B2(n_1717),
.C(n_1683),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1716),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_R g1774 ( 
.A(n_1690),
.B(n_1713),
.Y(n_1774)
);

A2O1A1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1687),
.A2(n_1689),
.B(n_1698),
.C(n_1677),
.Y(n_1775)
);

INVx5_ASAP7_75t_L g1776 ( 
.A(n_1711),
.Y(n_1776)
);

AO32x2_ASAP7_75t_L g1777 ( 
.A1(n_1669),
.A2(n_1685),
.A3(n_1684),
.B1(n_1659),
.B2(n_1658),
.Y(n_1777)
);

OAI211xp5_ASAP7_75t_L g1778 ( 
.A1(n_1692),
.A2(n_1683),
.B(n_1676),
.C(n_1709),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1692),
.A2(n_1738),
.B1(n_1690),
.B2(n_1651),
.Y(n_1779)
);

NOR2x1_ASAP7_75t_SL g1780 ( 
.A(n_1716),
.B(n_1647),
.Y(n_1780)
);

AOI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1710),
.A2(n_1712),
.B1(n_1708),
.B2(n_1634),
.C(n_1704),
.Y(n_1781)
);

AO21x2_ASAP7_75t_L g1782 ( 
.A1(n_1633),
.A2(n_1661),
.B(n_1662),
.Y(n_1782)
);

OAI21xp33_ASAP7_75t_SL g1783 ( 
.A1(n_1634),
.A2(n_1689),
.B(n_1687),
.Y(n_1783)
);

AOI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1712),
.A2(n_1708),
.B1(n_1704),
.B2(n_1702),
.C(n_1653),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1737),
.Y(n_1785)
);

OA21x2_ASAP7_75t_L g1786 ( 
.A1(n_1640),
.A2(n_1677),
.B(n_1633),
.Y(n_1786)
);

OR2x6_ASAP7_75t_L g1787 ( 
.A(n_1728),
.B(n_1729),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1737),
.Y(n_1788)
);

AO21x2_ASAP7_75t_L g1789 ( 
.A1(n_1661),
.A2(n_1662),
.B(n_1640),
.Y(n_1789)
);

BUFx4f_ASAP7_75t_SL g1790 ( 
.A(n_1654),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1702),
.A2(n_1657),
.B1(n_1658),
.B2(n_1674),
.C(n_1673),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1698),
.A2(n_1703),
.B(n_1729),
.Y(n_1792)
);

AOI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1657),
.A2(n_1673),
.B1(n_1674),
.B2(n_1649),
.C(n_1667),
.Y(n_1793)
);

OA21x2_ASAP7_75t_L g1794 ( 
.A1(n_1703),
.A2(n_1728),
.B(n_1691),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1647),
.B(n_1701),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1733),
.B(n_1654),
.Y(n_1796)
);

AO21x2_ASAP7_75t_L g1797 ( 
.A1(n_1635),
.A2(n_1638),
.B(n_1644),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1731),
.A2(n_1651),
.B(n_1648),
.Y(n_1798)
);

AO32x2_ASAP7_75t_L g1799 ( 
.A1(n_1650),
.A2(n_1707),
.A3(n_1714),
.B1(n_1713),
.B2(n_1651),
.Y(n_1799)
);

A2O1A1Ixp33_ASAP7_75t_L g1800 ( 
.A1(n_1654),
.A2(n_1656),
.B(n_1649),
.C(n_1734),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1647),
.B(n_1643),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1656),
.B(n_1738),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1734),
.Y(n_1803)
);

INVx3_ASAP7_75t_SL g1804 ( 
.A(n_1730),
.Y(n_1804)
);

OAI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1648),
.A2(n_1705),
.B(n_1652),
.Y(n_1805)
);

OA21x2_ASAP7_75t_L g1806 ( 
.A1(n_1688),
.A2(n_1691),
.B(n_1705),
.Y(n_1806)
);

O2A1O1Ixp33_ASAP7_75t_SL g1807 ( 
.A1(n_1656),
.A2(n_1736),
.B(n_1650),
.C(n_1707),
.Y(n_1807)
);

AO32x2_ASAP7_75t_L g1808 ( 
.A1(n_1714),
.A2(n_1713),
.A3(n_1621),
.B1(n_1688),
.B2(n_1624),
.Y(n_1808)
);

CKINVDCx10_ASAP7_75t_R g1809 ( 
.A(n_1730),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1770),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1797),
.Y(n_1811)
);

NOR2x1p5_ASAP7_75t_L g1812 ( 
.A(n_1803),
.B(n_1678),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1798),
.B(n_1636),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1744),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1751),
.Y(n_1815)
);

INVxp67_ASAP7_75t_L g1816 ( 
.A(n_1806),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1773),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_SL g1818 ( 
.A1(n_1778),
.A2(n_1696),
.B1(n_1631),
.B2(n_1700),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1806),
.B(n_1636),
.Y(n_1819)
);

INVxp67_ASAP7_75t_L g1820 ( 
.A(n_1795),
.Y(n_1820)
);

INVxp67_ASAP7_75t_L g1821 ( 
.A(n_1763),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1759),
.B(n_1639),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1787),
.B(n_1637),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1754),
.A2(n_1722),
.B1(n_1725),
.B2(n_1726),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1801),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1808),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_1768),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1777),
.B(n_1642),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1808),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1799),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1799),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1777),
.B(n_1642),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1789),
.B(n_1626),
.Y(n_1833)
);

AND2x2_ASAP7_75t_SL g1834 ( 
.A(n_1739),
.B(n_1631),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1766),
.B(n_1624),
.Y(n_1835)
);

BUFx2_ASAP7_75t_L g1836 ( 
.A(n_1799),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1766),
.B(n_1630),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1760),
.B(n_1630),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1777),
.B(n_1641),
.Y(n_1839)
);

INVx1_ASAP7_75t_SL g1840 ( 
.A(n_1743),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1764),
.Y(n_1841)
);

BUFx2_ASAP7_75t_L g1842 ( 
.A(n_1749),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1764),
.B(n_1641),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1787),
.B(n_1637),
.Y(n_1844)
);

OAI222xp33_ASAP7_75t_L g1845 ( 
.A1(n_1740),
.A2(n_1716),
.B1(n_1711),
.B2(n_1675),
.C1(n_1695),
.C2(n_1694),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1791),
.B(n_1781),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1746),
.B(n_1755),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1742),
.B(n_1735),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1764),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1805),
.B(n_1646),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1840),
.B(n_1743),
.Y(n_1851)
);

BUFx3_ASAP7_75t_L g1852 ( 
.A(n_1817),
.Y(n_1852)
);

AND2x2_ASAP7_75t_SL g1853 ( 
.A(n_1834),
.B(n_1750),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1820),
.B(n_1794),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1846),
.A2(n_1740),
.B1(n_1754),
.B2(n_1757),
.Y(n_1855)
);

OR2x6_ASAP7_75t_L g1856 ( 
.A(n_1812),
.B(n_1748),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1821),
.Y(n_1857)
);

INVx3_ASAP7_75t_L g1858 ( 
.A(n_1823),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1810),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1820),
.B(n_1782),
.Y(n_1860)
);

BUFx2_ASAP7_75t_L g1861 ( 
.A(n_1842),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1821),
.Y(n_1862)
);

INVx5_ASAP7_75t_L g1863 ( 
.A(n_1830),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1842),
.B(n_1787),
.Y(n_1864)
);

AO21x2_ASAP7_75t_L g1865 ( 
.A1(n_1811),
.A2(n_1792),
.B(n_1775),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1835),
.B(n_1782),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1835),
.B(n_1792),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1839),
.Y(n_1868)
);

NOR2x1p5_ASAP7_75t_L g1869 ( 
.A(n_1846),
.B(n_1761),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1839),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1822),
.B(n_1805),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1823),
.B(n_1780),
.Y(n_1872)
);

INVxp67_ASAP7_75t_L g1873 ( 
.A(n_1825),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1833),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1814),
.Y(n_1875)
);

NAND3xp33_ASAP7_75t_L g1876 ( 
.A(n_1818),
.B(n_1742),
.C(n_1793),
.Y(n_1876)
);

CKINVDCx20_ASAP7_75t_R g1877 ( 
.A(n_1827),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1843),
.Y(n_1878)
);

OAI33xp33_ASAP7_75t_L g1879 ( 
.A1(n_1841),
.A2(n_1779),
.A3(n_1694),
.B1(n_1695),
.B2(n_1735),
.B3(n_1668),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_L g1880 ( 
.A(n_1847),
.B(n_1753),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1843),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1828),
.Y(n_1882)
);

INVxp67_ASAP7_75t_L g1883 ( 
.A(n_1838),
.Y(n_1883)
);

AOI33xp33_ASAP7_75t_L g1884 ( 
.A1(n_1818),
.A2(n_1793),
.A3(n_1758),
.B1(n_1791),
.B2(n_1781),
.B3(n_1772),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1815),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1819),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1837),
.B(n_1786),
.Y(n_1887)
);

AND2x4_ASAP7_75t_L g1888 ( 
.A(n_1823),
.B(n_1776),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1883),
.B(n_1841),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1875),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1875),
.Y(n_1891)
);

NOR2x1_ASAP7_75t_SL g1892 ( 
.A(n_1856),
.B(n_1848),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1887),
.B(n_1830),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1863),
.B(n_1831),
.Y(n_1894)
);

INVx4_ASAP7_75t_L g1895 ( 
.A(n_1856),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1859),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1860),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1863),
.B(n_1831),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1873),
.B(n_1849),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1886),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1886),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1863),
.B(n_1836),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1863),
.B(n_1836),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1876),
.B(n_1834),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1867),
.B(n_1849),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1863),
.B(n_1813),
.Y(n_1906)
);

OAI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1876),
.A2(n_1827),
.B1(n_1804),
.B2(n_1837),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1867),
.B(n_1828),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1886),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1863),
.B(n_1882),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1868),
.B(n_1870),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1878),
.B(n_1813),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1859),
.B(n_1832),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1874),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1860),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1887),
.B(n_1826),
.Y(n_1916)
);

INVx3_ASAP7_75t_L g1917 ( 
.A(n_1872),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1881),
.B(n_1850),
.Y(n_1918)
);

NAND3xp33_ASAP7_75t_L g1919 ( 
.A(n_1855),
.B(n_1772),
.C(n_1784),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1861),
.B(n_1850),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1861),
.B(n_1832),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1858),
.B(n_1823),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1858),
.B(n_1826),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1885),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1858),
.B(n_1829),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1874),
.Y(n_1926)
);

INVx1_ASAP7_75t_SL g1927 ( 
.A(n_1852),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1874),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1858),
.B(n_1844),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1905),
.B(n_1908),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1896),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1896),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1921),
.B(n_1864),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1921),
.B(n_1917),
.Y(n_1934)
);

INVxp33_ASAP7_75t_L g1935 ( 
.A(n_1904),
.Y(n_1935)
);

OAI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1919),
.A2(n_1869),
.B1(n_1800),
.B2(n_1834),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1904),
.B(n_1853),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1924),
.Y(n_1938)
);

INVxp67_ASAP7_75t_L g1939 ( 
.A(n_1905),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1924),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1907),
.B(n_1869),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1890),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1921),
.B(n_1864),
.Y(n_1943)
);

OAI22xp33_ASAP7_75t_SL g1944 ( 
.A1(n_1893),
.A2(n_1866),
.B1(n_1880),
.B2(n_1854),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1908),
.B(n_1866),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1900),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1900),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1927),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1900),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1917),
.B(n_1920),
.Y(n_1950)
);

NAND2x2_ASAP7_75t_L g1951 ( 
.A(n_1919),
.B(n_1765),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1917),
.B(n_1856),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1917),
.B(n_1920),
.Y(n_1953)
);

INVx2_ASAP7_75t_SL g1954 ( 
.A(n_1917),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1920),
.B(n_1856),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1900),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1907),
.B(n_1771),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1890),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1890),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1891),
.Y(n_1960)
);

NAND2x1p5_ASAP7_75t_L g1961 ( 
.A(n_1895),
.B(n_1853),
.Y(n_1961)
);

NOR3xp33_ASAP7_75t_L g1962 ( 
.A(n_1895),
.B(n_1779),
.C(n_1884),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1927),
.B(n_1871),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1891),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1889),
.B(n_1854),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1901),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1895),
.B(n_1856),
.Y(n_1967)
);

NAND2x1p5_ASAP7_75t_L g1968 ( 
.A(n_1895),
.B(n_1853),
.Y(n_1968)
);

INVxp67_ASAP7_75t_L g1969 ( 
.A(n_1899),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1901),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1889),
.B(n_1871),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1893),
.B(n_1899),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1895),
.B(n_1872),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1892),
.B(n_1906),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1891),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1892),
.B(n_1872),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1962),
.B(n_1918),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1935),
.B(n_1918),
.Y(n_1978)
);

NAND2x2_ASAP7_75t_L g1979 ( 
.A(n_1941),
.B(n_1785),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1976),
.B(n_1892),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1976),
.B(n_1894),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1957),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1931),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1931),
.Y(n_1984)
);

NOR3x1_ASAP7_75t_L g1985 ( 
.A(n_1937),
.B(n_1893),
.C(n_1916),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1974),
.B(n_1894),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1948),
.B(n_1918),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1932),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1932),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1955),
.B(n_1894),
.Y(n_1990)
);

BUFx3_ASAP7_75t_L g1991 ( 
.A(n_1948),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1942),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1939),
.B(n_1912),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1936),
.B(n_1912),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1969),
.B(n_1912),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1942),
.Y(n_1996)
);

AOI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1951),
.A2(n_1865),
.B1(n_1888),
.B2(n_1767),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1958),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1958),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1959),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1930),
.B(n_1916),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1959),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1974),
.B(n_1898),
.Y(n_2003)
);

INVx1_ASAP7_75t_SL g2004 ( 
.A(n_1973),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1960),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1944),
.B(n_1963),
.Y(n_2006)
);

NAND4xp25_ASAP7_75t_SL g2007 ( 
.A(n_1967),
.B(n_1898),
.C(n_1902),
.D(n_1903),
.Y(n_2007)
);

NAND2x1_ASAP7_75t_L g2008 ( 
.A(n_1955),
.B(n_1910),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1930),
.B(n_1916),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1944),
.B(n_1857),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1961),
.B(n_1898),
.Y(n_2011)
);

INVxp67_ASAP7_75t_SL g2012 ( 
.A(n_1961),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1951),
.A2(n_1865),
.B1(n_1888),
.B2(n_1767),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1961),
.B(n_1902),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1933),
.B(n_1862),
.Y(n_2015)
);

OAI222xp33_ASAP7_75t_L g2016 ( 
.A1(n_2006),
.A2(n_1968),
.B1(n_1967),
.B2(n_1973),
.C1(n_1972),
.C2(n_1903),
.Y(n_2016)
);

AOI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1982),
.A2(n_1951),
.B1(n_1968),
.B2(n_1952),
.Y(n_2017)
);

AOI21x1_ASAP7_75t_L g2018 ( 
.A1(n_2008),
.A2(n_1940),
.B(n_1938),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1998),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1991),
.B(n_1933),
.Y(n_2020)
);

OAI221xp5_ASAP7_75t_L g2021 ( 
.A1(n_1979),
.A2(n_2010),
.B1(n_1977),
.B2(n_1994),
.C(n_1968),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_SL g2022 ( 
.A(n_1991),
.B(n_1774),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1998),
.Y(n_2023)
);

AOI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_1979),
.A2(n_1865),
.B1(n_1879),
.B2(n_1903),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_2004),
.B(n_1943),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1990),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1990),
.B(n_1943),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_L g2028 ( 
.A(n_2007),
.B(n_1672),
.Y(n_2028)
);

OAI33xp33_ASAP7_75t_L g2029 ( 
.A1(n_1984),
.A2(n_1940),
.A3(n_1938),
.B1(n_1972),
.B2(n_1965),
.B3(n_1975),
.Y(n_2029)
);

OR2x2_ASAP7_75t_L g2030 ( 
.A(n_1978),
.B(n_1971),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1984),
.Y(n_2031)
);

OAI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_2012),
.A2(n_1902),
.B(n_1952),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1988),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1988),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1989),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1990),
.B(n_1950),
.Y(n_2036)
);

OAI221xp5_ASAP7_75t_L g2037 ( 
.A1(n_1997),
.A2(n_1945),
.B1(n_1965),
.B2(n_1954),
.C(n_1950),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1986),
.B(n_1953),
.Y(n_2038)
);

INVx2_ASAP7_75t_SL g2039 ( 
.A(n_2008),
.Y(n_2039)
);

O2A1O1Ixp33_ASAP7_75t_L g2040 ( 
.A1(n_1987),
.A2(n_1745),
.B(n_1954),
.C(n_1945),
.Y(n_2040)
);

AOI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_2013),
.A2(n_1672),
.B(n_1730),
.Y(n_2041)
);

OR2x2_ASAP7_75t_L g2042 ( 
.A(n_2015),
.B(n_1953),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_SL g2043 ( 
.A1(n_2011),
.A2(n_1910),
.B1(n_1906),
.B2(n_1877),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_L g2044 ( 
.A(n_1995),
.B(n_1809),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2019),
.Y(n_2045)
);

AOI221x1_ASAP7_75t_SL g2046 ( 
.A1(n_2020),
.A2(n_1983),
.B1(n_1993),
.B2(n_1989),
.C(n_2005),
.Y(n_2046)
);

NOR3xp33_ASAP7_75t_L g2047 ( 
.A(n_2021),
.B(n_2014),
.C(n_2011),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_2039),
.Y(n_2048)
);

OAI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_2043),
.A2(n_1980),
.B1(n_2003),
.B2(n_1986),
.Y(n_2049)
);

INVx1_ASAP7_75t_SL g2050 ( 
.A(n_2036),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2023),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2031),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_2043),
.B(n_2014),
.Y(n_2053)
);

INVxp67_ASAP7_75t_SL g2054 ( 
.A(n_2018),
.Y(n_2054)
);

AOI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_2022),
.A2(n_1980),
.B1(n_2003),
.B2(n_1981),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_L g2056 ( 
.A(n_2044),
.B(n_1809),
.Y(n_2056)
);

NAND3xp33_ASAP7_75t_L g2057 ( 
.A(n_2032),
.B(n_1996),
.C(n_1992),
.Y(n_2057)
);

A2O1A1Ixp33_ASAP7_75t_L g2058 ( 
.A1(n_2040),
.A2(n_1985),
.B(n_2001),
.C(n_2009),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2033),
.Y(n_2059)
);

O2A1O1Ixp33_ASAP7_75t_L g2060 ( 
.A1(n_2016),
.A2(n_2002),
.B(n_2000),
.C(n_1999),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2026),
.B(n_1981),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_2044),
.B(n_2001),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_2028),
.B(n_1934),
.Y(n_2063)
);

INVxp67_ASAP7_75t_L g2064 ( 
.A(n_2028),
.Y(n_2064)
);

OAI221xp5_ASAP7_75t_L g2065 ( 
.A1(n_2017),
.A2(n_2009),
.B1(n_1824),
.B2(n_1934),
.C(n_1964),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_SL g2066 ( 
.A1(n_2037),
.A2(n_1906),
.B1(n_1790),
.B2(n_1762),
.Y(n_2066)
);

AOI21xp33_ASAP7_75t_SL g2067 ( 
.A1(n_2027),
.A2(n_1730),
.B(n_1802),
.Y(n_2067)
);

INVxp33_ASAP7_75t_SL g2068 ( 
.A(n_2056),
.Y(n_2068)
);

INVxp67_ASAP7_75t_L g2069 ( 
.A(n_2056),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2045),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_2064),
.B(n_2041),
.Y(n_2071)
);

INVxp67_ASAP7_75t_L g2072 ( 
.A(n_2062),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2051),
.Y(n_2073)
);

AOI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_2053),
.A2(n_2029),
.B1(n_2038),
.B2(n_2042),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_2058),
.A2(n_2024),
.B1(n_2025),
.B2(n_2030),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_2062),
.B(n_2029),
.Y(n_2076)
);

INVxp67_ASAP7_75t_L g2077 ( 
.A(n_2053),
.Y(n_2077)
);

AOI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_2054),
.A2(n_2024),
.B(n_2034),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2052),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2059),
.Y(n_2080)
);

OAI221xp5_ASAP7_75t_L g2081 ( 
.A1(n_2046),
.A2(n_2035),
.B1(n_1915),
.B2(n_1897),
.C(n_1975),
.Y(n_2081)
);

OAI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_2055),
.A2(n_1788),
.B1(n_1910),
.B2(n_1852),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2072),
.B(n_2050),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2069),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2070),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2071),
.B(n_2063),
.Y(n_2086)
);

NAND3xp33_ASAP7_75t_L g2087 ( 
.A(n_2076),
.B(n_2047),
.C(n_2048),
.Y(n_2087)
);

OAI221xp5_ASAP7_75t_L g2088 ( 
.A1(n_2077),
.A2(n_2066),
.B1(n_2049),
.B2(n_2057),
.C(n_2065),
.Y(n_2088)
);

NOR2x1_ASAP7_75t_L g2089 ( 
.A(n_2078),
.B(n_2060),
.Y(n_2089)
);

AOI221xp5_ASAP7_75t_L g2090 ( 
.A1(n_2075),
.A2(n_2061),
.B1(n_2067),
.B2(n_1915),
.C(n_1897),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2074),
.B(n_1911),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2073),
.Y(n_2092)
);

NAND4xp25_ASAP7_75t_L g2093 ( 
.A(n_2068),
.B(n_1796),
.C(n_1756),
.D(n_1752),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_SL g2094 ( 
.A(n_2082),
.B(n_1774),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2079),
.B(n_1922),
.Y(n_2095)
);

NOR2x1_ASAP7_75t_L g2096 ( 
.A(n_2080),
.B(n_1730),
.Y(n_2096)
);

NAND4xp25_ASAP7_75t_L g2097 ( 
.A(n_2081),
.B(n_1741),
.C(n_1747),
.D(n_1970),
.Y(n_2097)
);

NOR2xp67_ASAP7_75t_L g2098 ( 
.A(n_2082),
.B(n_1960),
.Y(n_2098)
);

OAI221xp5_ASAP7_75t_L g2099 ( 
.A1(n_2089),
.A2(n_1970),
.B1(n_1966),
.B2(n_1946),
.C(n_1956),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2083),
.Y(n_2100)
);

NOR4xp75_ASAP7_75t_L g2101 ( 
.A(n_2088),
.B(n_1762),
.C(n_1851),
.D(n_1913),
.Y(n_2101)
);

OAI221xp5_ASAP7_75t_L g2102 ( 
.A1(n_2087),
.A2(n_1970),
.B1(n_1966),
.B2(n_1956),
.C(n_1949),
.Y(n_2102)
);

AOI222xp33_ASAP7_75t_L g2103 ( 
.A1(n_2091),
.A2(n_1964),
.B1(n_1966),
.B2(n_1956),
.C1(n_1949),
.C2(n_1947),
.Y(n_2103)
);

NOR3xp33_ASAP7_75t_L g2104 ( 
.A(n_2084),
.B(n_2086),
.C(n_2090),
.Y(n_2104)
);

AOI221xp5_ASAP7_75t_SL g2105 ( 
.A1(n_2097),
.A2(n_1949),
.B1(n_1947),
.B2(n_1946),
.C(n_1911),
.Y(n_2105)
);

OAI211xp5_ASAP7_75t_L g2106 ( 
.A1(n_2096),
.A2(n_1769),
.B(n_1946),
.C(n_1947),
.Y(n_2106)
);

AOI211xp5_ASAP7_75t_L g2107 ( 
.A1(n_2098),
.A2(n_1807),
.B(n_1783),
.C(n_1845),
.Y(n_2107)
);

AOI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_2094),
.A2(n_1888),
.B1(n_1783),
.B2(n_1872),
.Y(n_2108)
);

OAI22xp5_ASAP7_75t_L g2109 ( 
.A1(n_2100),
.A2(n_2108),
.B1(n_2098),
.B2(n_2104),
.Y(n_2109)
);

AOI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_2106),
.A2(n_2095),
.B1(n_2105),
.B2(n_2093),
.Y(n_2110)
);

AOI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_2107),
.A2(n_2092),
.B1(n_2085),
.B2(n_1929),
.Y(n_2111)
);

OAI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_2102),
.A2(n_1929),
.B(n_1922),
.Y(n_2112)
);

AOI221xp5_ASAP7_75t_L g2113 ( 
.A1(n_2099),
.A2(n_1911),
.B1(n_1852),
.B2(n_1816),
.C(n_1928),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_2103),
.A2(n_1926),
.B(n_1914),
.Y(n_2114)
);

AOI221x1_ASAP7_75t_SL g2115 ( 
.A1(n_2101),
.A2(n_1913),
.B1(n_1928),
.B2(n_1926),
.C(n_1914),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_2100),
.Y(n_2116)
);

NOR2x1_ASAP7_75t_L g2117 ( 
.A(n_2109),
.B(n_1922),
.Y(n_2117)
);

AND2x4_ASAP7_75t_L g2118 ( 
.A(n_2116),
.B(n_1922),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_2111),
.B(n_1922),
.Y(n_2119)
);

NOR2x1_ASAP7_75t_L g2120 ( 
.A(n_2112),
.B(n_2114),
.Y(n_2120)
);

INVxp67_ASAP7_75t_L g2121 ( 
.A(n_2110),
.Y(n_2121)
);

INVx1_ASAP7_75t_SL g2122 ( 
.A(n_2115),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_2118),
.B(n_1914),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2120),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2119),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2117),
.Y(n_2126)
);

NOR3x2_ASAP7_75t_L g2127 ( 
.A(n_2124),
.B(n_2121),
.C(n_2122),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_2126),
.A2(n_2113),
.B(n_1926),
.Y(n_2128)
);

AOI211xp5_ASAP7_75t_L g2129 ( 
.A1(n_2128),
.A2(n_2125),
.B(n_2123),
.C(n_1845),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_SL g2130 ( 
.A1(n_2129),
.A2(n_2125),
.B1(n_2127),
.B2(n_2123),
.Y(n_2130)
);

OAI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_2129),
.A2(n_1928),
.B1(n_1926),
.B2(n_1914),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2130),
.Y(n_2132)
);

AO22x1_ASAP7_75t_L g2133 ( 
.A1(n_2131),
.A2(n_1922),
.B1(n_1929),
.B2(n_1727),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2132),
.Y(n_2134)
);

AOI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_2133),
.A2(n_1928),
.B(n_1909),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2134),
.Y(n_2136)
);

O2A1O1Ixp33_ASAP7_75t_L g2137 ( 
.A1(n_2136),
.A2(n_2135),
.B(n_1711),
.C(n_1719),
.Y(n_2137)
);

BUFx2_ASAP7_75t_L g2138 ( 
.A(n_2137),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_2138),
.A2(n_1925),
.B1(n_1923),
.B2(n_1901),
.Y(n_2139)
);

AOI211xp5_ASAP7_75t_L g2140 ( 
.A1(n_2139),
.A2(n_1680),
.B(n_1925),
.C(n_1923),
.Y(n_2140)
);


endmodule