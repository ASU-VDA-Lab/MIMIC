module fake_jpeg_11619_n_508 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_508);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_508;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_51),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_62),
.Y(n_115)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_32),
.B(n_9),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_66),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_9),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_60),
.B(n_86),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_30),
.B(n_9),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_72),
.A2(n_37),
.B1(n_23),
.B2(n_44),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_36),
.B(n_8),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_36),
.B(n_8),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_18),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_7),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_96),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g143 ( 
.A(n_88),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_90),
.Y(n_133)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_93),
.A2(n_21),
.B1(n_17),
.B2(n_38),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_10),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

BUFx4f_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_105),
.B(n_124),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_106),
.A2(n_138),
.B1(n_140),
.B2(n_72),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_69),
.A2(n_34),
.B1(n_17),
.B2(n_21),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_116),
.A2(n_134),
.B1(n_70),
.B2(n_77),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_37),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_122),
.B(n_47),
.Y(n_175)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_51),
.A2(n_21),
.B1(n_17),
.B2(n_47),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_147),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_91),
.A2(n_41),
.B1(n_46),
.B2(n_26),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_55),
.Y(n_158)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_110),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_174),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_120),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_102),
.B(n_38),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_163),
.B(n_164),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_26),
.Y(n_164)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_166),
.Y(n_240)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_40),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_168),
.B(n_170),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_103),
.B(n_40),
.Y(n_170)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_22),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_173),
.B(n_179),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_175),
.B(n_191),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_176),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_22),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_104),
.Y(n_180)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_181),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_140),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_193),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_138),
.A2(n_94),
.B1(n_74),
.B2(n_90),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_188),
.A2(n_133),
.B1(n_137),
.B2(n_113),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_190),
.A2(n_203),
.B1(n_204),
.B2(n_206),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_27),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_192),
.A2(n_196),
.B1(n_199),
.B2(n_205),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_120),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_146),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_194),
.B(n_198),
.Y(n_219)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_106),
.A2(n_89),
.B1(n_79),
.B2(n_78),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

OR2x2_ASAP7_75t_SL g210 ( 
.A(n_197),
.B(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_109),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_45),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_202),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_118),
.B(n_45),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_127),
.B(n_42),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_113),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_117),
.A2(n_84),
.B1(n_82),
.B2(n_92),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_128),
.B1(n_109),
.B2(n_142),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_161),
.A2(n_165),
.B(n_173),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_211),
.A2(n_180),
.B(n_208),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_116),
.B1(n_134),
.B2(n_132),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_212),
.A2(n_243),
.B1(n_248),
.B2(n_48),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_170),
.A2(n_114),
.B(n_132),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_220),
.A2(n_184),
.B(n_185),
.Y(n_262)
);

OAI32xp33_ASAP7_75t_L g221 ( 
.A1(n_163),
.A2(n_153),
.A3(n_57),
.B1(n_61),
.B2(n_73),
.Y(n_221)
);

AOI32xp33_ASAP7_75t_L g277 ( 
.A1(n_221),
.A2(n_48),
.A3(n_35),
.B1(n_67),
.B2(n_29),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_231),
.B1(n_235),
.B2(n_241),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_187),
.A2(n_133),
.B1(n_137),
.B2(n_128),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_159),
.B(n_65),
.C(n_123),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_220),
.C(n_209),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_192),
.A2(n_123),
.B1(n_54),
.B2(n_63),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_196),
.A2(n_111),
.B1(n_125),
.B2(n_142),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_164),
.A2(n_41),
.B1(n_46),
.B2(n_125),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_204),
.A2(n_46),
.B1(n_111),
.B2(n_42),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_178),
.B1(n_207),
.B2(n_182),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_168),
.A2(n_46),
.B1(n_47),
.B2(n_35),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_186),
.B1(n_143),
.B2(n_145),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_179),
.A2(n_19),
.B1(n_27),
.B2(n_80),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_162),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_250),
.B(n_251),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_171),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_249),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_258),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_237),
.A2(n_205),
.B1(n_167),
.B2(n_172),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_254),
.A2(n_257),
.B1(n_264),
.B2(n_266),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_255),
.B(n_276),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_213),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_256),
.B(n_278),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_189),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_215),
.Y(n_259)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_259),
.Y(n_291)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_217),
.Y(n_260)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_262),
.A2(n_263),
.B(n_268),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_226),
.A2(n_166),
.B(n_199),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_237),
.A2(n_183),
.B1(n_181),
.B2(n_197),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_211),
.A2(n_200),
.B1(n_169),
.B2(n_208),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_219),
.A2(n_198),
.B(n_195),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_267),
.A2(n_280),
.B(n_236),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_169),
.B1(n_177),
.B2(n_176),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_272),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_270),
.A2(n_277),
.B1(n_281),
.B2(n_285),
.Y(n_290)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_177),
.Y(n_272)
);

OA21x2_ASAP7_75t_L g273 ( 
.A1(n_241),
.A2(n_101),
.B(n_143),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_273),
.B(n_274),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_235),
.A2(n_48),
.B1(n_35),
.B2(n_64),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_222),
.B(n_64),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_236),
.C(n_230),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_222),
.B(n_218),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_244),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_224),
.B(n_0),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_282),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_219),
.A2(n_0),
.B(n_1),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_227),
.A2(n_48),
.B1(n_35),
.B2(n_29),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_224),
.B(n_0),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_221),
.A2(n_48),
.B1(n_35),
.B2(n_29),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_284),
.Y(n_289)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_231),
.A2(n_3),
.B(n_29),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_279),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_299),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_319),
.Y(n_333)
);

AOI32xp33_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_210),
.A3(n_246),
.B1(n_234),
.B2(n_247),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_294),
.A2(n_273),
.B(n_286),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_298),
.B(n_245),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_282),
.Y(n_299)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_303),
.Y(n_322)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_269),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_313),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_230),
.C(n_223),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_223),
.C(n_245),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_267),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_307),
.B(n_310),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_285),
.A2(n_229),
.B1(n_210),
.B2(n_246),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_309),
.A2(n_320),
.B1(n_273),
.B2(n_254),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_256),
.B(n_240),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_251),
.B(n_250),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_312),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_271),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_258),
.B(n_240),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_321),
.Y(n_350)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_283),
.Y(n_316)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_316),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_252),
.A2(n_246),
.B1(n_214),
.B2(n_216),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_257),
.Y(n_321)
);

OAI32xp33_ASAP7_75t_L g323 ( 
.A1(n_296),
.A2(n_253),
.A3(n_268),
.B1(n_277),
.B2(n_262),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_323),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_325),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_301),
.A2(n_252),
.B1(n_278),
.B2(n_255),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_326),
.A2(n_329),
.B1(n_340),
.B2(n_309),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_287),
.B(n_275),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_330),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_301),
.A2(n_261),
.B1(n_270),
.B2(n_284),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_287),
.B(n_263),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_319),
.A2(n_280),
.B(n_264),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_332),
.A2(n_334),
.B(n_336),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_333),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_281),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_335),
.B(n_339),
.C(n_344),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_302),
.A2(n_273),
.B(n_261),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_292),
.Y(n_337)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_337),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_290),
.A2(n_286),
.B1(n_261),
.B2(n_274),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_338),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_289),
.A2(n_307),
.B1(n_305),
.B2(n_296),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_290),
.A2(n_286),
.B1(n_260),
.B2(n_283),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_341),
.A2(n_321),
.B1(n_317),
.B2(n_320),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_288),
.B(n_260),
.Y(n_342)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_342),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_299),
.B(n_225),
.Y(n_343)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_343),
.Y(n_370)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_291),
.Y(n_347)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_291),
.Y(n_348)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_348),
.Y(n_377)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_295),
.Y(n_349)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_349),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_308),
.B(n_225),
.C(n_216),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_297),
.C(n_304),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_228),
.Y(n_353)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_313),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_303),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_298),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_366),
.C(n_368),
.Y(n_391)
);

BUFx4f_ASAP7_75t_L g359 ( 
.A(n_354),
.Y(n_359)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_343),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_364),
.B(n_369),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_365),
.A2(n_378),
.B1(n_385),
.B2(n_346),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_306),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_331),
.B(n_311),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_328),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_371),
.A2(n_325),
.B1(n_341),
.B2(n_338),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_333),
.B(n_314),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_372),
.B(n_295),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_294),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_375),
.C(n_379),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_326),
.A2(n_340),
.B1(n_332),
.B2(n_329),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_314),
.Y(n_379)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_380),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_344),
.B(n_353),
.C(n_333),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_384),
.C(n_324),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_330),
.B(n_293),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_342),
.A2(n_317),
.B1(n_318),
.B2(n_297),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_386),
.A2(n_367),
.B1(n_362),
.B2(n_363),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_334),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_379),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_R g390 ( 
.A(n_357),
.B(n_384),
.C(n_370),
.Y(n_390)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_390),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_383),
.B(n_345),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_392),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_361),
.A2(n_350),
.B1(n_318),
.B2(n_336),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_393),
.A2(n_397),
.B1(n_404),
.B2(n_406),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_351),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_394),
.B(n_403),
.Y(n_423)
);

AO21x1_ASAP7_75t_L g395 ( 
.A1(n_378),
.A2(n_323),
.B(n_348),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_395),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_361),
.A2(n_349),
.B1(n_347),
.B2(n_322),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_408),
.C(n_411),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_324),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_399),
.Y(n_415)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_400),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_322),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_401),
.A2(n_407),
.B1(n_7),
.B2(n_11),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_402),
.B(n_29),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_242),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_373),
.B(n_346),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_373),
.B(n_316),
.C(n_337),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_409),
.A2(n_410),
.B1(n_412),
.B2(n_382),
.Y(n_427)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_359),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_374),
.B(n_292),
.C(n_228),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_367),
.A2(n_300),
.B1(n_228),
.B2(n_217),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_417),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_389),
.B(n_366),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_414),
.B(n_416),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_381),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_372),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_356),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_429),
.Y(n_442)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_425),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_395),
.A2(n_362),
.B1(n_371),
.B2(n_363),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_426),
.A2(n_407),
.B1(n_401),
.B2(n_392),
.Y(n_437)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_427),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_355),
.C(n_217),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_433),
.C(n_387),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_300),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_405),
.A2(n_242),
.B(n_4),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_400),
.C(n_387),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_432),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_24),
.C(n_3),
.Y(n_433)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_422),
.Y(n_435)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_435),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_418),
.B(n_388),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_436),
.B(n_446),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_450),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_411),
.C(n_401),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_444),
.B(n_447),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_423),
.B(n_399),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_402),
.C(n_410),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_415),
.Y(n_448)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_448),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_449),
.B(n_433),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_413),
.B(n_390),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_451),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g452 ( 
.A1(n_420),
.A2(n_412),
.B1(n_7),
.B2(n_11),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_452),
.A2(n_432),
.B(n_431),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_419),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_465),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_434),
.Y(n_459)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_459),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_447),
.B(n_424),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_442),
.Y(n_472)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_443),
.Y(n_463)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_463),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_439),
.B(n_420),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_464),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_425),
.Y(n_466)
);

OAI21x1_ASAP7_75t_L g471 ( 
.A1(n_466),
.A2(n_459),
.B(n_464),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_468),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_414),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_453),
.A2(n_441),
.B(n_416),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_469),
.A2(n_479),
.B(n_438),
.Y(n_487)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_471),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_472),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_442),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_476),
.Y(n_486)
);

AO21x1_ASAP7_75t_L g475 ( 
.A1(n_462),
.A2(n_452),
.B(n_445),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_475),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_429),
.Y(n_476)
);

AO21x1_ASAP7_75t_L g477 ( 
.A1(n_462),
.A2(n_454),
.B(n_455),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_SL g490 ( 
.A1(n_477),
.A2(n_467),
.B(n_445),
.C(n_468),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_SL g479 ( 
.A(n_461),
.B(n_417),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_438),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_481),
.B(n_480),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_477),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_485),
.B(n_488),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_487),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_482),
.B(n_454),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_490),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_491),
.B(n_492),
.C(n_470),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_478),
.A2(n_11),
.B(n_12),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_485),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_474),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_497),
.A2(n_498),
.B(n_475),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_483),
.A2(n_481),
.B(n_480),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_495),
.B(n_484),
.C(n_489),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_499),
.B(n_501),
.C(n_502),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_500),
.A2(n_496),
.B(n_490),
.Y(n_504)
);

BUFx24_ASAP7_75t_SL g502 ( 
.A(n_494),
.Y(n_502)
);

OAI321xp33_ASAP7_75t_L g505 ( 
.A1(n_504),
.A2(n_12),
.A3(n_13),
.B1(n_15),
.B2(n_24),
.C(n_3),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_505),
.A2(n_503),
.B(n_13),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_506),
.A2(n_12),
.B1(n_15),
.B2(n_24),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_507),
.B(n_24),
.Y(n_508)
);


endmodule