module fake_jpeg_20345_n_290 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_290);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVxp67_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_6),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_20),
.B1(n_25),
.B2(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_20),
.B1(n_23),
.B2(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_31),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_60),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_39),
.B1(n_43),
.B2(n_36),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_60),
.Y(n_83)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_78),
.B1(n_82),
.B2(n_86),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_22),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_13),
.C(n_22),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_36),
.B1(n_43),
.B2(n_39),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_39),
.B1(n_27),
.B2(n_45),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_39),
.B1(n_27),
.B2(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_80),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_36),
.B1(n_38),
.B2(n_41),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_66),
.B1(n_78),
.B2(n_75),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_59),
.B1(n_47),
.B2(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_90),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_49),
.B(n_61),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_105),
.B(n_12),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_41),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_86),
.A2(n_50),
.B1(n_64),
.B2(n_62),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_92),
.B1(n_107),
.B2(n_73),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_50),
.B1(n_53),
.B2(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_96),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_13),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_87),
.C(n_85),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_48),
.C(n_29),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_101),
.A2(n_74),
.B1(n_68),
.B2(n_73),
.Y(n_116)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_21),
.B(n_8),
.Y(n_105)
);

XOR2x1_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_75),
.Y(n_108)
);

XNOR2x1_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_118),
.Y(n_150)
);

BUFx8_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_115),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_21),
.B1(n_20),
.B2(n_74),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_128),
.B1(n_18),
.B2(n_28),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_113),
.A2(n_121),
.B1(n_18),
.B2(n_16),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_117),
.Y(n_151)
);

AO22x1_ASAP7_75t_SL g117 ( 
.A1(n_106),
.A2(n_29),
.B1(n_26),
.B2(n_34),
.Y(n_117)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_98),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_119),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_32),
.A3(n_30),
.B1(n_28),
.B2(n_26),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_68),
.B1(n_23),
.B2(n_30),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_106),
.A2(n_32),
.B1(n_26),
.B2(n_29),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_28),
.B1(n_69),
.B2(n_70),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_92),
.B1(n_107),
.B2(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_89),
.A2(n_16),
.B(n_70),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_107),
.B(n_96),
.Y(n_144)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_134),
.B(n_136),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_100),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_139),
.C(n_141),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_100),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_90),
.C(n_101),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_153),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_108),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_149),
.C(n_124),
.Y(n_176)
);

AOI21x1_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_88),
.B(n_93),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_146),
.A2(n_150),
.B1(n_6),
.B2(n_10),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_70),
.B(n_93),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_154),
.B(n_120),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_18),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_152),
.A2(n_163),
.B1(n_129),
.B2(n_126),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_69),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_9),
.B(n_11),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_69),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_159),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_114),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_113),
.A2(n_23),
.B1(n_18),
.B2(n_19),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_161),
.Y(n_185)
);

AO22x1_ASAP7_75t_SL g162 ( 
.A1(n_117),
.A2(n_24),
.B1(n_19),
.B2(n_16),
.Y(n_162)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_131),
.B1(n_127),
.B2(n_114),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_165),
.A2(n_172),
.B1(n_173),
.B2(n_162),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_166),
.A2(n_177),
.B(n_162),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_188),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_147),
.B(n_115),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_170),
.B(n_180),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_127),
.B1(n_117),
.B2(n_119),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_124),
.B1(n_109),
.B2(n_24),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_145),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_109),
.B(n_7),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_6),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_24),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_186),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_135),
.A2(n_6),
.B(n_10),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_5),
.B1(n_10),
.B2(n_9),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_163),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_138),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_156),
.A2(n_144),
.B1(n_140),
.B2(n_142),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_0),
.C(n_1),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_154),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_148),
.B(n_158),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_177),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_194),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_176),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_168),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_197),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_137),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_152),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_189),
.B(n_146),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_203),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_209),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_0),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_211),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_184),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_188),
.C(n_184),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_212),
.B(n_215),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_183),
.C(n_164),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_205),
.B(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_191),
.A2(n_185),
.B1(n_178),
.B2(n_167),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_226),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_190),
.A2(n_185),
.B1(n_178),
.B2(n_167),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_179),
.B1(n_169),
.B2(n_172),
.Y(n_228)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

BUFx24_ASAP7_75t_SL g230 ( 
.A(n_224),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_238),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_193),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_225),
.Y(n_244)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_237),
.Y(n_252)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_243),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_197),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_192),
.B(n_202),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_210),
.B(n_179),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_207),
.B1(n_204),
.B2(n_203),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_201),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_221),
.B1(n_213),
.B2(n_229),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_248),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_225),
.C(n_215),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_246),
.B(n_250),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_233),
.B1(n_229),
.B2(n_199),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_223),
.C(n_220),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_223),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_251),
.B(n_254),
.Y(n_266)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_243),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_181),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_246),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_234),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_262),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_211),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_251),
.B1(n_3),
.B2(n_4),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_250),
.A2(n_3),
.B(n_4),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_265),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_3),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_267),
.B(n_5),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_264),
.B(n_254),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_271),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_270),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_258),
.B(n_3),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_4),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_2),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_273),
.A2(n_266),
.B(n_261),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_276),
.A2(n_273),
.B(n_7),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_275),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_281),
.C(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_283),
.A2(n_278),
.B(n_277),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_285),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_286),
.B(n_284),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_7),
.B(n_8),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_2),
.B1(n_11),
.B2(n_209),
.Y(n_290)
);


endmodule