module fake_netlist_6_1816_n_1065 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1065);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1065;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_760;
wire n_741;
wire n_680;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_832;
wire n_280;
wire n_287;
wire n_685;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_222;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_989;
wire n_843;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_962;
wire n_824;
wire n_1000;
wire n_279;
wire n_796;
wire n_686;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_984;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_939;
wire n_819;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_964;
wire n_802;
wire n_982;
wire n_831;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g190 ( 
.A(n_76),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_73),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_98),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_122),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_68),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_120),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_88),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_61),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_16),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_159),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_173),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_43),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_54),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_179),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_36),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_48),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_5),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_9),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_106),
.Y(n_213)
);

BUFx8_ASAP7_75t_SL g214 ( 
.A(n_186),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_123),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_143),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_67),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_18),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_69),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_72),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_175),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_117),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_56),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_104),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_70),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_126),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_119),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_14),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_52),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_74),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_165),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_51),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_89),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_62),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_7),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_35),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_181),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_95),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_114),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_118),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_169),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_34),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_50),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_105),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_59),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_184),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_183),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_155),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_141),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_100),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_23),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_29),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_25),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_41),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_180),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_176),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_134),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_46),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_212),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_208),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_211),
.Y(n_264)
);

BUFx2_ASAP7_75t_SL g265 ( 
.A(n_227),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_217),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_209),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_193),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_192),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

INVxp33_ASAP7_75t_SL g273 ( 
.A(n_200),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_190),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_191),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_193),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g278 ( 
.A(n_214),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_210),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_196),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_228),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_196),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_229),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_240),
.Y(n_285)
);

INVxp33_ASAP7_75t_SL g286 ( 
.A(n_253),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_227),
.Y(n_287)
);

INVxp33_ASAP7_75t_SL g288 ( 
.A(n_194),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_195),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_256),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_234),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_239),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_256),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_242),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_240),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_240),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_257),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_224),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_224),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_231),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_255),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_255),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_216),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_241),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_198),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_197),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_199),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_249),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_269),
.Y(n_312)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_263),
.A2(n_202),
.B(n_201),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_263),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_285),
.A2(n_231),
.B1(n_244),
.B2(n_250),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_268),
.Y(n_317)
);

BUFx8_ASAP7_75t_SL g318 ( 
.A(n_287),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_271),
.B(n_203),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_280),
.Y(n_322)
);

OAI22x1_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_236),
.B1(n_248),
.B2(n_252),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_260),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_270),
.B(n_249),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

AND2x6_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_30),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_264),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_274),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_266),
.A2(n_244),
.B1(n_250),
.B2(n_254),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_289),
.B(n_307),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_285),
.A2(n_296),
.B1(n_273),
.B2(n_286),
.Y(n_332)
);

OA21x2_ASAP7_75t_L g333 ( 
.A1(n_274),
.A2(n_276),
.B(n_275),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_275),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_262),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_276),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_279),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_299),
.B(n_258),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_296),
.A2(n_247),
.B1(n_246),
.B2(n_245),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_283),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_284),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_284),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_290),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_290),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_292),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_292),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_308),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_291),
.B(n_204),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_293),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_301),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_291),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_267),
.A2(n_243),
.B1(n_238),
.B2(n_237),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_265),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_298),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_281),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_295),
.B(n_206),
.Y(n_361)
);

AND2x6_ASAP7_75t_L g362 ( 
.A(n_297),
.B(n_31),
.Y(n_362)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_297),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_322),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_R g365 ( 
.A(n_355),
.B(n_297),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_R g366 ( 
.A(n_355),
.B(n_207),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_318),
.Y(n_367)
);

BUFx10_ASAP7_75t_L g368 ( 
.A(n_328),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_310),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_288),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_322),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_318),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_358),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_310),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_310),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_R g376 ( 
.A(n_331),
.B(n_213),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_358),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_R g378 ( 
.A(n_321),
.B(n_215),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_330),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_357),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_340),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_335),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_360),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_310),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_341),
.B(n_261),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_332),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_316),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_334),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_309),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_311),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_319),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_323),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_346),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_339),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_348),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_323),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_325),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_R g400 ( 
.A(n_340),
.B(n_219),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_325),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_352),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_361),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_337),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_278),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_361),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_351),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_313),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_353),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_313),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_353),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_313),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_337),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_R g417 ( 
.A(n_340),
.B(n_220),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_363),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_333),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_R g420 ( 
.A(n_333),
.B(n_0),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_363),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_R g422 ( 
.A(n_356),
.B(n_221),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_356),
.B(n_280),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_363),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_363),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_326),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_337),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_326),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_356),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_362),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_319),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_333),
.Y(n_432)
);

BUFx10_ASAP7_75t_L g433 ( 
.A(n_367),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_423),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_432),
.A2(n_265),
.B1(n_223),
.B2(n_225),
.Y(n_435)
);

AND2x2_ASAP7_75t_SL g436 ( 
.A(n_390),
.B(n_282),
.Y(n_436)
);

OR2x6_ASAP7_75t_L g437 ( 
.A(n_388),
.B(n_277),
.Y(n_437)
);

OR2x6_ASAP7_75t_L g438 ( 
.A(n_385),
.B(n_414),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_389),
.B(n_342),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g440 ( 
.A(n_429),
.B(n_362),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_423),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_423),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_426),
.Y(n_443)
);

AND2x4_ASAP7_75t_SL g444 ( 
.A(n_368),
.B(n_282),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_429),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_364),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_394),
.B(n_336),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_381),
.B(n_342),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_419),
.B(n_342),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_396),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_404),
.B(n_342),
.Y(n_454)
);

OAI22x1_ASAP7_75t_L g455 ( 
.A1(n_379),
.A2(n_303),
.B1(n_302),
.B2(n_305),
.Y(n_455)
);

AND2x2_ASAP7_75t_SL g456 ( 
.A(n_401),
.B(n_294),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_407),
.B(n_345),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_365),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_391),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_409),
.B(n_277),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_391),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_403),
.B(n_222),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_428),
.B(n_345),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_399),
.B(n_232),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_372),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_366),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_392),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_411),
.B(n_413),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_376),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_398),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_398),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_431),
.B(n_336),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_378),
.B(n_345),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_369),
.Y(n_474)
);

OR2x6_ASAP7_75t_L g475 ( 
.A(n_406),
.B(n_294),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_369),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_418),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_368),
.B(n_262),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_370),
.B(n_345),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_374),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_383),
.B(n_302),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_374),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_375),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_408),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_373),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_377),
.B(n_350),
.Y(n_488)
);

CKINVDCx6p67_ASAP7_75t_R g489 ( 
.A(n_386),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_395),
.B(n_233),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_416),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_427),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_412),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_393),
.B(n_303),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_415),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_430),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_424),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_397),
.B(n_329),
.Y(n_499)
);

BUFx4f_ASAP7_75t_L g500 ( 
.A(n_421),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_425),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_387),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_420),
.B(n_362),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_380),
.B(n_304),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_400),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_481),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_460),
.B(n_304),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_499),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_434),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_502),
.A2(n_305),
.B1(n_420),
.B2(n_298),
.Y(n_510)
);

A2O1A1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_439),
.A2(n_315),
.B(n_338),
.C(n_359),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_434),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_478),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_329),
.Y(n_514)
);

OAI221xp5_ASAP7_75t_L g515 ( 
.A1(n_448),
.A2(n_300),
.B1(n_359),
.B2(n_338),
.C(n_349),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_443),
.B(n_417),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_442),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_442),
.Y(n_518)
);

NAND2x1p5_ASAP7_75t_L g519 ( 
.A(n_443),
.B(n_324),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_436),
.B(n_343),
.Y(n_520)
);

AO22x2_ASAP7_75t_L g521 ( 
.A1(n_493),
.A2(n_300),
.B1(n_1),
.B2(n_2),
.Y(n_521)
);

OAI221xp5_ASAP7_75t_L g522 ( 
.A1(n_494),
.A2(n_349),
.B1(n_344),
.B2(n_347),
.C(n_343),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_441),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_453),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_472),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_504),
.B(n_344),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_472),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_485),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_468),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_469),
.Y(n_530)
);

OR2x2_ASAP7_75t_SL g531 ( 
.A(n_496),
.B(n_347),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_485),
.Y(n_532)
);

BUFx8_ASAP7_75t_L g533 ( 
.A(n_487),
.Y(n_533)
);

A2O1A1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_462),
.A2(n_315),
.B(n_312),
.C(n_320),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_467),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_503),
.B(n_327),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_486),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_449),
.B(n_327),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_471),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_471),
.Y(n_540)
);

AO22x2_ASAP7_75t_L g541 ( 
.A1(n_497),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_486),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_466),
.Y(n_543)
);

CKINVDCx14_ASAP7_75t_R g544 ( 
.A(n_465),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_503),
.B(n_327),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_456),
.B(n_422),
.Y(n_546)
);

NAND2x1p5_ASAP7_75t_L g547 ( 
.A(n_445),
.B(n_324),
.Y(n_547)
);

NAND3x1_ASAP7_75t_L g548 ( 
.A(n_495),
.B(n_315),
.C(n_324),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_491),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_444),
.B(n_314),
.Y(n_550)
);

OAI221xp5_ASAP7_75t_L g551 ( 
.A1(n_446),
.A2(n_320),
.B1(n_317),
.B2(n_314),
.C(n_326),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_449),
.B(n_317),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_468),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_489),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_452),
.B(n_32),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_482),
.Y(n_556)
);

AO22x2_ASAP7_75t_L g557 ( 
.A1(n_497),
.A2(n_435),
.B1(n_505),
.B2(n_447),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_482),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_437),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_491),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_453),
.B(n_319),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_451),
.B(n_33),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_458),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_464),
.B(n_3),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_437),
.Y(n_565)
);

AO22x2_ASAP7_75t_L g566 ( 
.A1(n_498),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_520),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_533),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_514),
.B(n_453),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_524),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_508),
.B(n_475),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_538),
.B(n_498),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_535),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_533),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_562),
.A2(n_450),
.B(n_479),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_529),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_506),
.B(n_475),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_526),
.B(n_500),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_524),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_510),
.A2(n_455),
.B1(n_454),
.B2(n_457),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_539),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_507),
.B(n_500),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_536),
.A2(n_463),
.B(n_473),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_524),
.B(n_501),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_564),
.B(n_488),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_528),
.B(n_501),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_553),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_517),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_518),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_562),
.A2(n_484),
.B(n_476),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_510),
.B(n_477),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_546),
.B(n_477),
.Y(n_592)
);

BUFx6f_ASAP7_75t_SL g593 ( 
.A(n_565),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_545),
.A2(n_483),
.B(n_459),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_532),
.B(n_484),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_563),
.B(n_438),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_509),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_537),
.B(n_459),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_540),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_552),
.B(n_483),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_511),
.A2(n_440),
.B(n_461),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_542),
.B(n_470),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_556),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_525),
.A2(n_492),
.B1(n_440),
.B2(n_438),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_555),
.A2(n_527),
.B1(n_557),
.B2(n_523),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_550),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_549),
.B(n_474),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_560),
.B(n_480),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_513),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_552),
.B(n_440),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_555),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_530),
.B(n_478),
.Y(n_612)
);

O2A1O1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_516),
.A2(n_522),
.B(n_515),
.C(n_534),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_513),
.B(n_433),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_561),
.A2(n_38),
.B(n_37),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_512),
.A2(n_40),
.B(n_39),
.Y(n_616)
);

INVx11_ASAP7_75t_L g617 ( 
.A(n_544),
.Y(n_617)
);

AO21x1_ASAP7_75t_L g618 ( 
.A1(n_558),
.A2(n_519),
.B(n_547),
.Y(n_618)
);

OAI21x1_ASAP7_75t_L g619 ( 
.A1(n_548),
.A2(n_44),
.B(n_42),
.Y(n_619)
);

NAND2x1p5_ASAP7_75t_L g620 ( 
.A(n_570),
.B(n_513),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_567),
.B(n_557),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_573),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_588),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_617),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_587),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_578),
.B(n_543),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_567),
.B(n_559),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_606),
.B(n_521),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_611),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_589),
.Y(n_630)
);

A2O1A1Ixp33_ASAP7_75t_SL g631 ( 
.A1(n_613),
.A2(n_522),
.B(n_515),
.C(n_551),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_571),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_611),
.A2(n_531),
.B1(n_566),
.B2(n_541),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_606),
.B(n_554),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_582),
.B(n_433),
.Y(n_635)
);

AND2x2_ASAP7_75t_SL g636 ( 
.A(n_605),
.B(n_566),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_577),
.A2(n_541),
.B1(n_521),
.B2(n_7),
.Y(n_637)
);

INVx3_ASAP7_75t_SL g638 ( 
.A(n_587),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_611),
.B(n_4),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_581),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_580),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_641)
);

A2O1A1Ixp33_ASAP7_75t_SL g642 ( 
.A1(n_601),
.A2(n_112),
.B(n_188),
.C(n_187),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_SL g643 ( 
.A1(n_580),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_643)
);

O2A1O1Ixp33_ASAP7_75t_L g644 ( 
.A1(n_591),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_585),
.B(n_586),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_605),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_587),
.B(n_45),
.Y(n_647)
);

NAND3xp33_ASAP7_75t_L g648 ( 
.A(n_569),
.B(n_13),
.C(n_14),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_575),
.A2(n_116),
.B(n_185),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_599),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_612),
.B(n_15),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_596),
.B(n_15),
.Y(n_652)
);

AND2x4_ASAP7_75t_SL g653 ( 
.A(n_570),
.B(n_47),
.Y(n_653)
);

O2A1O1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_592),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_654)
);

O2A1O1Ixp33_ASAP7_75t_L g655 ( 
.A1(n_584),
.A2(n_17),
.B(n_19),
.C(n_20),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_614),
.B(n_19),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_568),
.B(n_49),
.Y(n_657)
);

INVx5_ASAP7_75t_L g658 ( 
.A(n_572),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_603),
.B(n_20),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_604),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_572),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_583),
.A2(n_129),
.B(n_182),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_576),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_597),
.B(n_24),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_574),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_610),
.B(n_25),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_572),
.B(n_26),
.Y(n_667)
);

OAI22xp33_ASAP7_75t_L g668 ( 
.A1(n_609),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_597),
.B(n_27),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_602),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_607),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_608),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_595),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_598),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_600),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_590),
.A2(n_131),
.B(n_53),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_593),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_638),
.Y(n_678)
);

CKINVDCx11_ASAP7_75t_R g679 ( 
.A(n_625),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_625),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_658),
.B(n_572),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_623),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_630),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_658),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_625),
.Y(n_685)
);

BUFx2_ASAP7_75t_SL g686 ( 
.A(n_658),
.Y(n_686)
);

CKINVDCx11_ASAP7_75t_R g687 ( 
.A(n_657),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_622),
.Y(n_688)
);

BUFx8_ASAP7_75t_L g689 ( 
.A(n_651),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_621),
.Y(n_690)
);

NAND2x1p5_ASAP7_75t_L g691 ( 
.A(n_629),
.B(n_579),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_650),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_640),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_620),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_629),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_672),
.Y(n_696)
);

INVx3_ASAP7_75t_SL g697 ( 
.A(n_624),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_645),
.B(n_579),
.Y(n_698)
);

BUFx6f_ASAP7_75t_SL g699 ( 
.A(n_657),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_673),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_647),
.Y(n_701)
);

CKINVDCx8_ASAP7_75t_R g702 ( 
.A(n_665),
.Y(n_702)
);

INVx5_ASAP7_75t_L g703 ( 
.A(n_647),
.Y(n_703)
);

BUFx6f_ASAP7_75t_SL g704 ( 
.A(n_675),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_674),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_653),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_677),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_670),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_627),
.Y(n_709)
);

INVx8_ASAP7_75t_L g710 ( 
.A(n_663),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_626),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_671),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_632),
.B(n_615),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_634),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_659),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_635),
.B(n_616),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_628),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_667),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_633),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_636),
.B(n_619),
.Y(n_720)
);

INVx5_ASAP7_75t_L g721 ( 
.A(n_642),
.Y(n_721)
);

BUFx12f_ASAP7_75t_L g722 ( 
.A(n_656),
.Y(n_722)
);

BUFx4_ASAP7_75t_SL g723 ( 
.A(n_648),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_664),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_666),
.Y(n_725)
);

NAND2x1p5_ASAP7_75t_L g726 ( 
.A(n_641),
.B(n_639),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_652),
.Y(n_727)
);

BUFx10_ASAP7_75t_L g728 ( 
.A(n_654),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_669),
.B(n_594),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_643),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_646),
.Y(n_731)
);

INVxp67_ASAP7_75t_SL g732 ( 
.A(n_643),
.Y(n_732)
);

INVxp67_ASAP7_75t_SL g733 ( 
.A(n_644),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_660),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_637),
.B(n_28),
.Y(n_735)
);

BUFx2_ASAP7_75t_SL g736 ( 
.A(n_662),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_661),
.B(n_55),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_655),
.Y(n_738)
);

BUFx12f_ASAP7_75t_L g739 ( 
.A(n_668),
.Y(n_739)
);

BUFx4f_ASAP7_75t_SL g740 ( 
.A(n_649),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_702),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_732),
.A2(n_730),
.B1(n_703),
.B2(n_701),
.Y(n_742)
);

OAI21x1_ASAP7_75t_SL g743 ( 
.A1(n_712),
.A2(n_618),
.B(n_676),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_682),
.Y(n_744)
);

OAI21x1_ASAP7_75t_L g745 ( 
.A1(n_683),
.A2(n_631),
.B(n_593),
.Y(n_745)
);

OAI21x1_ASAP7_75t_L g746 ( 
.A1(n_683),
.A2(n_57),
.B(n_58),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_701),
.B(n_60),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_708),
.A2(n_63),
.B(n_64),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_716),
.A2(n_65),
.B(n_66),
.Y(n_749)
);

AO31x2_ASAP7_75t_L g750 ( 
.A1(n_738),
.A2(n_71),
.A3(n_75),
.B(n_77),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_701),
.B(n_78),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_701),
.B(n_79),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_708),
.B(n_80),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_690),
.B(n_81),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_700),
.A2(n_82),
.B(n_83),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_714),
.B(n_84),
.Y(n_756)
);

BUFx8_ASAP7_75t_L g757 ( 
.A(n_699),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_684),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_703),
.B(n_85),
.Y(n_759)
);

OAI21x1_ASAP7_75t_L g760 ( 
.A1(n_700),
.A2(n_86),
.B(n_87),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_698),
.A2(n_90),
.B(n_91),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_690),
.B(n_92),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_692),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_696),
.Y(n_764)
);

AO21x2_ASAP7_75t_L g765 ( 
.A1(n_733),
.A2(n_93),
.B(n_94),
.Y(n_765)
);

NAND3xp33_ASAP7_75t_L g766 ( 
.A(n_732),
.B(n_96),
.C(n_97),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_717),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_717),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_703),
.B(n_712),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_705),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_713),
.A2(n_99),
.B(n_101),
.Y(n_771)
);

AO21x2_ASAP7_75t_L g772 ( 
.A1(n_733),
.A2(n_103),
.B(n_107),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_711),
.B(n_108),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_693),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_695),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_724),
.B(n_109),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_698),
.A2(n_110),
.B(n_111),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_739),
.A2(n_113),
.B1(n_115),
.B2(n_121),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_727),
.B(n_718),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_725),
.A2(n_124),
.B(n_125),
.Y(n_780)
);

OAI21x1_ASAP7_75t_L g781 ( 
.A1(n_725),
.A2(n_127),
.B(n_128),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_718),
.Y(n_782)
);

AOI21x1_ASAP7_75t_L g783 ( 
.A1(n_729),
.A2(n_130),
.B(n_132),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_715),
.B(n_133),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_688),
.Y(n_785)
);

OA21x2_ASAP7_75t_L g786 ( 
.A1(n_729),
.A2(n_720),
.B(n_734),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_695),
.Y(n_787)
);

NAND4xp25_ASAP7_75t_L g788 ( 
.A(n_735),
.B(n_135),
.C(n_136),
.D(n_137),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_704),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_719),
.B(n_138),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_721),
.A2(n_139),
.B(n_140),
.Y(n_791)
);

OA21x2_ASAP7_75t_L g792 ( 
.A1(n_729),
.A2(n_142),
.B(n_144),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_704),
.Y(n_793)
);

OAI21x1_ASAP7_75t_SL g794 ( 
.A1(n_731),
.A2(n_145),
.B(n_147),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_768),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_749),
.A2(n_726),
.B(n_737),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_763),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_768),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_744),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_786),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_786),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_774),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_785),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_769),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_764),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_782),
.B(n_727),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_757),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_779),
.B(n_709),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_770),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_788),
.A2(n_739),
.B1(n_726),
.B2(n_740),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_767),
.Y(n_811)
);

INVxp33_ASAP7_75t_L g812 ( 
.A(n_773),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_775),
.B(n_734),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_787),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_745),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_754),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_754),
.B(n_688),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_792),
.B(n_721),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_792),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_750),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_750),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_750),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_753),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_753),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_778),
.A2(n_699),
.B1(n_740),
.B2(n_722),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_748),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_769),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_765),
.Y(n_828)
);

AO21x1_ASAP7_75t_L g829 ( 
.A1(n_742),
.A2(n_723),
.B(n_684),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_758),
.Y(n_830)
);

AO21x2_ASAP7_75t_L g831 ( 
.A1(n_743),
.A2(n_721),
.B(n_736),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_742),
.Y(n_832)
);

OAI21x1_ASAP7_75t_L g833 ( 
.A1(n_783),
.A2(n_691),
.B(n_721),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_778),
.A2(n_703),
.B1(n_722),
.B2(n_706),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_765),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_772),
.Y(n_836)
);

AO21x1_ASAP7_75t_SL g837 ( 
.A1(n_777),
.A2(n_723),
.B(n_728),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_757),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_789),
.B(n_793),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_772),
.B(n_790),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_788),
.A2(n_728),
.B1(n_687),
.B2(n_689),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_816),
.B(n_761),
.Y(n_842)
);

OR2x6_ASAP7_75t_L g843 ( 
.A(n_800),
.B(n_791),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_823),
.B(n_761),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_807),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_808),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_807),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_800),
.B(n_762),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_823),
.B(n_756),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_841),
.A2(n_766),
.B1(n_777),
.B2(n_790),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_800),
.B(n_771),
.Y(n_851)
);

AND2x2_ASAP7_75t_SL g852 ( 
.A(n_840),
.B(n_747),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_805),
.Y(n_853)
);

CKINVDCx16_ASAP7_75t_R g854 ( 
.A(n_838),
.Y(n_854)
);

NAND2xp33_ASAP7_75t_R g855 ( 
.A(n_839),
.B(n_747),
.Y(n_855)
);

BUFx12f_ASAP7_75t_L g856 ( 
.A(n_838),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_802),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_837),
.A2(n_766),
.B1(n_728),
.B2(n_687),
.Y(n_858)
);

OR2x6_ASAP7_75t_L g859 ( 
.A(n_815),
.B(n_791),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_802),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_795),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_801),
.B(n_776),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_839),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_799),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_R g865 ( 
.A(n_804),
.B(n_741),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_SL g866 ( 
.A1(n_796),
.A2(n_749),
.B1(n_752),
.B2(n_751),
.Y(n_866)
);

NOR3xp33_ASAP7_75t_SL g867 ( 
.A(n_834),
.B(n_689),
.C(n_702),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_799),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_805),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_804),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_810),
.A2(n_759),
.B(n_751),
.C(n_752),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_825),
.A2(n_759),
.B(n_746),
.C(n_781),
.Y(n_872)
);

AO21x2_ASAP7_75t_L g873 ( 
.A1(n_828),
.A2(n_794),
.B(n_780),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_870),
.B(n_801),
.Y(n_874)
);

AND2x4_ASAP7_75t_SL g875 ( 
.A(n_867),
.B(n_827),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_857),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_870),
.B(n_839),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_861),
.B(n_798),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_857),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_848),
.B(n_803),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_848),
.B(n_804),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_856),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_851),
.B(n_815),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_850),
.A2(n_837),
.B1(n_829),
.B2(n_812),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_860),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_862),
.B(n_806),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_860),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_851),
.B(n_827),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_862),
.B(n_806),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_863),
.B(n_811),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_864),
.B(n_820),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_864),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_868),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_863),
.B(n_811),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_853),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_868),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_884),
.A2(n_858),
.B(n_871),
.C(n_866),
.Y(n_897)
);

OAI211xp5_ASAP7_75t_L g898 ( 
.A1(n_878),
.A2(n_849),
.B(n_842),
.C(n_844),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_881),
.B(n_863),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_891),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_881),
.B(n_863),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_880),
.B(n_846),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_895),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_895),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_891),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_890),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_882),
.A2(n_871),
.B(n_872),
.C(n_840),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_878),
.Y(n_908)
);

NAND4xp25_ASAP7_75t_L g909 ( 
.A(n_882),
.B(n_817),
.C(n_832),
.D(n_845),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_886),
.B(n_889),
.Y(n_910)
);

NOR3xp33_ASAP7_75t_L g911 ( 
.A(n_882),
.B(n_854),
.C(n_872),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_903),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_906),
.B(n_888),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_904),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_SL g915 ( 
.A(n_907),
.B(n_856),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_910),
.B(n_888),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_908),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_911),
.B(n_875),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_899),
.B(n_888),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_900),
.Y(n_920)
);

AOI221xp5_ASAP7_75t_SL g921 ( 
.A1(n_897),
.A2(n_909),
.B1(n_902),
.B2(n_911),
.C(n_890),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_900),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_901),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_923),
.B(n_898),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_921),
.B(n_905),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_915),
.B(n_865),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_920),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_919),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_912),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_919),
.B(n_888),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_914),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_925),
.A2(n_926),
.B(n_918),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_928),
.B(n_918),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_930),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_925),
.B(n_917),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_927),
.B(n_924),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_929),
.B(n_922),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_931),
.B(n_918),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_938),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_933),
.B(n_916),
.Y(n_940)
);

OAI221xp5_ASAP7_75t_L g941 ( 
.A1(n_932),
.A2(n_847),
.B1(n_845),
.B2(n_817),
.C(n_855),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_936),
.B(n_847),
.Y(n_942)
);

INVx1_ASAP7_75t_SL g943 ( 
.A(n_935),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_937),
.Y(n_944)
);

AOI221xp5_ASAP7_75t_L g945 ( 
.A1(n_934),
.A2(n_913),
.B1(n_905),
.B2(n_883),
.C(n_829),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_934),
.B(n_916),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_937),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_937),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_937),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_943),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_940),
.B(n_913),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_946),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_942),
.B(n_697),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_943),
.B(n_944),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_947),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_939),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_948),
.B(n_894),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_946),
.B(n_875),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_956),
.B(n_949),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_950),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_952),
.B(n_941),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_954),
.Y(n_962)
);

OAI221xp5_ASAP7_75t_L g963 ( 
.A1(n_953),
.A2(n_945),
.B1(n_707),
.B2(n_697),
.C(n_678),
.Y(n_963)
);

NAND2xp33_ASAP7_75t_SL g964 ( 
.A(n_958),
.B(n_877),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_957),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_955),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_951),
.B(n_894),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_960),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_959),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_962),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_966),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_965),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_961),
.B(n_958),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_967),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_964),
.B(n_886),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_963),
.A2(n_852),
.B1(n_689),
.B2(n_678),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_969),
.B(n_968),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_970),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_973),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_971),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_976),
.A2(n_710),
.B(n_836),
.C(n_835),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_972),
.B(n_880),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_974),
.B(n_877),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_975),
.B(n_889),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_973),
.B(n_710),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_969),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_979),
.B(n_983),
.Y(n_987)
);

AOI211xp5_ASAP7_75t_SL g988 ( 
.A1(n_986),
.A2(n_784),
.B(n_679),
.C(n_758),
.Y(n_988)
);

NAND4xp25_ASAP7_75t_L g989 ( 
.A(n_985),
.B(n_706),
.C(n_694),
.D(n_685),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_982),
.B(n_710),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_977),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_978),
.Y(n_992)
);

NOR2xp67_ASAP7_75t_L g993 ( 
.A(n_980),
.B(n_706),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_984),
.B(n_883),
.Y(n_994)
);

NOR3x1_ASAP7_75t_L g995 ( 
.A(n_981),
.B(n_679),
.C(n_760),
.Y(n_995)
);

NOR4xp25_ASAP7_75t_L g996 ( 
.A(n_992),
.B(n_874),
.C(n_885),
.D(n_887),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_993),
.B(n_883),
.Y(n_997)
);

NAND3xp33_ASAP7_75t_L g998 ( 
.A(n_987),
.B(n_680),
.C(n_685),
.Y(n_998)
);

AOI21xp33_ASAP7_75t_SL g999 ( 
.A1(n_991),
.A2(n_148),
.B(n_149),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_988),
.A2(n_694),
.B(n_835),
.C(n_828),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_990),
.A2(n_836),
.B(n_852),
.Y(n_1001)
);

OAI22xp33_ASAP7_75t_SL g1002 ( 
.A1(n_997),
.A2(n_994),
.B1(n_995),
.B2(n_989),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_998),
.A2(n_883),
.B1(n_874),
.B2(n_680),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_SL g1004 ( 
.A1(n_1001),
.A2(n_150),
.B(n_151),
.C(n_152),
.Y(n_1004)
);

AOI211xp5_ASAP7_75t_L g1005 ( 
.A1(n_999),
.A2(n_755),
.B(n_681),
.C(n_818),
.Y(n_1005)
);

AOI221xp5_ASAP7_75t_L g1006 ( 
.A1(n_1000),
.A2(n_887),
.B1(n_885),
.B2(n_822),
.C(n_821),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_996),
.Y(n_1007)
);

AO21x1_ASAP7_75t_L g1008 ( 
.A1(n_997),
.A2(n_691),
.B(n_827),
.Y(n_1008)
);

AOI221x1_ASAP7_75t_L g1009 ( 
.A1(n_999),
.A2(n_686),
.B1(n_821),
.B2(n_820),
.C(n_822),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_997),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_1000),
.A2(n_859),
.B(n_831),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_1002),
.B(n_896),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_1010),
.B(n_1007),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1003),
.A2(n_843),
.B1(n_892),
.B2(n_859),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1008),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1004),
.B(n_896),
.Y(n_1016)
);

AOI321xp33_ASAP7_75t_L g1017 ( 
.A1(n_1011),
.A2(n_818),
.A3(n_681),
.B1(n_824),
.B2(n_813),
.C(n_830),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1009),
.Y(n_1018)
);

AOI211xp5_ASAP7_75t_L g1019 ( 
.A1(n_1005),
.A2(n_681),
.B(n_797),
.C(n_869),
.Y(n_1019)
);

AOI222xp33_ASAP7_75t_L g1020 ( 
.A1(n_1006),
.A2(n_893),
.B1(n_879),
.B2(n_876),
.C1(n_819),
.C2(n_809),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_1013),
.A2(n_833),
.B(n_843),
.Y(n_1021)
);

NOR3xp33_ASAP7_75t_L g1022 ( 
.A(n_1012),
.B(n_830),
.C(n_824),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_1015),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1016),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_1018),
.A2(n_843),
.B1(n_893),
.B2(n_876),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1019),
.B(n_879),
.Y(n_1026)
);

NAND4xp25_ASAP7_75t_L g1027 ( 
.A(n_1017),
.B(n_830),
.C(n_813),
.D(n_814),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_1014),
.A2(n_859),
.B(n_831),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_1020),
.B(n_873),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_1013),
.A2(n_843),
.B(n_859),
.C(n_156),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1013),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1015),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1013),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_1031),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1023),
.Y(n_1035)
);

CKINVDCx16_ASAP7_75t_R g1036 ( 
.A(n_1033),
.Y(n_1036)
);

AOI221xp5_ASAP7_75t_L g1037 ( 
.A1(n_1032),
.A2(n_809),
.B1(n_814),
.B2(n_826),
.C(n_819),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_1024),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_1026),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_1022),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1025),
.A2(n_1029),
.B1(n_1027),
.B2(n_1028),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_1030),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1036),
.B(n_1021),
.Y(n_1043)
);

AOI22x1_ASAP7_75t_L g1044 ( 
.A1(n_1035),
.A2(n_153),
.B1(n_154),
.B2(n_157),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1038),
.Y(n_1045)
);

OAI22x1_ASAP7_75t_L g1046 ( 
.A1(n_1034),
.A2(n_826),
.B1(n_161),
.B2(n_162),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_SL g1047 ( 
.A1(n_1041),
.A2(n_1039),
.B(n_1040),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1042),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1037),
.B(n_873),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1045),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1048),
.B(n_873),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1043),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_1050),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_1053),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_1054),
.A2(n_1052),
.B1(n_1047),
.B2(n_1046),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1055),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1055),
.Y(n_1057)
);

OAI211xp5_ASAP7_75t_L g1058 ( 
.A1(n_1056),
.A2(n_1051),
.B(n_1044),
.C(n_1049),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1057),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_SL g1060 ( 
.A1(n_1059),
.A2(n_160),
.B1(n_164),
.B2(n_166),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1058),
.Y(n_1061)
);

OR2x6_ASAP7_75t_L g1062 ( 
.A(n_1061),
.B(n_167),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1060),
.A2(n_831),
.B1(n_170),
.B2(n_171),
.Y(n_1063)
);

NAND4xp25_ASAP7_75t_L g1064 ( 
.A(n_1063),
.B(n_168),
.C(n_172),
.D(n_174),
.Y(n_1064)
);

AOI211xp5_ASAP7_75t_L g1065 ( 
.A1(n_1064),
.A2(n_1062),
.B(n_177),
.C(n_178),
.Y(n_1065)
);


endmodule