module fake_netlist_5_1938_n_349 (n_91, n_82, n_10, n_24, n_86, n_83, n_61, n_90, n_75, n_65, n_78, n_74, n_57, n_96, n_37, n_31, n_13, n_66, n_60, n_16, n_43, n_0, n_58, n_9, n_69, n_18, n_42, n_22, n_1, n_45, n_46, n_21, n_94, n_38, n_80, n_4, n_35, n_73, n_17, n_92, n_19, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_62, n_71, n_85, n_95, n_59, n_26, n_55, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_36, n_76, n_87, n_27, n_64, n_77, n_81, n_28, n_89, n_70, n_68, n_93, n_72, n_32, n_41, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_349);

input n_91;
input n_82;
input n_10;
input n_24;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_65;
input n_78;
input n_74;
input n_57;
input n_96;
input n_37;
input n_31;
input n_13;
input n_66;
input n_60;
input n_16;
input n_43;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_42;
input n_22;
input n_1;
input n_45;
input n_46;
input n_21;
input n_94;
input n_38;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_62;
input n_71;
input n_85;
input n_95;
input n_59;
input n_26;
input n_55;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_81;
input n_28;
input n_89;
input n_70;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;

output n_349;

wire n_137;
wire n_294;
wire n_318;
wire n_194;
wire n_316;
wire n_248;
wire n_124;
wire n_146;
wire n_136;
wire n_315;
wire n_268;
wire n_127;
wire n_235;
wire n_226;
wire n_111;
wire n_155;
wire n_116;
wire n_284;
wire n_245;
wire n_139;
wire n_105;
wire n_280;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_244;
wire n_173;
wire n_198;
wire n_247;
wire n_314;
wire n_321;
wire n_292;
wire n_100;
wire n_212;
wire n_119;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_147;
wire n_307;
wire n_150;
wire n_106;
wire n_209;
wire n_259;
wire n_301;
wire n_186;
wire n_134;
wire n_191;
wire n_171;
wire n_153;
wire n_341;
wire n_204;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_122;
wire n_282;
wire n_331;
wire n_325;
wire n_132;
wire n_101;
wire n_281;
wire n_240;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_152;
wire n_317;
wire n_323;
wire n_195;
wire n_227;
wire n_271;
wire n_335;
wire n_123;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_267;
wire n_297;
wire n_156;
wire n_225;
wire n_219;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_158;
wire n_138;
wire n_264;
wire n_109;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_196;
wire n_211;
wire n_218;
wire n_181;
wire n_290;
wire n_221;
wire n_178;
wire n_287;
wire n_344;
wire n_104;
wire n_141;
wire n_336;
wire n_145;
wire n_337;
wire n_313;
wire n_216;
wire n_168;
wire n_164;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_296;
wire n_241;
wire n_184;
wire n_144;
wire n_114;
wire n_165;
wire n_213;
wire n_129;
wire n_342;
wire n_98;
wire n_197;
wire n_107;
wire n_236;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_277;
wire n_338;
wire n_149;
wire n_333;
wire n_309;
wire n_130;
wire n_322;
wire n_258;
wire n_151;
wire n_306;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_224;
wire n_228;
wire n_283;
wire n_112;
wire n_239;
wire n_310;
wire n_170;
wire n_332;
wire n_102;
wire n_161;
wire n_273;
wire n_270;
wire n_230;
wire n_118;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_312;
wire n_345;
wire n_210;
wire n_176;
wire n_182;
wire n_143;
wire n_237;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_229;
wire n_108;
wire n_177;
wire n_117;
wire n_326;
wire n_233;
wire n_205;
wire n_113;
wire n_246;
wire n_179;
wire n_125;
wire n_269;
wire n_128;
wire n_285;
wire n_120;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_193;
wire n_251;
wire n_160;
wire n_154;
wire n_148;
wire n_300;
wire n_159;
wire n_334;
wire n_175;
wire n_262;
wire n_238;
wire n_99;
wire n_319;
wire n_121;
wire n_242;
wire n_200;
wire n_162;
wire n_222;
wire n_115;
wire n_324;
wire n_199;
wire n_187;
wire n_103;
wire n_348;
wire n_166;
wire n_256;
wire n_305;
wire n_278;
wire n_110;

INVx1_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_11),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_66),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_54),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_1),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_14),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_21),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_8),
.Y(n_113)
);

INVxp67_ASAP7_75t_SL g114 ( 
.A(n_13),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_71),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_72),
.Y(n_120)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_90),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_56),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_0),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_31),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_5),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_69),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_46),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_27),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_4),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_0),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

NOR2xp67_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_1),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_2),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_105),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_131),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_2),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_112),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_3),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_138),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_103),
.B1(n_100),
.B2(n_130),
.Y(n_155)
);

OAI221xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_114),
.B1(n_115),
.B2(n_120),
.C(n_121),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

OR2x2_ASAP7_75t_SL g158 ( 
.A(n_147),
.B(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

AND2x4_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_114),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_106),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_101),
.Y(n_169)
);

AND2x4_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_120),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_102),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_121),
.Y(n_173)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_108),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_101),
.Y(n_176)
);

NAND2x1p5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_109),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_170),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_127),
.B1(n_133),
.B2(n_132),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_129),
.B(n_119),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_118),
.B(n_117),
.C(n_126),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_138),
.B(n_4),
.C(n_6),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_3),
.B(n_6),
.C(n_7),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_172),
.B(n_7),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_173),
.B(n_8),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_9),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_174),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_174),
.B(n_10),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_176),
.Y(n_196)
);

BUFx6f_ASAP7_75t_SL g197 ( 
.A(n_176),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_12),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_164),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_22),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_25),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_32),
.B(n_34),
.Y(n_208)
);

NOR2xp67_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_36),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_155),
.B(n_41),
.Y(n_212)
);

CKINVDCx6p67_ASAP7_75t_R g213 ( 
.A(n_197),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_42),
.B(n_43),
.Y(n_214)
);

AO21x2_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_44),
.B(n_45),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_178),
.A2(n_47),
.B(n_48),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_50),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_51),
.Y(n_218)
);

AO31x2_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_55),
.A3(n_57),
.B(n_58),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_59),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_204),
.Y(n_226)
);

AO21x2_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_61),
.B(n_62),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_63),
.B(n_64),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_181),
.A2(n_65),
.B(n_67),
.C(n_68),
.Y(n_230)
);

BUFx4f_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

AO31x2_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_70),
.A3(n_73),
.B(n_74),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

OAI21x1_ASAP7_75t_SL g234 ( 
.A1(n_180),
.A2(n_76),
.B(n_78),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g235 ( 
.A1(n_192),
.A2(n_79),
.B(n_80),
.Y(n_235)
);

OA21x2_ASAP7_75t_L g236 ( 
.A1(n_191),
.A2(n_81),
.B(n_82),
.Y(n_236)
);

OAI221xp5_ASAP7_75t_L g237 ( 
.A1(n_179),
.A2(n_182),
.B1(n_212),
.B2(n_188),
.C(n_186),
.Y(n_237)
);

AND2x4_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_199),
.Y(n_238)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_187),
.B(n_83),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_196),
.A2(n_197),
.B1(n_189),
.B2(n_200),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

NOR4xp25_ASAP7_75t_L g242 ( 
.A(n_184),
.B(n_86),
.C(n_89),
.D(n_91),
.Y(n_242)
);

AOI21x1_ASAP7_75t_L g243 ( 
.A1(n_201),
.A2(n_92),
.B(n_93),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_183),
.Y(n_244)
);

OAI21x1_ASAP7_75t_L g245 ( 
.A1(n_206),
.A2(n_94),
.B(n_95),
.Y(n_245)
);

BUFx2_ASAP7_75t_SL g246 ( 
.A(n_197),
.Y(n_246)
);

AO31x2_ASAP7_75t_L g247 ( 
.A1(n_208),
.A2(n_207),
.A3(n_211),
.B(n_206),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_SL g248 ( 
.A(n_217),
.B(n_223),
.Y(n_248)
);

CKINVDCx12_ASAP7_75t_R g249 ( 
.A(n_213),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_237),
.B1(n_233),
.B2(n_225),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

OR2x6_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_244),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_216),
.A2(n_227),
.B1(n_241),
.B2(n_238),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_231),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_218),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_240),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_R g265 ( 
.A(n_231),
.B(n_243),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_218),
.A2(n_230),
.B(n_236),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_221),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_R g269 ( 
.A(n_228),
.B(n_242),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_228),
.B(n_247),
.Y(n_270)
);

NOR3xp33_ASAP7_75t_SL g271 ( 
.A(n_229),
.B(n_242),
.C(n_219),
.Y(n_271)
);

AOI211xp5_ASAP7_75t_SL g272 ( 
.A1(n_219),
.A2(n_234),
.B(n_232),
.C(n_247),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_228),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_235),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_215),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_254),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_219),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_232),
.B(n_215),
.C(n_214),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_267),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_257),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_259),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_270),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_250),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_264),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_252),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_260),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_253),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_287),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_290),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_294),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

NAND2x1p5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_286),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

AND3x1_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_271),
.C(n_288),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

AO21x2_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_281),
.B(n_269),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_289),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_278),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_293),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_314),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_315),
.Y(n_320)
);

A2O1A1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_311),
.A2(n_248),
.B(n_271),
.C(n_272),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

NOR3xp33_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_291),
.C(n_300),
.Y(n_323)
);

AOI221xp5_ASAP7_75t_L g324 ( 
.A1(n_304),
.A2(n_292),
.B1(n_266),
.B2(n_269),
.C(n_281),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_304),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_302),
.A2(n_265),
.B1(n_252),
.B2(n_288),
.Y(n_326)
);

NOR3xp33_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_279),
.C(n_268),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_252),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_312),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_308),
.A2(n_249),
.B1(n_275),
.B2(n_274),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_319),
.B(n_309),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_309),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_310),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_309),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_316),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_322),
.Y(n_336)
);

NAND2x1_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_329),
.Y(n_337)
);

OAI211xp5_ASAP7_75t_SL g338 ( 
.A1(n_331),
.A2(n_326),
.B(n_330),
.C(n_323),
.Y(n_338)
);

NOR3xp33_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_334),
.C(n_321),
.Y(n_339)
);

A2O1A1Ixp33_ASAP7_75t_L g340 ( 
.A1(n_337),
.A2(n_324),
.B(n_317),
.C(n_333),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_339),
.Y(n_342)
);

NAND4xp25_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_324),
.C(n_332),
.D(n_327),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_341),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_344),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_343),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_345),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_346),
.B1(n_318),
.B2(n_310),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_348),
.A2(n_318),
.B1(n_310),
.B2(n_335),
.Y(n_349)
);


endmodule