module fake_ariane_243_n_1995 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1995);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1995;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_925;
wire n_246;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_77),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_36),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_17),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_131),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_13),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_116),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_187),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_11),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_14),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_90),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_174),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_7),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_97),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_40),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_84),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_78),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_2),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_107),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_0),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_132),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_41),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_65),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_47),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_94),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_85),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_81),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_11),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_69),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_57),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_126),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_111),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_13),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_143),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_44),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_102),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_38),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_152),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_34),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_46),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_62),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_144),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_42),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_83),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_67),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_1),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_109),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_24),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_36),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_135),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_50),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_91),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_21),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_69),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_67),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_44),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_57),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_142),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_34),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_189),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_60),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_68),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_74),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_153),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_66),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_114),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_177),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_117),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_25),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_93),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_79),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_65),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_26),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_168),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_156),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_32),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_73),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_18),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_60),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_146),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_161),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_48),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_26),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_75),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_38),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_186),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_101),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_62),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_42),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_80),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_139),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_166),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_47),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_119),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_179),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_88),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_130),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_3),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_188),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_72),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_59),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_183),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_105),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_92),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_127),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_165),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_54),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_182),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_76),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_155),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_82),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_157),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_129),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_21),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_173),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_104),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_70),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_6),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_2),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_0),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_52),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_25),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_7),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_16),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_54),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_33),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_61),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_9),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_178),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_68),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_86),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_5),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_120),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_18),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_20),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_46),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_134),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_106),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_171),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_28),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_49),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_115),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_8),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_23),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_140),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_108),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_103),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_51),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_71),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_43),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_110),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_66),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_113),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_145),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_95),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_87),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_19),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_43),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_64),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_61),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_159),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_35),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_180),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_89),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_48),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_160),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_141),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_24),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_128),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_10),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_31),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_55),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_122),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_19),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_118),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_32),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_28),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_175),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_151),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_37),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_154),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_49),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_52),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_198),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_215),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_212),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_339),
.B(n_1),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_212),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_212),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_323),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_308),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_323),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_286),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_309),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_274),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_286),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_274),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_339),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_204),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_352),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_352),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_201),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_352),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_328),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_352),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_230),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_204),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_201),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_330),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_216),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_R g409 ( 
.A(n_360),
.B(n_137),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_315),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_230),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_311),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_315),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_250),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_208),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_208),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_311),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_236),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_236),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_192),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_241),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_332),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_241),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_266),
.Y(n_424)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_238),
.B(n_345),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_266),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_341),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_275),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_290),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_275),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_351),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_290),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_276),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_276),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_290),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_238),
.B(n_3),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_351),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_194),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_282),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_205),
.B(n_4),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_340),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_196),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_199),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_340),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_282),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_295),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_295),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_298),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_290),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_340),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_205),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_298),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_316),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_214),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_340),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_223),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_224),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_200),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_200),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_225),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_316),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_200),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_228),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_217),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_318),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_217),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_217),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_318),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_207),
.B(n_4),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_232),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_234),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_324),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_324),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_207),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_209),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_429),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_471),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_400),
.B(n_406),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_400),
.B(n_290),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_429),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_432),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_432),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_406),
.B(n_345),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_451),
.B(n_331),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_435),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_435),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_383),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_385),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_386),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_404),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_387),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_451),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_474),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_388),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_474),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_475),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_398),
.B(n_211),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_475),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_390),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_449),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_L g501 ( 
.A(n_384),
.B(n_219),
.Y(n_501)
);

CKINVDCx11_ASAP7_75t_R g502 ( 
.A(n_414),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_415),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_419),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_391),
.B(n_306),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_421),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_423),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_396),
.B(n_350),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_404),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_394),
.B(n_331),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_424),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_426),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_428),
.Y(n_513)
);

AND2x6_ASAP7_75t_L g514 ( 
.A(n_440),
.B(n_193),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_410),
.B(n_333),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_434),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_431),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_439),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_413),
.B(n_333),
.Y(n_520)
);

OA21x2_ASAP7_75t_L g521 ( 
.A1(n_446),
.A2(n_221),
.B(n_209),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_452),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_453),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_461),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_465),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_381),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_468),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_411),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_473),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_469),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_398),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_425),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_436),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_416),
.B(n_221),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_418),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_430),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_411),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_445),
.B(n_337),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_447),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_SL g540 ( 
.A(n_396),
.B(n_235),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_448),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_412),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_472),
.B(n_337),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_L g544 ( 
.A(n_399),
.B(n_219),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_437),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_412),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_399),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_401),
.B(n_211),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_405),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_401),
.B(n_226),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_403),
.B(n_267),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_405),
.B(n_354),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_403),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_408),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_547),
.B(n_393),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_542),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_531),
.B(n_226),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_492),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_492),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_500),
.B(n_393),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_492),
.Y(n_561)
);

INVxp67_ASAP7_75t_SL g562 ( 
.A(n_492),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_547),
.B(n_395),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_492),
.Y(n_564)
);

BUFx10_ASAP7_75t_L g565 ( 
.A(n_531),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_500),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_492),
.Y(n_567)
);

OAI22xp33_ASAP7_75t_L g568 ( 
.A1(n_550),
.A2(n_395),
.B1(n_417),
.B2(n_441),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_492),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_492),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_492),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_493),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_493),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_547),
.B(n_420),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_531),
.B(n_227),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_536),
.Y(n_576)
);

INVx6_ASAP7_75t_L g577 ( 
.A(n_484),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_547),
.B(n_420),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_486),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_486),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_478),
.B(n_438),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_531),
.B(n_227),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_493),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_553),
.B(n_438),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_476),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_500),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_486),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_495),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_478),
.B(n_442),
.Y(n_589)
);

BUFx4f_ASAP7_75t_L g590 ( 
.A(n_531),
.Y(n_590)
);

INVxp33_ASAP7_75t_L g591 ( 
.A(n_477),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_495),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_530),
.A2(n_397),
.B1(n_409),
.B2(n_417),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_478),
.B(n_442),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_478),
.B(n_536),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_486),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_495),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_481),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_494),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_494),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_484),
.B(n_354),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_553),
.B(n_443),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_542),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_542),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_481),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_530),
.A2(n_362),
.B1(n_369),
.B2(n_356),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_496),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_481),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_484),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_482),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_531),
.B(n_231),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_482),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_482),
.Y(n_613)
);

INVx8_ASAP7_75t_L g614 ( 
.A(n_514),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_549),
.B(n_443),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_536),
.B(n_356),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_553),
.B(n_454),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_485),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g619 ( 
.A1(n_550),
.A2(n_456),
.B1(n_457),
.B2(n_454),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_497),
.B(n_456),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_549),
.B(n_457),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_553),
.B(n_460),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_485),
.Y(n_623)
);

AND2x2_ASAP7_75t_SL g624 ( 
.A(n_544),
.B(n_521),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_500),
.B(n_460),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_530),
.A2(n_369),
.B1(n_362),
.B2(n_444),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_496),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_530),
.B(n_463),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_484),
.B(n_242),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_494),
.Y(n_630)
);

INVxp33_ASAP7_75t_L g631 ( 
.A(n_477),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_514),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_494),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_494),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_553),
.B(n_463),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_508),
.A2(n_349),
.B1(n_218),
.B2(n_244),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_496),
.Y(n_637)
);

BUFx4f_ASAP7_75t_L g638 ( 
.A(n_531),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_536),
.B(n_470),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_498),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_502),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_485),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_498),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_497),
.B(n_470),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_498),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_503),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_553),
.B(n_240),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_508),
.A2(n_321),
.B1(n_245),
.B2(n_247),
.Y(n_648)
);

AND3x2_ASAP7_75t_L g649 ( 
.A(n_546),
.B(n_312),
.C(n_249),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_533),
.B(n_260),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_484),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_548),
.B(n_450),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_494),
.Y(n_653)
);

INVx4_ASAP7_75t_SL g654 ( 
.A(n_514),
.Y(n_654)
);

INVx5_ASAP7_75t_L g655 ( 
.A(n_514),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_539),
.B(n_455),
.Y(n_656)
);

BUFx4f_ASAP7_75t_L g657 ( 
.A(n_531),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_476),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_476),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_476),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_484),
.B(n_242),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_546),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_531),
.B(n_535),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_517),
.Y(n_664)
);

CKINVDCx11_ASAP7_75t_R g665 ( 
.A(n_502),
.Y(n_665)
);

INVx6_ASAP7_75t_L g666 ( 
.A(n_479),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_533),
.B(n_261),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_476),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_539),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_517),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_514),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_476),
.Y(n_672)
);

OR2x6_ASAP7_75t_L g673 ( 
.A(n_483),
.B(n_334),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_R g674 ( 
.A(n_546),
.B(n_382),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_517),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_518),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_517),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_476),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_514),
.A2(n_375),
.B1(n_336),
.B2(n_334),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_526),
.Y(n_680)
);

OAI21xp33_ASAP7_75t_L g681 ( 
.A1(n_534),
.A2(n_249),
.B(n_231),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_539),
.B(n_251),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_476),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_539),
.B(n_252),
.Y(n_684)
);

NOR3xp33_ASAP7_75t_L g685 ( 
.A(n_540),
.B(n_254),
.C(n_253),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_517),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_533),
.B(n_281),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_535),
.B(n_281),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_535),
.B(n_256),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_541),
.B(n_284),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_476),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_548),
.B(n_458),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_517),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_527),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_541),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_541),
.B(n_284),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_527),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_549),
.B(n_258),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_551),
.B(n_459),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_551),
.B(n_554),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_527),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_527),
.B(n_296),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_527),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_480),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_480),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_527),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_554),
.B(n_259),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_566),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_676),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_676),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_574),
.B(n_554),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_628),
.B(n_555),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_566),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_680),
.Y(n_714)
);

NOR3xp33_ASAP7_75t_L g715 ( 
.A(n_556),
.B(n_540),
.C(n_509),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_601),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_620),
.A2(n_544),
.B1(n_514),
.B2(n_509),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_586),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_695),
.B(n_538),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_572),
.Y(n_720)
);

BUFx5_ASAP7_75t_L g721 ( 
.A(n_565),
.Y(n_721)
);

AND2x6_ASAP7_75t_SL g722 ( 
.A(n_665),
.B(n_552),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_586),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_590),
.B(n_490),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_695),
.B(n_538),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_556),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_603),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_644),
.A2(n_514),
.B1(n_528),
.B2(n_490),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_572),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_579),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_573),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_590),
.B(n_528),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_579),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_603),
.B(n_537),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_625),
.B(n_537),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_635),
.B(n_578),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_604),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_580),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_590),
.B(n_552),
.Y(n_739)
);

NOR2x1p5_ASAP7_75t_L g740 ( 
.A(n_641),
.B(n_552),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_L g741 ( 
.A1(n_636),
.A2(n_534),
.B1(n_504),
.B2(n_506),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_604),
.Y(n_742)
);

BUFx10_ASAP7_75t_L g743 ( 
.A(n_641),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_573),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_576),
.B(n_538),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_576),
.B(n_538),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_583),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_580),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_669),
.B(n_543),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_L g750 ( 
.A(n_557),
.B(n_514),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_638),
.B(n_657),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_560),
.B(n_563),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_669),
.B(n_543),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_584),
.B(n_505),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_602),
.B(n_505),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_638),
.B(n_552),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_583),
.Y(n_757)
);

BUFx6f_ASAP7_75t_SL g758 ( 
.A(n_616),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_577),
.A2(n_504),
.B1(n_506),
.B2(n_503),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_588),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_587),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_601),
.B(n_552),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_588),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_617),
.B(n_552),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_638),
.B(n_479),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_592),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_622),
.B(n_543),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_614),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_662),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_592),
.A2(n_504),
.B(n_506),
.C(n_503),
.Y(n_770)
);

BUFx5_ASAP7_75t_L g771 ( 
.A(n_565),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_639),
.B(n_543),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_L g773 ( 
.A(n_557),
.B(n_514),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_681),
.A2(n_511),
.B(n_512),
.C(n_507),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_577),
.A2(n_511),
.B1(n_512),
.B2(n_507),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_L g776 ( 
.A1(n_636),
.A2(n_511),
.B1(n_512),
.B2(n_507),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_639),
.B(n_513),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_609),
.B(n_513),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_681),
.A2(n_514),
.B1(n_521),
.B2(n_483),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_595),
.B(n_513),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_587),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_595),
.B(n_519),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_682),
.B(n_519),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_609),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_682),
.B(n_519),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_597),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_684),
.B(n_522),
.Y(n_787)
);

INVx8_ASAP7_75t_L g788 ( 
.A(n_614),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_609),
.B(n_522),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_662),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_614),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_L g792 ( 
.A(n_557),
.B(n_514),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_596),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_651),
.B(n_522),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_684),
.B(n_523),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_646),
.B(n_523),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_651),
.B(n_523),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_674),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_646),
.B(n_524),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_581),
.B(n_524),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_581),
.B(n_524),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_589),
.B(n_529),
.Y(n_802)
);

BUFx6f_ASAP7_75t_SL g803 ( 
.A(n_616),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_657),
.B(n_479),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_597),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_651),
.B(n_529),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_SL g807 ( 
.A(n_689),
.B(n_529),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_589),
.B(n_545),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_596),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_594),
.B(n_483),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_619),
.B(n_515),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_594),
.B(n_483),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_601),
.B(n_545),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_650),
.B(n_483),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_577),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_667),
.B(n_483),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_577),
.A2(n_279),
.B1(n_262),
.B2(n_269),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_700),
.B(n_515),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_689),
.B(n_479),
.Y(n_819)
);

AND2x4_ASAP7_75t_SL g820 ( 
.A(n_656),
.B(n_389),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_679),
.A2(n_521),
.B1(n_515),
.B2(n_525),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_607),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_656),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_616),
.B(n_479),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_601),
.B(n_545),
.Y(n_825)
);

NAND3x1_ASAP7_75t_L g826 ( 
.A(n_648),
.B(n_427),
.C(n_422),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_657),
.B(n_479),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_607),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_627),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_627),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_637),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_637),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_601),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_666),
.B(n_515),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_624),
.B(n_525),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_616),
.B(n_525),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_675),
.B(n_525),
.Y(n_837)
);

AND2x4_ASAP7_75t_SL g838 ( 
.A(n_629),
.B(n_392),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_675),
.B(n_487),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_629),
.A2(n_273),
.B1(n_270),
.B2(n_280),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_615),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_615),
.B(n_518),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_640),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_624),
.B(n_487),
.Y(n_844)
);

OAI22xp33_ASAP7_75t_L g845 ( 
.A1(n_648),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.Y(n_845)
);

INVxp33_ASAP7_75t_L g846 ( 
.A(n_591),
.Y(n_846)
);

BUFx8_ASAP7_75t_L g847 ( 
.A(n_621),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_640),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_666),
.B(n_487),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_643),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_624),
.B(n_565),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_621),
.B(n_545),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_643),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_645),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_645),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_629),
.A2(n_320),
.B1(n_304),
.B2(n_327),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_675),
.B(n_697),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_666),
.B(n_488),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_SL g859 ( 
.A(n_652),
.B(n_518),
.Y(n_859)
);

NAND2xp33_ASAP7_75t_L g860 ( 
.A(n_557),
.B(n_488),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_697),
.B(n_488),
.Y(n_861)
);

AOI221xp5_ASAP7_75t_L g862 ( 
.A1(n_626),
.A2(n_510),
.B1(n_516),
.B2(n_520),
.C(n_285),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_697),
.B(n_489),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_598),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_666),
.B(n_489),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_614),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_664),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_629),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_598),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_664),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_701),
.B(n_489),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_L g872 ( 
.A(n_568),
.B(n_477),
.C(n_526),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_670),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_565),
.B(n_491),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_614),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_707),
.B(n_701),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_701),
.B(n_491),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_629),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_661),
.A2(n_501),
.B1(n_521),
.B2(n_520),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_712),
.A2(n_692),
.B1(n_699),
.B2(n_593),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_712),
.A2(n_661),
.B1(n_673),
.B2(n_647),
.Y(n_881)
);

O2A1O1Ixp5_ASAP7_75t_L g882 ( 
.A1(n_751),
.A2(n_663),
.B(n_690),
.C(n_688),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_822),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_730),
.Y(n_884)
);

OAI21x1_ASAP7_75t_SL g885 ( 
.A1(n_770),
.A2(n_632),
.B(n_671),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_735),
.B(n_698),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_741),
.A2(n_661),
.B1(n_673),
.B2(n_685),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_751),
.A2(n_562),
.B(n_670),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_733),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_857),
.A2(n_686),
.B(n_677),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_735),
.B(n_698),
.Y(n_891)
);

AND2x2_ASAP7_75t_SL g892 ( 
.A(n_762),
.B(n_521),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_711),
.B(n_706),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_762),
.B(n_654),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_772),
.B(n_696),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_734),
.B(n_631),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_738),
.Y(n_897)
);

O2A1O1Ixp5_ASAP7_75t_L g898 ( 
.A1(n_811),
.A2(n_702),
.B(n_677),
.C(n_693),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_772),
.A2(n_706),
.B(n_606),
.C(n_693),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_768),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_719),
.B(n_687),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_742),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_841),
.B(n_706),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_725),
.B(n_754),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_752),
.B(n_599),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_874),
.A2(n_694),
.B(n_686),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_811),
.A2(n_703),
.B(n_694),
.C(n_600),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_874),
.A2(n_703),
.B(n_661),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_754),
.B(n_599),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_741),
.A2(n_661),
.B1(n_673),
.B2(n_402),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_764),
.A2(n_600),
.B(n_630),
.C(n_599),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_755),
.B(n_600),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_835),
.A2(n_633),
.B(n_630),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_721),
.B(n_632),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_784),
.A2(n_630),
.B1(n_634),
.B2(n_633),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_752),
.B(n_633),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_SL g917 ( 
.A(n_714),
.B(n_407),
.Y(n_917)
);

OAI321xp33_ASAP7_75t_L g918 ( 
.A1(n_776),
.A2(n_673),
.A3(n_532),
.B1(n_353),
.B2(n_296),
.C(n_297),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_839),
.A2(n_653),
.B(n_634),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_828),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_861),
.A2(n_871),
.B(n_863),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_755),
.B(n_634),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_764),
.A2(n_653),
.B(n_499),
.C(n_491),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_829),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_709),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_721),
.B(n_632),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_L g927 ( 
.A(n_769),
.B(n_317),
.C(n_314),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_837),
.A2(n_653),
.B(n_567),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_777),
.B(n_800),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_L g930 ( 
.A1(n_767),
.A2(n_322),
.B(n_319),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_768),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_721),
.B(n_632),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_736),
.B(n_673),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_776),
.A2(n_521),
.B1(n_608),
.B2(n_610),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_801),
.B(n_649),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_802),
.B(n_605),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_721),
.B(n_671),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_767),
.B(n_605),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_852),
.B(n_745),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_746),
.B(n_608),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_765),
.A2(n_827),
.B(n_804),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_835),
.A2(n_567),
.B(n_561),
.Y(n_942)
);

NAND3xp33_ASAP7_75t_L g943 ( 
.A(n_726),
.B(n_501),
.C(n_671),
.Y(n_943)
);

O2A1O1Ixp5_ASAP7_75t_L g944 ( 
.A1(n_724),
.A2(n_569),
.B(n_559),
.C(n_564),
.Y(n_944)
);

NAND2x1_ASAP7_75t_L g945 ( 
.A(n_866),
.B(n_569),
.Y(n_945)
);

BUFx4f_ASAP7_75t_L g946 ( 
.A(n_727),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_710),
.B(n_510),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_749),
.B(n_610),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_765),
.A2(n_571),
.B(n_561),
.Y(n_949)
);

AOI21xp33_ASAP7_75t_L g950 ( 
.A1(n_842),
.A2(n_613),
.B(n_612),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_748),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_804),
.A2(n_571),
.B(n_559),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_753),
.B(n_612),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_827),
.A2(n_564),
.B(n_558),
.Y(n_954)
);

AO21x1_ASAP7_75t_L g955 ( 
.A1(n_844),
.A2(n_299),
.B(n_297),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_844),
.A2(n_558),
.B(n_569),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_737),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_790),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_761),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_783),
.B(n_613),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_785),
.B(n_618),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_787),
.B(n_618),
.Y(n_962)
);

NAND2x1p5_ASAP7_75t_L g963 ( 
.A(n_815),
.B(n_655),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_795),
.B(n_623),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_877),
.A2(n_575),
.B(n_557),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_810),
.A2(n_499),
.B(n_491),
.C(n_623),
.Y(n_966)
);

AOI21x1_ASAP7_75t_L g967 ( 
.A1(n_739),
.A2(n_659),
.B(n_658),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_815),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_851),
.A2(n_659),
.B(n_658),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_808),
.B(n_510),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_819),
.B(n_642),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_851),
.A2(n_672),
.B(n_660),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_778),
.A2(n_570),
.B1(n_655),
.B2(n_347),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_812),
.A2(n_499),
.B(n_642),
.C(n_516),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_736),
.A2(n_672),
.B(n_660),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_721),
.B(n_570),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_877),
.A2(n_704),
.B(n_691),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_778),
.B(n_789),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_739),
.A2(n_704),
.B(n_691),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_789),
.B(n_557),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_823),
.B(n_705),
.Y(n_981)
);

AO21x1_ASAP7_75t_L g982 ( 
.A1(n_807),
.A2(n_302),
.B(n_299),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_813),
.B(n_654),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_794),
.A2(n_575),
.B(n_557),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_813),
.B(n_654),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_794),
.A2(n_582),
.B(n_575),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_721),
.B(n_570),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_797),
.B(n_575),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_797),
.B(n_575),
.Y(n_989)
);

AOI21xp33_ASAP7_75t_L g990 ( 
.A1(n_859),
.A2(n_464),
.B(n_462),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_756),
.A2(n_705),
.B(n_570),
.Y(n_991)
);

OAI321xp33_ASAP7_75t_L g992 ( 
.A1(n_717),
.A2(n_532),
.A3(n_358),
.B1(n_353),
.B2(n_326),
.C(n_302),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_806),
.A2(n_570),
.B1(n_655),
.B2(n_374),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_830),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_820),
.B(n_510),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_781),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_850),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_825),
.B(n_499),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_806),
.B(n_575),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_756),
.A2(n_668),
.B(n_585),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_825),
.B(n_466),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_728),
.A2(n_575),
.B1(n_582),
.B2(n_611),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_793),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_771),
.B(n_655),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_780),
.A2(n_520),
.B(n_516),
.C(n_326),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_782),
.A2(n_520),
.B(n_516),
.C(n_358),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_862),
.A2(n_521),
.B1(n_582),
.B2(n_611),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_796),
.A2(n_668),
.B(n_585),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_809),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_814),
.B(n_582),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_716),
.B(n_833),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_838),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_853),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_743),
.Y(n_1014)
);

AOI21x1_ASAP7_75t_L g1015 ( 
.A1(n_720),
.A2(n_278),
.B(n_267),
.Y(n_1015)
);

INVx3_ASAP7_75t_SL g1016 ( 
.A(n_743),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_799),
.A2(n_732),
.B(n_724),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_732),
.A2(n_668),
.B(n_585),
.Y(n_1018)
);

AOI21x1_ASAP7_75t_L g1019 ( 
.A1(n_729),
.A2(n_344),
.B(n_278),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_867),
.A2(n_668),
.B(n_585),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_864),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_870),
.A2(n_668),
.B(n_585),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_869),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_779),
.A2(n_611),
.B1(n_582),
.B2(n_532),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_716),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_873),
.A2(n_683),
.B(n_678),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_759),
.A2(n_376),
.B(n_378),
.C(n_344),
.Y(n_1027)
);

OAI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_833),
.A2(n_325),
.B1(n_359),
.B2(n_357),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_731),
.A2(n_831),
.B(n_757),
.C(n_843),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_758),
.Y(n_1030)
);

INVx5_ASAP7_75t_L g1031 ( 
.A(n_788),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_816),
.B(n_582),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_768),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_744),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_846),
.B(n_467),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_834),
.B(n_582),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_876),
.B(n_655),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_847),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_834),
.B(n_611),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_768),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_798),
.B(n_329),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_849),
.B(n_858),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_876),
.B(n_655),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_849),
.B(n_858),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_758),
.B(n_683),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_775),
.A2(n_376),
.B(n_378),
.C(n_355),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_708),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_747),
.A2(n_683),
.B(n_678),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_826),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_865),
.B(n_611),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_840),
.A2(n_338),
.B(n_346),
.C(n_365),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_771),
.B(n_791),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_865),
.B(n_611),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_713),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_803),
.B(n_683),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_771),
.B(n_683),
.Y(n_1056)
);

AOI33xp33_ASAP7_75t_L g1057 ( 
.A1(n_760),
.A2(n_367),
.A3(n_368),
.B1(n_371),
.B2(n_373),
.B3(n_377),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_818),
.A2(n_611),
.B(n_654),
.Y(n_1058)
);

NOR2x1_ASAP7_75t_L g1059 ( 
.A(n_740),
.B(n_678),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_763),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_766),
.A2(n_678),
.B(n_191),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_715),
.B(n_379),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_718),
.Y(n_1063)
);

AOI21xp33_ASAP7_75t_L g1064 ( 
.A1(n_856),
.A2(n_380),
.B(n_678),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_824),
.B(n_195),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_818),
.A2(n_277),
.B(n_372),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_847),
.Y(n_1067)
);

OAI321xp33_ASAP7_75t_L g1068 ( 
.A1(n_779),
.A2(n_480),
.A3(n_364),
.B1(n_343),
.B2(n_291),
.C(n_243),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_868),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_786),
.B(n_197),
.Y(n_1070)
);

NOR2x1_ASAP7_75t_R g1071 ( 
.A(n_722),
.B(n_202),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_805),
.A2(n_848),
.B(n_832),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_854),
.A2(n_283),
.B(n_370),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_894),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_883),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_SL g1076 ( 
.A(n_1014),
.B(n_817),
.C(n_855),
.Y(n_1076)
);

AO32x1_ASAP7_75t_L g1077 ( 
.A1(n_920),
.A2(n_723),
.A3(n_845),
.B1(n_774),
.B2(n_879),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_978),
.A2(n_886),
.B1(n_891),
.B2(n_880),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_924),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_886),
.A2(n_872),
.B(n_774),
.C(n_878),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_946),
.B(n_868),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_891),
.A2(n_878),
.B(n_845),
.C(n_836),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_933),
.A2(n_792),
.B(n_773),
.C(n_750),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_933),
.A2(n_860),
.B(n_821),
.C(n_788),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_904),
.B(n_821),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_929),
.A2(n_788),
.B(n_866),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1013),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_910),
.A2(n_803),
.B1(n_875),
.B2(n_791),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_970),
.B(n_791),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_896),
.B(n_791),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_1016),
.Y(n_1091)
);

AND3x1_ASAP7_75t_SL g1092 ( 
.A(n_1034),
.B(n_5),
.C(n_6),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1042),
.A2(n_771),
.B(n_875),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1044),
.A2(n_771),
.B(n_875),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_894),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_994),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_895),
.B(n_875),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_902),
.Y(n_1098)
);

OAI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_887),
.A2(n_917),
.B1(n_881),
.B2(n_946),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_995),
.B(n_8),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_958),
.Y(n_1101)
);

BUFx4f_ASAP7_75t_L g1102 ( 
.A(n_1016),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_939),
.B(n_947),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_1051),
.A2(n_9),
.B(n_10),
.C(n_12),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_1038),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_930),
.A2(n_12),
.B(n_14),
.C(n_15),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_1025),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_1031),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_1067),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_1025),
.Y(n_1110)
);

INVxp67_ASAP7_75t_L g1111 ( 
.A(n_1001),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_889),
.Y(n_1112)
);

AO32x2_ASAP7_75t_L g1113 ( 
.A1(n_915),
.A2(n_480),
.A3(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_1113)
);

INVx5_ASAP7_75t_L g1114 ( 
.A(n_983),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_901),
.A2(n_15),
.B(n_22),
.C(n_23),
.Y(n_1115)
);

AND2x6_ASAP7_75t_SL g1116 ( 
.A(n_1001),
.B(n_22),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_1035),
.Y(n_1117)
);

BUFx8_ASAP7_75t_L g1118 ( 
.A(n_1012),
.Y(n_1118)
);

XOR2xp5_ASAP7_75t_L g1119 ( 
.A(n_1030),
.B(n_203),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_905),
.B(n_771),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_921),
.A2(n_206),
.B(n_366),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_957),
.B(n_210),
.Y(n_1122)
);

OR2x6_ASAP7_75t_L g1123 ( 
.A(n_983),
.B(n_480),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_905),
.A2(n_287),
.B1(n_213),
.B2(n_363),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_1069),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_934),
.A2(n_288),
.B1(n_220),
.B2(n_361),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_1011),
.B(n_222),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_916),
.B(n_1011),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1030),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_916),
.B(n_903),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_990),
.B(n_229),
.Y(n_1131)
);

OAI22x1_ASAP7_75t_L g1132 ( 
.A1(n_1049),
.A2(n_1062),
.B1(n_935),
.B2(n_925),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_893),
.A2(n_293),
.B1(n_233),
.B2(n_348),
.Y(n_1133)
);

BUFx8_ASAP7_75t_L g1134 ( 
.A(n_1041),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_1028),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_893),
.A2(n_289),
.B(n_237),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_903),
.B(n_27),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1060),
.B(n_29),
.Y(n_1138)
);

NAND2x1p5_ASAP7_75t_L g1139 ( 
.A(n_985),
.B(n_480),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1028),
.A2(n_1046),
.B(n_1029),
.C(n_911),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_892),
.A2(n_294),
.B1(n_255),
.B2(n_239),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_960),
.A2(n_292),
.B(n_246),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_985),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_1031),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_SL g1145 ( 
.A(n_892),
.B(n_248),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_909),
.A2(n_300),
.B1(n_257),
.B2(n_263),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_961),
.A2(n_303),
.B(n_264),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1059),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_962),
.A2(n_305),
.B(n_265),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1031),
.B(n_301),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_997),
.B(n_912),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1031),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_964),
.A2(n_307),
.B(n_268),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_SL g1154 ( 
.A1(n_1005),
.A2(n_30),
.B(n_31),
.C(n_33),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_968),
.Y(n_1155)
);

BUFx8_ASAP7_75t_L g1156 ( 
.A(n_1071),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_941),
.A2(n_480),
.B(n_310),
.C(n_271),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_968),
.B(n_922),
.Y(n_1158)
);

NAND2x1p5_ASAP7_75t_L g1159 ( 
.A(n_1033),
.B(n_480),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_889),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1056),
.A2(n_313),
.B(n_272),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_951),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_951),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1056),
.A2(n_335),
.B(n_342),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_998),
.B(n_35),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1029),
.A2(n_37),
.B(n_39),
.C(n_40),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_918),
.B(n_39),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1047),
.B(n_41),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1021),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1023),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_934),
.A2(n_480),
.B1(n_364),
.B2(n_343),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_998),
.B(n_45),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_980),
.A2(n_364),
.B(n_343),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_938),
.B(n_45),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_988),
.A2(n_364),
.B(n_343),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_911),
.A2(n_50),
.B(n_51),
.C(n_53),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_900),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_989),
.A2(n_364),
.B(n_343),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_884),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_936),
.B(n_1072),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_999),
.A2(n_291),
.B(n_243),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_897),
.Y(n_1182)
);

AOI33xp33_ASAP7_75t_L g1183 ( 
.A1(n_1006),
.A2(n_53),
.A3(n_55),
.B1(n_56),
.B2(n_58),
.B3(n_59),
.Y(n_1183)
);

AOI21xp33_ASAP7_75t_L g1184 ( 
.A1(n_1066),
.A2(n_992),
.B(n_974),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1009),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1007),
.A2(n_291),
.B1(n_243),
.B2(n_193),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_927),
.B(n_56),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_976),
.A2(n_291),
.B(n_243),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_900),
.Y(n_1189)
);

NAND2x1p5_ASAP7_75t_L g1190 ( 
.A(n_1033),
.B(n_243),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1057),
.B(n_58),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1009),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1045),
.B(n_63),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1054),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1045),
.Y(n_1195)
);

NOR3xp33_ASAP7_75t_SL g1196 ( 
.A(n_1073),
.B(n_63),
.C(n_64),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_959),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_996),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1063),
.A2(n_193),
.B1(n_219),
.B2(n_70),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_900),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1055),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1003),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_981),
.Y(n_1203)
);

AND2x6_ASAP7_75t_L g1204 ( 
.A(n_931),
.B(n_193),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_1055),
.B(n_193),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_976),
.A2(n_138),
.B(n_96),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_931),
.B(n_219),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_942),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_981),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_940),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_SL g1211 ( 
.A(n_984),
.B(n_219),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1068),
.A2(n_219),
.B(n_71),
.C(n_99),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_987),
.A2(n_98),
.B(n_100),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1015),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_948),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_907),
.A2(n_219),
.B(n_121),
.C(n_124),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1019),
.Y(n_1217)
);

OAI21xp33_ASAP7_75t_SL g1218 ( 
.A1(n_986),
.A2(n_219),
.B(n_125),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_SL g1219 ( 
.A1(n_913),
.A2(n_219),
.B(n_133),
.C(n_136),
.Y(n_1219)
);

BUFx2_ASAP7_75t_SL g1220 ( 
.A(n_931),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1040),
.B(n_112),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1017),
.A2(n_899),
.B(n_908),
.C(n_1007),
.Y(n_1222)
);

INVxp67_ASAP7_75t_L g1223 ( 
.A(n_1070),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_953),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_987),
.A2(n_147),
.B(n_148),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_SL g1226 ( 
.A1(n_1024),
.A2(n_149),
.B1(n_150),
.B2(n_158),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1040),
.B(n_170),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_914),
.A2(n_172),
.B(n_176),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_899),
.A2(n_181),
.B1(n_184),
.B2(n_1024),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_982),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_950),
.A2(n_1065),
.B1(n_1064),
.B2(n_971),
.Y(n_1231)
);

NOR3xp33_ASAP7_75t_SL g1232 ( 
.A(n_1057),
.B(n_907),
.C(n_906),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1002),
.A2(n_965),
.B1(n_943),
.B2(n_1039),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_931),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_966),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1036),
.A2(n_1053),
.B1(n_1050),
.B2(n_923),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_914),
.A2(n_926),
.B(n_932),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1078),
.A2(n_1052),
.B(n_932),
.Y(n_1238)
);

OR2x6_ASAP7_75t_L g1239 ( 
.A(n_1123),
.B(n_963),
.Y(n_1239)
);

CKINVDCx11_ASAP7_75t_R g1240 ( 
.A(n_1098),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1103),
.B(n_923),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1237),
.A2(n_972),
.B(n_967),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1210),
.B(n_975),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1120),
.A2(n_1052),
.B(n_926),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1091),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1102),
.Y(n_1246)
);

NOR2xp67_ASAP7_75t_L g1247 ( 
.A(n_1200),
.B(n_1000),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1180),
.A2(n_937),
.B(n_1008),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1075),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1215),
.B(n_1037),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1143),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1184),
.A2(n_1027),
.B(n_1043),
.C(n_1037),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1102),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1099),
.B(n_1043),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1125),
.B(n_1032),
.Y(n_1255)
);

O2A1O1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1104),
.A2(n_993),
.B(n_973),
.C(n_882),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1211),
.A2(n_937),
.B(n_1048),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1114),
.B(n_1058),
.Y(n_1258)
);

INVxp67_ASAP7_75t_SL g1259 ( 
.A(n_1128),
.Y(n_1259)
);

AO32x2_ASAP7_75t_L g1260 ( 
.A1(n_1186),
.A2(n_955),
.A3(n_944),
.B1(n_898),
.B2(n_969),
.Y(n_1260)
);

AO21x1_ASAP7_75t_L g1261 ( 
.A1(n_1186),
.A2(n_1010),
.B(n_1018),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1145),
.A2(n_956),
.B1(n_919),
.B2(n_963),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1222),
.A2(n_1020),
.B(n_1022),
.Y(n_1263)
);

AOI221xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1135),
.A2(n_890),
.B1(n_1061),
.B2(n_928),
.C(n_949),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1214),
.A2(n_1026),
.B(n_977),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1118),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1079),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1211),
.A2(n_1004),
.B(n_888),
.Y(n_1268)
);

AOI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1217),
.A2(n_979),
.B(n_991),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1096),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1087),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1093),
.A2(n_1004),
.B(n_954),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1223),
.A2(n_885),
.B(n_952),
.C(n_945),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1229),
.A2(n_1218),
.B(n_1236),
.Y(n_1274)
);

AO31x2_ASAP7_75t_L g1275 ( 
.A1(n_1208),
.A2(n_1229),
.A3(n_1171),
.B(n_1212),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1145),
.A2(n_1111),
.B1(n_1141),
.B2(n_1124),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1094),
.A2(n_1130),
.B(n_1086),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1218),
.A2(n_1085),
.B(n_1140),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1101),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1107),
.B(n_1110),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1100),
.B(n_1193),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_SL g1282 ( 
.A1(n_1097),
.A2(n_1219),
.B(n_1137),
.C(n_1154),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1083),
.A2(n_1233),
.B(n_1084),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1167),
.A2(n_1080),
.B(n_1082),
.C(n_1106),
.Y(n_1284)
);

CKINVDCx8_ASAP7_75t_R g1285 ( 
.A(n_1116),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1117),
.B(n_1193),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1173),
.A2(n_1181),
.B(n_1178),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1175),
.A2(n_1230),
.A3(n_1157),
.B(n_1235),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1188),
.A2(n_1162),
.A3(n_1192),
.B(n_1112),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1160),
.A2(n_1185),
.A3(n_1163),
.B(n_1132),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1131),
.A2(n_1226),
.B1(n_1141),
.B2(n_1134),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1216),
.A2(n_1190),
.B(n_1206),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1174),
.A2(n_1231),
.B(n_1076),
.C(n_1158),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1197),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1233),
.A2(n_1226),
.B(n_1224),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1190),
.A2(n_1213),
.B(n_1225),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1108),
.Y(n_1297)
);

BUFx4_ASAP7_75t_SL g1298 ( 
.A(n_1105),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1089),
.A2(n_1209),
.B(n_1203),
.Y(n_1299)
);

AOI222xp33_ASAP7_75t_L g1300 ( 
.A1(n_1187),
.A2(n_1134),
.B1(n_1191),
.B2(n_1172),
.C1(n_1165),
.C2(n_1116),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1169),
.Y(n_1301)
);

AO22x2_ASAP7_75t_L g1302 ( 
.A1(n_1151),
.A2(n_1202),
.B1(n_1170),
.B2(n_1198),
.Y(n_1302)
);

OA22x2_ASAP7_75t_L g1303 ( 
.A1(n_1088),
.A2(n_1119),
.B1(n_1127),
.B2(n_1109),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1195),
.B(n_1201),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1129),
.B(n_1143),
.Y(n_1305)
);

AOI221x1_ASAP7_75t_L g1306 ( 
.A1(n_1126),
.A2(n_1168),
.B1(n_1138),
.B2(n_1121),
.C(n_1228),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1077),
.A2(n_1123),
.B(n_1159),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1166),
.A2(n_1176),
.B(n_1124),
.C(n_1115),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1081),
.B(n_1090),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1077),
.A2(n_1179),
.A3(n_1182),
.B(n_1126),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1143),
.B(n_1095),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1118),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1194),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1183),
.A2(n_1088),
.B(n_1196),
.C(n_1136),
.Y(n_1314)
);

INVxp67_ASAP7_75t_SL g1315 ( 
.A(n_1139),
.Y(n_1315)
);

O2A1O1Ixp5_ASAP7_75t_L g1316 ( 
.A1(n_1150),
.A2(n_1234),
.B(n_1200),
.C(n_1146),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1095),
.B(n_1074),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1114),
.B(n_1074),
.Y(n_1318)
);

NOR2xp67_ASAP7_75t_SL g1319 ( 
.A(n_1220),
.B(n_1108),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1074),
.B(n_1114),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1077),
.A2(n_1123),
.B(n_1153),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1144),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1142),
.A2(n_1149),
.B(n_1147),
.Y(n_1323)
);

AO32x2_ASAP7_75t_L g1324 ( 
.A1(n_1113),
.A2(n_1148),
.A3(n_1133),
.B1(n_1232),
.B2(n_1092),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1155),
.B(n_1144),
.Y(n_1325)
);

AO32x2_ASAP7_75t_L g1326 ( 
.A1(n_1113),
.A2(n_1205),
.A3(n_1199),
.B1(n_1204),
.B2(n_1234),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1152),
.B(n_1227),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1221),
.B(n_1227),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1221),
.Y(n_1329)
);

AOI221xp5_ASAP7_75t_L g1330 ( 
.A1(n_1122),
.A2(n_1164),
.B1(n_1161),
.B2(n_1113),
.C(n_1177),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1177),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1205),
.B(n_1139),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1152),
.A2(n_1204),
.B(n_1177),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1205),
.A2(n_1189),
.B(n_1204),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1204),
.A2(n_1189),
.B(n_1156),
.Y(n_1335)
);

CKINVDCx11_ASAP7_75t_R g1336 ( 
.A(n_1156),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1189),
.Y(n_1337)
);

AO31x2_ASAP7_75t_L g1338 ( 
.A1(n_1186),
.A2(n_1208),
.A3(n_1222),
.B(n_1217),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1078),
.A2(n_638),
.B(n_590),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1078),
.B(n_886),
.Y(n_1340)
);

AOI221x1_ASAP7_75t_L g1341 ( 
.A1(n_1078),
.A2(n_1186),
.B1(n_1229),
.B2(n_1226),
.C(n_1167),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1237),
.A2(n_972),
.B(n_942),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1125),
.B(n_842),
.Y(n_1343)
);

AOI31xp67_ASAP7_75t_L g1344 ( 
.A1(n_1214),
.A2(n_1217),
.A3(n_1208),
.B(n_1056),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1102),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1078),
.A2(n_638),
.B(n_590),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1075),
.Y(n_1347)
);

OAI22x1_ASAP7_75t_L g1348 ( 
.A1(n_1088),
.A2(n_880),
.B1(n_910),
.B2(n_636),
.Y(n_1348)
);

INVx3_ASAP7_75t_L g1349 ( 
.A(n_1108),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1078),
.A2(n_638),
.B(n_590),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1078),
.A2(n_638),
.B(n_590),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1078),
.B(n_886),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1075),
.Y(n_1353)
);

OAI22x1_ASAP7_75t_L g1354 ( 
.A1(n_1088),
.A2(n_880),
.B1(n_910),
.B2(n_636),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1078),
.A2(n_638),
.B(n_590),
.Y(n_1355)
);

O2A1O1Ixp5_ASAP7_75t_SL g1356 ( 
.A1(n_1186),
.A2(n_1078),
.B(n_1207),
.C(n_1235),
.Y(n_1356)
);

AO31x2_ASAP7_75t_L g1357 ( 
.A1(n_1186),
.A2(n_1208),
.A3(n_1222),
.B(n_1217),
.Y(n_1357)
);

O2A1O1Ixp5_ASAP7_75t_SL g1358 ( 
.A1(n_1186),
.A2(n_1078),
.B(n_1207),
.C(n_1235),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1078),
.A2(n_891),
.B(n_886),
.C(n_711),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1091),
.Y(n_1360)
);

BUFx12f_ASAP7_75t_L g1361 ( 
.A(n_1091),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1091),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_SL g1363 ( 
.A1(n_1078),
.A2(n_978),
.B(n_1130),
.C(n_904),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1078),
.B(n_886),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_SL g1365 ( 
.A(n_1145),
.B(n_1226),
.Y(n_1365)
);

A2O1A1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1078),
.A2(n_880),
.B(n_891),
.C(n_886),
.Y(n_1366)
);

AO21x2_ASAP7_75t_L g1367 ( 
.A1(n_1186),
.A2(n_1208),
.B(n_1222),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1078),
.A2(n_638),
.B(n_590),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1186),
.A2(n_1208),
.A3(n_1222),
.B(n_1217),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1078),
.A2(n_638),
.B(n_590),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1143),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1237),
.A2(n_972),
.B(n_942),
.Y(n_1372)
);

NAND2x1p5_ASAP7_75t_L g1373 ( 
.A(n_1114),
.B(n_894),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1237),
.A2(n_972),
.B(n_942),
.Y(n_1374)
);

NOR2x1_ASAP7_75t_R g1375 ( 
.A(n_1091),
.B(n_665),
.Y(n_1375)
);

NOR2x1_ASAP7_75t_L g1376 ( 
.A(n_1099),
.B(n_1130),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1078),
.A2(n_886),
.B1(n_891),
.B2(n_880),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1091),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_1128),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1087),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1078),
.A2(n_638),
.B(n_590),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1075),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1078),
.A2(n_978),
.B1(n_891),
.B2(n_886),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1078),
.A2(n_880),
.B(n_891),
.C(n_886),
.Y(n_1384)
);

O2A1O1Ixp5_ASAP7_75t_SL g1385 ( 
.A1(n_1186),
.A2(n_1078),
.B(n_1207),
.C(n_1235),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1078),
.A2(n_638),
.B(n_590),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1078),
.B(n_886),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1222),
.A2(n_1217),
.B(n_1214),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1075),
.Y(n_1389)
);

BUFx10_ASAP7_75t_L g1390 ( 
.A(n_1091),
.Y(n_1390)
);

AOI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1214),
.A2(n_1019),
.B(n_1015),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1078),
.A2(n_880),
.B(n_891),
.C(n_886),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1078),
.A2(n_638),
.B(n_590),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1125),
.B(n_842),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1186),
.A2(n_1208),
.B(n_1222),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1078),
.B(n_904),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1222),
.A2(n_1217),
.B(n_1214),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_SL g1398 ( 
.A1(n_1078),
.A2(n_978),
.B(n_1130),
.C(n_904),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1237),
.A2(n_972),
.B(n_942),
.Y(n_1399)
);

BUFx4f_ASAP7_75t_SL g1400 ( 
.A(n_1118),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_SL g1401 ( 
.A1(n_1078),
.A2(n_978),
.B(n_1130),
.C(n_904),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1078),
.A2(n_891),
.B(n_886),
.C(n_711),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1102),
.Y(n_1403)
);

A2O1A1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1078),
.A2(n_880),
.B(n_891),
.C(n_886),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1237),
.A2(n_972),
.B(n_942),
.Y(n_1405)
);

INVx5_ASAP7_75t_L g1406 ( 
.A(n_1204),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1365),
.A2(n_1348),
.B1(n_1354),
.B2(n_1291),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1366),
.A2(n_1392),
.B(n_1384),
.Y(n_1408)
);

INVx8_ASAP7_75t_L g1409 ( 
.A(n_1361),
.Y(n_1409)
);

OAI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1365),
.A2(n_1377),
.B1(n_1341),
.B2(n_1285),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1377),
.A2(n_1352),
.B1(n_1340),
.B2(n_1387),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1300),
.A2(n_1276),
.B1(n_1376),
.B2(n_1254),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1383),
.A2(n_1364),
.B1(n_1274),
.B2(n_1303),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1404),
.A2(n_1383),
.B(n_1300),
.Y(n_1414)
);

INVx6_ASAP7_75t_L g1415 ( 
.A(n_1390),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1267),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1270),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1336),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1396),
.A2(n_1402),
.B1(n_1359),
.B2(n_1274),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1312),
.Y(n_1420)
);

INVx6_ASAP7_75t_L g1421 ( 
.A(n_1390),
.Y(n_1421)
);

OAI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1295),
.A2(n_1396),
.B1(n_1376),
.B2(n_1394),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1302),
.A2(n_1278),
.B1(n_1379),
.B2(n_1259),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1380),
.Y(n_1424)
);

OAI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1328),
.A2(n_1250),
.B1(n_1329),
.B2(n_1301),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1240),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_1400),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1363),
.B(n_1398),
.Y(n_1428)
);

CKINVDCx11_ASAP7_75t_R g1429 ( 
.A(n_1345),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1347),
.Y(n_1430)
);

INVx4_ASAP7_75t_L g1431 ( 
.A(n_1403),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1353),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1245),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1302),
.A2(n_1278),
.B1(n_1271),
.B2(n_1286),
.Y(n_1434)
);

CKINVDCx6p67_ASAP7_75t_R g1435 ( 
.A(n_1343),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1308),
.A2(n_1284),
.B1(n_1314),
.B2(n_1293),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1360),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1382),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1281),
.A2(n_1258),
.B1(n_1309),
.B2(n_1389),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1280),
.B(n_1304),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1290),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1279),
.B(n_1305),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1258),
.A2(n_1241),
.B1(n_1313),
.B2(n_1255),
.Y(n_1443)
);

INVx4_ASAP7_75t_L g1444 ( 
.A(n_1362),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1378),
.Y(n_1445)
);

NAND2x1p5_ASAP7_75t_L g1446 ( 
.A(n_1406),
.B(n_1335),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1283),
.A2(n_1252),
.B1(n_1406),
.B2(n_1299),
.Y(n_1447)
);

CKINVDCx11_ASAP7_75t_R g1448 ( 
.A(n_1375),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1325),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1332),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1325),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1290),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1266),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1337),
.Y(n_1454)
);

BUFx4f_ASAP7_75t_SL g1455 ( 
.A(n_1246),
.Y(n_1455)
);

BUFx10_ASAP7_75t_L g1456 ( 
.A(n_1331),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1327),
.Y(n_1457)
);

INVx6_ASAP7_75t_L g1458 ( 
.A(n_1251),
.Y(n_1458)
);

INVx6_ASAP7_75t_L g1459 ( 
.A(n_1251),
.Y(n_1459)
);

BUFx8_ASAP7_75t_L g1460 ( 
.A(n_1375),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1243),
.Y(n_1461)
);

CKINVDCx11_ASAP7_75t_R g1462 ( 
.A(n_1371),
.Y(n_1462)
);

CKINVDCx8_ASAP7_75t_R g1463 ( 
.A(n_1371),
.Y(n_1463)
);

NAND2x1p5_ASAP7_75t_L g1464 ( 
.A(n_1406),
.B(n_1327),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1367),
.A2(n_1395),
.B1(n_1330),
.B2(n_1321),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_SL g1466 ( 
.A1(n_1367),
.A2(n_1395),
.B1(n_1326),
.B2(n_1324),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1401),
.B(n_1310),
.Y(n_1467)
);

CKINVDCx6p67_ASAP7_75t_R g1468 ( 
.A(n_1298),
.Y(n_1468)
);

INVx3_ASAP7_75t_SL g1469 ( 
.A(n_1311),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1261),
.A2(n_1307),
.B1(n_1239),
.B2(n_1320),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1239),
.A2(n_1370),
.B1(n_1393),
.B2(n_1386),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1373),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1289),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1310),
.B(n_1315),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1388),
.A2(n_1397),
.B1(n_1323),
.B2(n_1317),
.Y(n_1475)
);

OAI22x1_ASAP7_75t_L g1476 ( 
.A1(n_1324),
.A2(n_1326),
.B1(n_1318),
.B2(n_1397),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1339),
.A2(n_1346),
.B1(n_1350),
.B2(n_1351),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1355),
.A2(n_1368),
.B1(n_1381),
.B2(n_1238),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1256),
.A2(n_1262),
.B1(n_1324),
.B2(n_1349),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1297),
.A2(n_1322),
.B1(n_1349),
.B2(n_1326),
.Y(n_1480)
);

BUFx4f_ASAP7_75t_SL g1481 ( 
.A(n_1322),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1388),
.A2(n_1334),
.B1(n_1263),
.B2(n_1244),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1333),
.Y(n_1483)
);

OAI21xp33_ASAP7_75t_L g1484 ( 
.A1(n_1356),
.A2(n_1385),
.B(n_1358),
.Y(n_1484)
);

CKINVDCx11_ASAP7_75t_R g1485 ( 
.A(n_1319),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1310),
.B(n_1338),
.Y(n_1486)
);

BUFx10_ASAP7_75t_L g1487 ( 
.A(n_1316),
.Y(n_1487)
);

CKINVDCx10_ASAP7_75t_R g1488 ( 
.A(n_1306),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1344),
.Y(n_1489)
);

BUFx2_ASAP7_75t_SL g1490 ( 
.A(n_1247),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1275),
.A2(n_1292),
.B1(n_1263),
.B2(n_1268),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1248),
.A2(n_1277),
.B1(n_1247),
.B2(n_1257),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1272),
.A2(n_1265),
.B1(n_1296),
.B2(n_1405),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1275),
.A2(n_1260),
.B1(n_1338),
.B2(n_1369),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1288),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_SL g1496 ( 
.A(n_1282),
.Y(n_1496)
);

INVx6_ASAP7_75t_SL g1497 ( 
.A(n_1273),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1342),
.A2(n_1399),
.B1(n_1374),
.B2(n_1372),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1357),
.B(n_1369),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1369),
.B(n_1275),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1269),
.A2(n_1391),
.B1(n_1264),
.B2(n_1260),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1264),
.A2(n_1287),
.B1(n_1242),
.B2(n_1260),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1288),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1288),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1280),
.Y(n_1505)
);

INVx6_ASAP7_75t_L g1506 ( 
.A(n_1390),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1249),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1365),
.A2(n_880),
.B1(n_910),
.B2(n_1377),
.Y(n_1508)
);

CKINVDCx14_ASAP7_75t_R g1509 ( 
.A(n_1336),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1280),
.Y(n_1510)
);

INVx3_ASAP7_75t_SL g1511 ( 
.A(n_1245),
.Y(n_1511)
);

INVx6_ASAP7_75t_L g1512 ( 
.A(n_1390),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1249),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1249),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1312),
.Y(n_1515)
);

CKINVDCx8_ASAP7_75t_R g1516 ( 
.A(n_1245),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1249),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1249),
.Y(n_1518)
);

BUFx12f_ASAP7_75t_L g1519 ( 
.A(n_1336),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1249),
.Y(n_1520)
);

INVx5_ASAP7_75t_L g1521 ( 
.A(n_1406),
.Y(n_1521)
);

BUFx10_ASAP7_75t_L g1522 ( 
.A(n_1245),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1365),
.A2(n_1186),
.B1(n_1145),
.B2(n_1383),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1365),
.A2(n_1354),
.B1(n_1348),
.B2(n_1291),
.Y(n_1524)
);

CKINVDCx11_ASAP7_75t_R g1525 ( 
.A(n_1336),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1365),
.A2(n_891),
.B1(n_886),
.B2(n_1099),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1294),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1377),
.A2(n_1352),
.B1(n_1364),
.B2(n_1340),
.Y(n_1528)
);

INVx2_ASAP7_75t_SL g1529 ( 
.A(n_1298),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1253),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1249),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1377),
.A2(n_1352),
.B1(n_1364),
.B2(n_1340),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1253),
.Y(n_1533)
);

BUFx10_ASAP7_75t_L g1534 ( 
.A(n_1245),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1365),
.A2(n_1186),
.B1(n_1145),
.B2(n_1383),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_1336),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1249),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1336),
.Y(n_1538)
);

BUFx8_ASAP7_75t_L g1539 ( 
.A(n_1361),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1294),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1365),
.A2(n_1354),
.B1(n_1348),
.B2(n_1291),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1249),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1365),
.A2(n_891),
.B1(n_886),
.B2(n_1099),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1249),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1365),
.A2(n_1354),
.B1(n_1348),
.B2(n_1291),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1249),
.Y(n_1546)
);

BUFx8_ASAP7_75t_L g1547 ( 
.A(n_1361),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1365),
.A2(n_1354),
.B1(n_1348),
.B2(n_1291),
.Y(n_1548)
);

OAI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1365),
.A2(n_880),
.B1(n_910),
.B2(n_1377),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1249),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1249),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1280),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1483),
.B(n_1500),
.Y(n_1553)
);

AO21x2_ASAP7_75t_L g1554 ( 
.A1(n_1499),
.A2(n_1504),
.B(n_1503),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1489),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1528),
.B(n_1532),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1461),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1474),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1528),
.B(n_1532),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1473),
.Y(n_1560)
);

OA21x2_ASAP7_75t_L g1561 ( 
.A1(n_1465),
.A2(n_1486),
.B(n_1502),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1449),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1497),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1505),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1441),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1452),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1456),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1510),
.B(n_1411),
.Y(n_1568)
);

AO21x2_ASAP7_75t_L g1569 ( 
.A1(n_1499),
.A2(n_1467),
.B(n_1486),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1474),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1467),
.Y(n_1571)
);

OA21x2_ASAP7_75t_L g1572 ( 
.A1(n_1492),
.A2(n_1493),
.B(n_1484),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1523),
.A2(n_1535),
.B1(n_1413),
.B2(n_1549),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1435),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1416),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1417),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1430),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1521),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1497),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1511),
.B(n_1444),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1521),
.B(n_1495),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1432),
.Y(n_1582)
);

INVx4_ASAP7_75t_L g1583 ( 
.A(n_1521),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1495),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1464),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1466),
.B(n_1438),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1466),
.B(n_1507),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1513),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1514),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1517),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1470),
.B(n_1408),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1451),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1518),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1414),
.A2(n_1543),
.B(n_1526),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1456),
.Y(n_1595)
);

O2A1O1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1414),
.A2(n_1508),
.B(n_1410),
.C(n_1436),
.Y(n_1596)
);

NOR2x1_ASAP7_75t_L g1597 ( 
.A(n_1422),
.B(n_1447),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1520),
.B(n_1531),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1552),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1477),
.A2(n_1478),
.B(n_1471),
.Y(n_1600)
);

AO21x2_ASAP7_75t_L g1601 ( 
.A1(n_1501),
.A2(n_1479),
.B(n_1477),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1537),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1551),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1542),
.B(n_1544),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1546),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1480),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1450),
.B(n_1419),
.Y(n_1607)
);

OR2x6_ASAP7_75t_L g1608 ( 
.A(n_1446),
.B(n_1476),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1550),
.Y(n_1609)
);

INVxp67_ASAP7_75t_L g1610 ( 
.A(n_1440),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1501),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1419),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1494),
.B(n_1408),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1413),
.B(n_1425),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1480),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1442),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1475),
.B(n_1482),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1494),
.Y(n_1618)
);

OA21x2_ASAP7_75t_L g1619 ( 
.A1(n_1498),
.A2(n_1428),
.B(n_1478),
.Y(n_1619)
);

AOI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1428),
.A2(n_1447),
.B(n_1479),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1523),
.A2(n_1535),
.B1(n_1412),
.B2(n_1436),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1424),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1454),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1471),
.A2(n_1446),
.B(n_1548),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1491),
.A2(n_1407),
.B(n_1524),
.Y(n_1625)
);

NAND2x1p5_ASAP7_75t_L g1626 ( 
.A(n_1450),
.B(n_1457),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1541),
.B(n_1545),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1434),
.A2(n_1423),
.B1(n_1439),
.B2(n_1443),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1527),
.Y(n_1629)
);

OA21x2_ASAP7_75t_L g1630 ( 
.A1(n_1540),
.A2(n_1491),
.B(n_1488),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1469),
.B(n_1487),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1487),
.B(n_1490),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1496),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1415),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_1463),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1496),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1415),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1421),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1481),
.Y(n_1639)
);

AOI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1485),
.A2(n_1458),
.B(n_1459),
.Y(n_1640)
);

AOI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1462),
.A2(n_1529),
.B(n_1472),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1530),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1431),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1420),
.A2(n_1515),
.B1(n_1429),
.B2(n_1533),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1506),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1533),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1506),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1431),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1512),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1512),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1455),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1433),
.B(n_1437),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1409),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1453),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1522),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1409),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1409),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1534),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1468),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1539),
.Y(n_1660)
);

AO31x2_ASAP7_75t_L g1661 ( 
.A1(n_1460),
.A2(n_1448),
.A3(n_1547),
.B(n_1539),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1547),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1460),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1516),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1564),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1594),
.B(n_1426),
.C(n_1509),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1616),
.B(n_1519),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1594),
.A2(n_1418),
.B1(n_1536),
.B2(n_1538),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1610),
.B(n_1525),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1556),
.B(n_1445),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1596),
.A2(n_1427),
.B(n_1621),
.C(n_1597),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1605),
.Y(n_1672)
);

AOI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1573),
.A2(n_1559),
.B1(n_1621),
.B2(n_1613),
.C(n_1612),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1612),
.B(n_1607),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_SL g1675 ( 
.A1(n_1591),
.A2(n_1614),
.B(n_1635),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1597),
.A2(n_1600),
.B(n_1601),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1607),
.B(n_1613),
.Y(n_1677)
);

A2O1A1Ixp33_ASAP7_75t_L g1678 ( 
.A1(n_1625),
.A2(n_1591),
.B(n_1627),
.C(n_1568),
.Y(n_1678)
);

AO32x2_ASAP7_75t_L g1679 ( 
.A1(n_1567),
.A2(n_1595),
.A3(n_1645),
.B1(n_1638),
.B2(n_1634),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1591),
.A2(n_1636),
.B(n_1633),
.C(n_1579),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1623),
.B(n_1599),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1553),
.B(n_1562),
.Y(n_1682)
);

AOI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1591),
.A2(n_1606),
.B1(n_1615),
.B2(n_1627),
.C(n_1618),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1592),
.B(n_1598),
.Y(n_1684)
);

OA21x2_ASAP7_75t_L g1685 ( 
.A1(n_1624),
.A2(n_1611),
.B(n_1558),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1557),
.B(n_1615),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1592),
.B(n_1598),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1592),
.B(n_1604),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1604),
.B(n_1631),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1631),
.B(n_1652),
.Y(n_1690)
);

O2A1O1Ixp33_ASAP7_75t_L g1691 ( 
.A1(n_1633),
.A2(n_1636),
.B(n_1579),
.C(n_1648),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1570),
.B(n_1571),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1570),
.B(n_1571),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1628),
.A2(n_1620),
.B1(n_1563),
.B2(n_1630),
.Y(n_1694)
);

AO32x2_ASAP7_75t_L g1695 ( 
.A1(n_1637),
.A2(n_1578),
.A3(n_1583),
.B1(n_1586),
.B2(n_1587),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1563),
.A2(n_1630),
.B1(n_1574),
.B2(n_1582),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1575),
.A2(n_1602),
.B1(n_1582),
.B2(n_1588),
.C(n_1589),
.Y(n_1697)
);

AND2x6_ASAP7_75t_L g1698 ( 
.A(n_1632),
.B(n_1585),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1630),
.A2(n_1603),
.B1(n_1576),
.B2(n_1577),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1553),
.B(n_1608),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1601),
.A2(n_1577),
.B1(n_1602),
.B2(n_1593),
.C(n_1590),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1572),
.A2(n_1619),
.B(n_1617),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1646),
.B(n_1643),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1664),
.B(n_1651),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1630),
.A2(n_1609),
.B1(n_1644),
.B2(n_1635),
.Y(n_1705)
);

CKINVDCx8_ASAP7_75t_R g1706 ( 
.A(n_1654),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_SL g1707 ( 
.A1(n_1617),
.A2(n_1601),
.B1(n_1561),
.B2(n_1608),
.Y(n_1707)
);

AO32x2_ASAP7_75t_L g1708 ( 
.A1(n_1626),
.A2(n_1569),
.A3(n_1561),
.B1(n_1622),
.B2(n_1629),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1569),
.A2(n_1617),
.B1(n_1642),
.B2(n_1655),
.C(n_1658),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1584),
.A2(n_1566),
.B(n_1565),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1674),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1700),
.B(n_1581),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1665),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1710),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1701),
.B(n_1619),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1673),
.A2(n_1561),
.B1(n_1572),
.B2(n_1608),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1672),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1673),
.A2(n_1619),
.B1(n_1561),
.B2(n_1655),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1686),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1677),
.B(n_1619),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1686),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1701),
.B(n_1572),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1695),
.B(n_1555),
.Y(n_1723)
);

NOR2x1_ASAP7_75t_L g1724 ( 
.A(n_1691),
.B(n_1658),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1683),
.A2(n_1572),
.B1(n_1662),
.B2(n_1660),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1695),
.B(n_1555),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1695),
.B(n_1555),
.Y(n_1727)
);

CKINVDCx20_ASAP7_75t_R g1728 ( 
.A(n_1706),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1692),
.B(n_1554),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1684),
.B(n_1554),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1698),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1683),
.A2(n_1662),
.B1(n_1660),
.B2(n_1654),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1687),
.B(n_1554),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1688),
.B(n_1554),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1689),
.B(n_1702),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1679),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1708),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1708),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1703),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1693),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1676),
.B(n_1560),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1685),
.Y(n_1742)
);

INVxp67_ASAP7_75t_SL g1743 ( 
.A(n_1742),
.Y(n_1743)
);

BUFx6f_ASAP7_75t_L g1744 ( 
.A(n_1731),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1720),
.B(n_1681),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1728),
.B(n_1660),
.Y(n_1746)
);

AOI21xp33_ASAP7_75t_L g1747 ( 
.A1(n_1722),
.A2(n_1671),
.B(n_1709),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1717),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1711),
.B(n_1697),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1717),
.Y(n_1750)
);

BUFx2_ASAP7_75t_L g1751 ( 
.A(n_1731),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1713),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1713),
.B(n_1668),
.Y(n_1753)
);

INVxp67_ASAP7_75t_SL g1754 ( 
.A(n_1742),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1724),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1735),
.B(n_1690),
.Y(n_1756)
);

OAI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1715),
.A2(n_1678),
.B1(n_1707),
.B2(n_1699),
.C(n_1696),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1731),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1732),
.A2(n_1694),
.B1(n_1699),
.B2(n_1705),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1723),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1719),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1735),
.B(n_1682),
.Y(n_1762)
);

OAI21xp33_ASAP7_75t_L g1763 ( 
.A1(n_1715),
.A2(n_1668),
.B(n_1666),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1735),
.B(n_1682),
.Y(n_1764)
);

OAI33xp33_ASAP7_75t_L g1765 ( 
.A1(n_1718),
.A2(n_1694),
.A3(n_1705),
.B1(n_1696),
.B2(n_1670),
.B3(n_1666),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1721),
.Y(n_1766)
);

INVx5_ASAP7_75t_L g1767 ( 
.A(n_1714),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1723),
.Y(n_1768)
);

AO21x2_ASAP7_75t_L g1769 ( 
.A1(n_1722),
.A2(n_1737),
.B(n_1738),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1736),
.B(n_1679),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1718),
.A2(n_1675),
.B1(n_1680),
.B2(n_1670),
.C(n_1704),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1721),
.Y(n_1772)
);

NAND2x1_ASAP7_75t_L g1773 ( 
.A(n_1723),
.B(n_1698),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1739),
.B(n_1679),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1743),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1760),
.B(n_1768),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1760),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1754),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1765),
.A2(n_1716),
.B1(n_1725),
.B2(n_1732),
.Y(n_1779)
);

INVx1_ASAP7_75t_SL g1780 ( 
.A(n_1751),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1760),
.B(n_1768),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1760),
.B(n_1768),
.Y(n_1782)
);

INVx2_ASAP7_75t_SL g1783 ( 
.A(n_1767),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1748),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1770),
.B(n_1726),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1751),
.Y(n_1786)
);

AND2x6_ASAP7_75t_SL g1787 ( 
.A(n_1746),
.B(n_1663),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1770),
.B(n_1726),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1761),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1749),
.B(n_1740),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1748),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1774),
.B(n_1727),
.Y(n_1792)
);

NAND2x1p5_ASAP7_75t_L g1793 ( 
.A(n_1767),
.B(n_1773),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1774),
.B(n_1727),
.Y(n_1794)
);

NOR2x1p5_ASAP7_75t_L g1795 ( 
.A(n_1773),
.B(n_1656),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1766),
.Y(n_1796)
);

NAND3xp33_ASAP7_75t_SL g1797 ( 
.A(n_1763),
.B(n_1725),
.C(n_1716),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1767),
.B(n_1727),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1756),
.B(n_1730),
.Y(n_1799)
);

NAND2xp33_ASAP7_75t_R g1800 ( 
.A(n_1749),
.B(n_1741),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1756),
.B(n_1730),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1767),
.B(n_1712),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1767),
.B(n_1730),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1772),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1750),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1772),
.B(n_1740),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1767),
.B(n_1733),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1769),
.B(n_1729),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1784),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1784),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1784),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1791),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1791),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1799),
.B(n_1762),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1791),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1799),
.B(n_1762),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1799),
.B(n_1764),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1805),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1789),
.Y(n_1819)
);

INVxp67_ASAP7_75t_L g1820 ( 
.A(n_1790),
.Y(n_1820)
);

AND4x1_ASAP7_75t_L g1821 ( 
.A(n_1779),
.B(n_1763),
.C(n_1771),
.D(n_1753),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1801),
.B(n_1758),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1790),
.B(n_1755),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1782),
.Y(n_1824)
);

OR2x6_ASAP7_75t_L g1825 ( 
.A(n_1793),
.B(n_1640),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1805),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1801),
.B(n_1758),
.Y(n_1827)
);

NAND2x1_ASAP7_75t_L g1828 ( 
.A(n_1802),
.B(n_1744),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1801),
.B(n_1795),
.Y(n_1829)
);

AOI32xp33_ASAP7_75t_L g1830 ( 
.A1(n_1779),
.A2(n_1792),
.A3(n_1794),
.B1(n_1785),
.B2(n_1788),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1806),
.B(n_1752),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1805),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1782),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1804),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1782),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1782),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1780),
.B(n_1734),
.Y(n_1837)
);

INVxp67_ASAP7_75t_L g1838 ( 
.A(n_1800),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1806),
.B(n_1789),
.Y(n_1839)
);

OAI21xp33_ASAP7_75t_SL g1840 ( 
.A1(n_1795),
.A2(n_1781),
.B(n_1776),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1804),
.Y(n_1841)
);

NAND2x2_ASAP7_75t_L g1842 ( 
.A(n_1795),
.B(n_1656),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1796),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1801),
.B(n_1802),
.Y(n_1844)
);

OAI21xp33_ASAP7_75t_L g1845 ( 
.A1(n_1797),
.A2(n_1747),
.B(n_1759),
.Y(n_1845)
);

OR2x6_ASAP7_75t_L g1846 ( 
.A(n_1793),
.B(n_1783),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1802),
.B(n_1758),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1780),
.B(n_1734),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1802),
.B(n_1785),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1796),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1786),
.B(n_1745),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1822),
.B(n_1786),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1845),
.B(n_1820),
.Y(n_1853)
);

INVx1_ASAP7_75t_SL g1854 ( 
.A(n_1847),
.Y(n_1854)
);

OAI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1838),
.A2(n_1797),
.B(n_1747),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1809),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1822),
.B(n_1802),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1823),
.A2(n_1757),
.B(n_1775),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1809),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1821),
.B(n_1775),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1839),
.B(n_1785),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1824),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1827),
.B(n_1802),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1827),
.B(n_1793),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1810),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1814),
.B(n_1793),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1830),
.B(n_1775),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1810),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1814),
.B(n_1793),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1811),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1849),
.B(n_1846),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1839),
.B(n_1831),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_SL g1873 ( 
.A1(n_1829),
.A2(n_1800),
.B1(n_1794),
.B2(n_1792),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1819),
.B(n_1778),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1811),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1812),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1831),
.B(n_1785),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1847),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1812),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1843),
.B(n_1788),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1843),
.B(n_1778),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1816),
.B(n_1803),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1840),
.B(n_1787),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1816),
.B(n_1803),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1817),
.B(n_1803),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1849),
.B(n_1783),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1850),
.B(n_1788),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1824),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1856),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1886),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1856),
.Y(n_1891)
);

NAND3x2_ASAP7_75t_L g1892 ( 
.A(n_1871),
.B(n_1778),
.C(n_1829),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1860),
.A2(n_1828),
.B(n_1846),
.Y(n_1893)
);

AOI211xp5_ASAP7_75t_L g1894 ( 
.A1(n_1855),
.A2(n_1803),
.B(n_1807),
.C(n_1783),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1859),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1858),
.A2(n_1853),
.B(n_1867),
.Y(n_1896)
);

AOI211xp5_ASAP7_75t_L g1897 ( 
.A1(n_1883),
.A2(n_1807),
.B(n_1783),
.C(n_1841),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1877),
.B(n_1850),
.Y(n_1898)
);

INVxp67_ASAP7_75t_L g1899 ( 
.A(n_1874),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1859),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1865),
.Y(n_1901)
);

AND2x4_ASAP7_75t_SL g1902 ( 
.A(n_1871),
.B(n_1667),
.Y(n_1902)
);

NAND3xp33_ASAP7_75t_L g1903 ( 
.A(n_1873),
.B(n_1881),
.C(n_1834),
.Y(n_1903)
);

AOI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1852),
.A2(n_1828),
.B(n_1846),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1872),
.B(n_1841),
.Y(n_1905)
);

NAND2x1_ASAP7_75t_L g1906 ( 
.A(n_1871),
.B(n_1846),
.Y(n_1906)
);

OAI31xp33_ASAP7_75t_L g1907 ( 
.A1(n_1880),
.A2(n_1808),
.A3(n_1794),
.B(n_1792),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1865),
.Y(n_1908)
);

OAI22xp33_ASAP7_75t_L g1909 ( 
.A1(n_1877),
.A2(n_1759),
.B1(n_1825),
.B2(n_1842),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1872),
.B(n_1788),
.Y(n_1910)
);

OAI332xp33_ASAP7_75t_L g1911 ( 
.A1(n_1861),
.A2(n_1887),
.A3(n_1880),
.B1(n_1854),
.B2(n_1878),
.B3(n_1808),
.C1(n_1888),
.C2(n_1862),
.Y(n_1911)
);

AOI21xp33_ASAP7_75t_L g1912 ( 
.A1(n_1868),
.A2(n_1808),
.B(n_1769),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1868),
.Y(n_1913)
);

AOI221xp5_ASAP7_75t_L g1914 ( 
.A1(n_1862),
.A2(n_1769),
.B1(n_1792),
.B2(n_1794),
.C(n_1837),
.Y(n_1914)
);

OAI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1896),
.A2(n_1852),
.B(n_1871),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1899),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1894),
.B(n_1886),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1905),
.Y(n_1918)
);

BUFx3_ASAP7_75t_L g1919 ( 
.A(n_1902),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1889),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1911),
.B(n_1861),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1890),
.B(n_1864),
.Y(n_1922)
);

OAI211xp5_ASAP7_75t_L g1923 ( 
.A1(n_1892),
.A2(n_1864),
.B(n_1887),
.C(n_1866),
.Y(n_1923)
);

AOI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1914),
.A2(n_1888),
.B1(n_1862),
.B2(n_1876),
.C(n_1870),
.Y(n_1924)
);

OAI32xp33_ASAP7_75t_L g1925 ( 
.A1(n_1903),
.A2(n_1866),
.A3(n_1869),
.B1(n_1857),
.B2(n_1863),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1891),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1895),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1910),
.B(n_1851),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1906),
.A2(n_1886),
.B(n_1875),
.Y(n_1929)
);

NAND2xp33_ASAP7_75t_SL g1930 ( 
.A(n_1905),
.B(n_1869),
.Y(n_1930)
);

AOI21xp33_ASAP7_75t_L g1931 ( 
.A1(n_1900),
.A2(n_1888),
.B(n_1875),
.Y(n_1931)
);

AOI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1909),
.A2(n_1825),
.B1(n_1737),
.B2(n_1738),
.Y(n_1932)
);

OAI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1912),
.A2(n_1886),
.B(n_1724),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1901),
.Y(n_1934)
);

NAND2xp33_ASAP7_75t_SL g1935 ( 
.A(n_1916),
.B(n_1898),
.Y(n_1935)
);

OAI21xp33_ASAP7_75t_L g1936 ( 
.A1(n_1921),
.A2(n_1910),
.B(n_1897),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1916),
.Y(n_1937)
);

INVxp67_ASAP7_75t_L g1938 ( 
.A(n_1919),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1915),
.B(n_1857),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1920),
.Y(n_1940)
);

XOR2x2_ASAP7_75t_L g1941 ( 
.A(n_1919),
.B(n_1641),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1926),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1927),
.Y(n_1943)
);

O2A1O1Ixp33_ASAP7_75t_L g1944 ( 
.A1(n_1918),
.A2(n_1912),
.B(n_1913),
.C(n_1908),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1931),
.B(n_1870),
.Y(n_1945)
);

OAI221xp5_ASAP7_75t_L g1946 ( 
.A1(n_1924),
.A2(n_1907),
.B1(n_1893),
.B2(n_1825),
.C(n_1904),
.Y(n_1946)
);

OAI211xp5_ASAP7_75t_SL g1947 ( 
.A1(n_1936),
.A2(n_1923),
.B(n_1917),
.C(n_1933),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1937),
.Y(n_1948)
);

A2O1A1Ixp33_ASAP7_75t_L g1949 ( 
.A1(n_1944),
.A2(n_1932),
.B(n_1930),
.C(n_1925),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1935),
.B(n_1928),
.Y(n_1950)
);

INVxp67_ASAP7_75t_SL g1951 ( 
.A(n_1938),
.Y(n_1951)
);

INVxp67_ASAP7_75t_SL g1952 ( 
.A(n_1945),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1939),
.B(n_1922),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1940),
.B(n_1934),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1941),
.Y(n_1955)
);

NAND3xp33_ASAP7_75t_L g1956 ( 
.A(n_1945),
.B(n_1930),
.C(n_1929),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1942),
.Y(n_1957)
);

AOI211xp5_ASAP7_75t_L g1958 ( 
.A1(n_1947),
.A2(n_1946),
.B(n_1917),
.C(n_1943),
.Y(n_1958)
);

AOI221xp5_ASAP7_75t_L g1959 ( 
.A1(n_1952),
.A2(n_1876),
.B1(n_1879),
.B2(n_1815),
.C(n_1813),
.Y(n_1959)
);

NOR3xp33_ASAP7_75t_L g1960 ( 
.A(n_1952),
.B(n_1641),
.C(n_1659),
.Y(n_1960)
);

AOI22xp33_ASAP7_75t_SL g1961 ( 
.A1(n_1956),
.A2(n_1825),
.B1(n_1879),
.B2(n_1863),
.Y(n_1961)
);

O2A1O1Ixp5_ASAP7_75t_L g1962 ( 
.A1(n_1949),
.A2(n_1951),
.B(n_1950),
.C(n_1953),
.Y(n_1962)
);

AOI211xp5_ASAP7_75t_L g1963 ( 
.A1(n_1955),
.A2(n_1885),
.B(n_1884),
.C(n_1882),
.Y(n_1963)
);

NAND4xp75_ASAP7_75t_L g1964 ( 
.A(n_1948),
.B(n_1954),
.C(n_1957),
.D(n_1885),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1951),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1965),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1963),
.B(n_1787),
.Y(n_1967)
);

NOR3xp33_ASAP7_75t_SL g1968 ( 
.A(n_1964),
.B(n_1580),
.C(n_1661),
.Y(n_1968)
);

OAI221xp5_ASAP7_75t_L g1969 ( 
.A1(n_1960),
.A2(n_1842),
.B1(n_1835),
.B2(n_1836),
.C(n_1833),
.Y(n_1969)
);

AOI211xp5_ASAP7_75t_L g1970 ( 
.A1(n_1958),
.A2(n_1656),
.B(n_1657),
.C(n_1884),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1962),
.B(n_1961),
.Y(n_1971)
);

AOI221xp5_ASAP7_75t_L g1972 ( 
.A1(n_1959),
.A2(n_1813),
.B1(n_1818),
.B2(n_1826),
.C(n_1832),
.Y(n_1972)
);

AOI221xp5_ASAP7_75t_L g1973 ( 
.A1(n_1962),
.A2(n_1832),
.B1(n_1818),
.B2(n_1826),
.C(n_1815),
.Y(n_1973)
);

NOR2x1_ASAP7_75t_L g1974 ( 
.A(n_1971),
.B(n_1657),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1966),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1967),
.Y(n_1976)
);

NAND4xp75_ASAP7_75t_L g1977 ( 
.A(n_1968),
.B(n_1973),
.C(n_1972),
.D(n_1970),
.Y(n_1977)
);

XNOR2xp5_ASAP7_75t_L g1978 ( 
.A(n_1969),
.B(n_1657),
.Y(n_1978)
);

XNOR2x1_ASAP7_75t_L g1979 ( 
.A(n_1966),
.B(n_1661),
.Y(n_1979)
);

O2A1O1Ixp33_ASAP7_75t_L g1980 ( 
.A1(n_1975),
.A2(n_1833),
.B(n_1836),
.C(n_1835),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1976),
.A2(n_1882),
.B1(n_1798),
.B2(n_1844),
.Y(n_1981)
);

OA22x2_ASAP7_75t_L g1982 ( 
.A1(n_1978),
.A2(n_1651),
.B1(n_1669),
.B2(n_1653),
.Y(n_1982)
);

HB1xp67_ASAP7_75t_L g1983 ( 
.A(n_1982),
.Y(n_1983)
);

OAI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1983),
.A2(n_1974),
.B1(n_1981),
.B2(n_1977),
.Y(n_1984)
);

AOI22x1_ASAP7_75t_L g1985 ( 
.A1(n_1984),
.A2(n_1979),
.B1(n_1980),
.B2(n_1651),
.Y(n_1985)
);

OAI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1984),
.A2(n_1844),
.B1(n_1848),
.B2(n_1777),
.Y(n_1986)
);

AOI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1986),
.A2(n_1777),
.B1(n_1653),
.B2(n_1798),
.Y(n_1987)
);

XNOR2xp5_ASAP7_75t_L g1988 ( 
.A(n_1985),
.B(n_1661),
.Y(n_1988)
);

OAI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1987),
.A2(n_1777),
.B1(n_1653),
.B2(n_1661),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1988),
.Y(n_1990)
);

XNOR2xp5_ASAP7_75t_L g1991 ( 
.A(n_1990),
.B(n_1661),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1991),
.A2(n_1989),
.B(n_1661),
.Y(n_1992)
);

CKINVDCx20_ASAP7_75t_R g1993 ( 
.A(n_1992),
.Y(n_1993)
);

AOI221xp5_ASAP7_75t_L g1994 ( 
.A1(n_1993),
.A2(n_1650),
.B1(n_1647),
.B2(n_1649),
.C(n_1639),
.Y(n_1994)
);

AOI211xp5_ASAP7_75t_L g1995 ( 
.A1(n_1994),
.A2(n_1639),
.B(n_1650),
.C(n_1647),
.Y(n_1995)
);


endmodule