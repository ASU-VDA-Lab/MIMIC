module fake_jpeg_2757_n_247 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_42),
.Y(n_113)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_2),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_58),
.Y(n_91)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_22),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_37),
.B1(n_36),
.B2(n_11),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_4),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_62),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_25),
.A2(n_6),
.B(n_7),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_57),
.B(n_30),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_23),
.B(n_33),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_21),
.A2(n_14),
.B1(n_15),
.B2(n_9),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_61),
.B1(n_69),
.B2(n_28),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_21),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_70),
.Y(n_96)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_76),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_17),
.A2(n_8),
.B1(n_11),
.B2(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_77),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_18),
.B(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_75),
.Y(n_102)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_11),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_20),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_63),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_32),
.B1(n_38),
.B2(n_26),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_80),
.A2(n_101),
.B1(n_109),
.B2(n_81),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_84),
.A2(n_114),
.B1(n_100),
.B2(n_82),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_37),
.B1(n_26),
.B2(n_28),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_89),
.A2(n_111),
.B(n_107),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_97),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_53),
.Y(n_97)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_30),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_35),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_116),
.Y(n_136)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_55),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_68),
.A2(n_19),
.B1(n_40),
.B2(n_56),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_79),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_51),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_118),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_44),
.B(n_66),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_91),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_122),
.B(n_125),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_124),
.A2(n_139),
.B1(n_142),
.B2(n_150),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_96),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_141),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_98),
.Y(n_130)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_130),
.B(n_152),
.CI(n_151),
.CON(n_165),
.SN(n_165)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_85),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_140),
.Y(n_161)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_87),
.B(n_113),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_82),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_84),
.A2(n_93),
.B1(n_110),
.B2(n_90),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_143),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_114),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_140),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_149),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_114),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_143),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_93),
.A2(n_110),
.B1(n_90),
.B2(n_100),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_151),
.Y(n_158)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_99),
.A2(n_89),
.B1(n_101),
.B2(n_104),
.Y(n_150)
);

OR2x4_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_95),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_154),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_104),
.A2(n_70),
.B1(n_75),
.B2(n_78),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_135),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_163),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_136),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_177),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_169),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_166),
.B(n_174),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_123),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_171),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_120),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_121),
.B(n_130),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_132),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_134),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_194),
.Y(n_204)
);

NAND2xp33_ASAP7_75t_SL g183 ( 
.A(n_155),
.B(n_142),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_192),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_197),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_129),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_186),
.B(n_191),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_129),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_193),
.C(n_196),
.Y(n_200)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_127),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_127),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_167),
.B1(n_161),
.B2(n_170),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_149),
.C(n_138),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_166),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_157),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_201),
.C(n_188),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_161),
.C(n_157),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_182),
.A2(n_172),
.B1(n_158),
.B2(n_176),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_208),
.Y(n_212)
);

A2O1A1O1Ixp25_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_165),
.B(n_177),
.C(n_160),
.D(n_158),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_185),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_158),
.B(n_164),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_194),
.A2(n_188),
.B1(n_181),
.B2(n_195),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_184),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_214),
.C(n_221),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_196),
.C(n_179),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_217),
.Y(n_223)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_183),
.B1(n_190),
.B2(n_189),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_220),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_185),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_218),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_219),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_165),
.C(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_228),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_212),
.A2(n_206),
.B(n_209),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_225),
.A2(n_204),
.B(n_209),
.Y(n_231)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_227),
.B1(n_209),
.B2(n_211),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_221),
.C(n_213),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_232),
.B(n_233),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_211),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_198),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_235),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_225),
.B(n_201),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_SL g236 ( 
.A(n_230),
.B(n_227),
.C(n_224),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_238),
.B(n_237),
.Y(n_242)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_230),
.A2(n_226),
.B(n_204),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_240),
.A2(n_205),
.B1(n_222),
.B2(n_202),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_241),
.A2(n_243),
.B(n_203),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_242),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_192),
.A3(n_203),
.B1(n_159),
.B2(n_160),
.C1(n_171),
.C2(n_173),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_239),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_245),
.Y(n_247)
);


endmodule