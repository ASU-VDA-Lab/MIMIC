module fake_jpeg_22094_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_SL g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_17),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_33),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_3),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_19),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_1),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_44),
.B1(n_23),
.B2(n_31),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_26),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_50),
.B(n_58),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_24),
.B(n_28),
.Y(n_50)
);

OR2x2_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_16),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_15),
.B(n_14),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_57),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_23),
.B1(n_27),
.B2(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_55),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_32),
.A2(n_33),
.B1(n_40),
.B2(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_20),
.B1(n_18),
.B2(n_27),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_62),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_33),
.A2(n_20),
.B1(n_21),
.B2(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_26),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_25),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_15),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_78),
.B(n_82),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_4),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_6),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_7),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_22),
.B(n_44),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_91),
.B(n_47),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_7),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_22),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_68),
.Y(n_110)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_10),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_92),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_47),
.A2(n_22),
.B(n_14),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_10),
.Y(n_92)
);

CKINVDCx10_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_100),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_55),
.C(n_69),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_102),
.C(n_83),
.Y(n_122)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_104),
.B(n_107),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_85),
.C(n_91),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_110),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_71),
.A2(n_63),
.B(n_45),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_68),
.B(n_22),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_75),
.B1(n_70),
.B2(n_79),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_116),
.B1(n_118),
.B2(n_98),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_75),
.B1(n_70),
.B2(n_56),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_88),
.B1(n_72),
.B2(n_87),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_118),
.B1(n_125),
.B2(n_122),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_72),
.B1(n_84),
.B2(n_77),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_72),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_122),
.C(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_121),
.A2(n_100),
.B1(n_105),
.B2(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_76),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_86),
.C(n_89),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_74),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_94),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_128),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_129),
.B(n_131),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_98),
.B(n_97),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_135),
.Y(n_138)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_94),
.B(n_86),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_137),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_117),
.B1(n_113),
.B2(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

OAI322xp33_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_112),
.A3(n_96),
.B1(n_106),
.B2(n_99),
.C1(n_111),
.C2(n_22),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_131),
.C(n_130),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_133),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_138),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_149),
.C(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

OAI21x1_ASAP7_75t_SL g154 ( 
.A1(n_151),
.A2(n_146),
.B(n_140),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_139),
.C(n_142),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_SL g160 ( 
.A1(n_154),
.A2(n_96),
.B(n_152),
.C(n_99),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_133),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_156),
.C(n_157),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_148),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_160),
.C(n_11),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_157),
.C(n_11),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.C(n_13),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_13),
.Y(n_164)
);


endmodule