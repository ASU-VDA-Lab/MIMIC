module fake_jpeg_2105_n_483 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_483);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_483;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_48),
.B(n_74),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g141 ( 
.A(n_50),
.Y(n_141)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_52),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_53),
.Y(n_134)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_56),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_61),
.Y(n_149)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g110 ( 
.A(n_65),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_82),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_72),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_27),
.B(n_14),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_36),
.B(n_7),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_84),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_41),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g144 ( 
.A(n_77),
.Y(n_144)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_43),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_18),
.B(n_8),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_37),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_97),
.Y(n_103)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_91),
.Y(n_133)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_18),
.B(n_8),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_96),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_37),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_37),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_72),
.A2(n_32),
.B1(n_46),
.B2(n_40),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_107),
.A2(n_117),
.B1(n_127),
.B2(n_143),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_53),
.B1(n_56),
.B2(n_59),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_109),
.A2(n_123),
.B1(n_128),
.B2(n_152),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_32),
.B1(n_46),
.B2(n_40),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_64),
.A2(n_32),
.B1(n_46),
.B2(n_29),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_61),
.A2(n_40),
.B1(n_45),
.B2(n_19),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_83),
.A2(n_29),
.B1(n_39),
.B2(n_26),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_76),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_63),
.A2(n_19),
.B1(n_45),
.B2(n_26),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_146),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_65),
.B(n_39),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_147),
.B(n_150),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_97),
.A2(n_31),
.B1(n_30),
.B2(n_42),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_57),
.B(n_42),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_66),
.A2(n_30),
.B1(n_31),
.B2(n_37),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_79),
.A2(n_47),
.B1(n_33),
.B2(n_28),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_158),
.Y(n_217)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_174),
.Y(n_215)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_161),
.Y(n_236)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_33),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_164),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_28),
.Y(n_164)
);

OR2x4_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_98),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_166),
.Y(n_238)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_100),
.B(n_87),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

INVx4_ASAP7_75t_SL g170 ( 
.A(n_110),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_125),
.A2(n_47),
.A3(n_96),
.B1(n_99),
.B2(n_89),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_171),
.A2(n_114),
.B(n_135),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_108),
.B(n_95),
.C(n_86),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_107),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_85),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_142),
.B(n_80),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_175),
.B(n_181),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_194),
.Y(n_214)
);

OR2x2_ASAP7_75t_SL g177 ( 
.A(n_112),
.B(n_49),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_177),
.Y(n_233)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_101),
.Y(n_178)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_118),
.B(n_0),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_183),
.Y(n_219)
);

INVx6_ASAP7_75t_SL g180 ( 
.A(n_101),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_180),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_133),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_0),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_124),
.B(n_73),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_190),
.Y(n_227)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_103),
.B(n_0),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_SL g207 ( 
.A(n_191),
.B(n_198),
.Y(n_207)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_193),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_68),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_197),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_0),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_203),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_114),
.B(n_9),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_200),
.B(n_202),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_122),
.A2(n_16),
.B1(n_20),
.B2(n_10),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_117),
.B1(n_153),
.B2(n_106),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_115),
.B(n_10),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_143),
.B(n_2),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_165),
.A2(n_127),
.B(n_148),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_206),
.A2(n_105),
.B(n_177),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_209),
.B(n_196),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_213),
.A2(n_223),
.B1(n_237),
.B2(n_198),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_228),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_160),
.A2(n_155),
.B1(n_130),
.B2(n_140),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_163),
.B(n_155),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_224),
.B(n_198),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_113),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_160),
.A2(n_130),
.B1(n_140),
.B2(n_119),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_239),
.Y(n_294)
);

BUFx12_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_184),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_241),
.B(n_261),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_242),
.B(n_260),
.Y(n_272)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_164),
.C(n_191),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_214),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_183),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_262),
.Y(n_271)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_219),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_257),
.C(n_233),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_226),
.A2(n_165),
.B1(n_195),
.B2(n_203),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_252),
.A2(n_253),
.B1(n_265),
.B2(n_267),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_226),
.A2(n_195),
.B1(n_176),
.B2(n_185),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_210),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_258),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_256),
.B(n_263),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_207),
.B(n_191),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_230),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_205),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_228),
.B(n_176),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_231),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_171),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_170),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_264),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_238),
.A2(n_195),
.B1(n_196),
.B2(n_166),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_205),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_266),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_268),
.A2(n_180),
.B(n_232),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_276),
.C(n_277),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_221),
.B1(n_237),
.B2(n_209),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_273),
.A2(n_274),
.B1(n_279),
.B2(n_280),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_221),
.B1(n_206),
.B2(n_233),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_214),
.C(n_172),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_214),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_285),
.C(n_291),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_248),
.A2(n_223),
.B1(n_227),
.B2(n_215),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_248),
.A2(n_263),
.B1(n_268),
.B2(n_258),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_227),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_261),
.A2(n_213),
.B1(n_215),
.B2(n_230),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_290),
.A2(n_296),
.B1(n_239),
.B2(n_216),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_244),
.B(n_249),
.C(n_245),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_242),
.B(n_222),
.C(n_204),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_276),
.C(n_278),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_252),
.A2(n_222),
.B1(n_231),
.B2(n_232),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_298),
.A2(n_158),
.B(n_168),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_243),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_300),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_266),
.Y(n_300)
);

AOI21xp33_ASAP7_75t_L g301 ( 
.A1(n_280),
.A2(n_253),
.B(n_246),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_301),
.A2(n_327),
.B(n_272),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_305),
.B(n_182),
.Y(n_352)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_283),
.B(n_265),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_313),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_218),
.C(n_260),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_269),
.C(n_277),
.Y(n_332)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_281),
.Y(n_309)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_240),
.B(n_250),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_288),
.Y(n_311)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_284),
.A2(n_262),
.B1(n_220),
.B2(n_240),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_324),
.B1(n_294),
.B2(n_286),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_259),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_271),
.B(n_247),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_315),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_218),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_295),
.B(n_240),
.Y(n_316)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_316),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_279),
.B(n_239),
.Y(n_317)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_317),
.Y(n_356)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_289),
.B(n_272),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_320),
.B(n_291),
.Y(n_334)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_292),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_321),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_322),
.A2(n_296),
.B1(n_286),
.B2(n_287),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_274),
.A2(n_212),
.B(n_229),
.C(n_220),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_L g339 ( 
.A1(n_323),
.A2(n_297),
.B(n_292),
.C(n_294),
.Y(n_339)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_270),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_287),
.B(n_229),
.Y(n_325)
);

XNOR2x2_ASAP7_75t_SL g333 ( 
.A(n_325),
.B(n_285),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_284),
.A2(n_234),
.B(n_105),
.Y(n_326)
);

OA21x2_ASAP7_75t_L g337 ( 
.A1(n_326),
.A2(n_273),
.B(n_290),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_297),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_328),
.A2(n_337),
.B(n_316),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_329),
.A2(n_348),
.B1(n_312),
.B2(n_356),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_338),
.C(n_344),
.Y(n_359)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_334),
.B(n_315),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_282),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_335),
.B(n_345),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_293),
.Y(n_338)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_339),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_341),
.A2(n_326),
.B1(n_327),
.B2(n_322),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_167),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_302),
.B(n_162),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_216),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_349),
.C(n_353),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_302),
.B(n_234),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_352),
.B(n_305),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_305),
.B(n_113),
.C(n_197),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_317),
.A2(n_186),
.B1(n_137),
.B2(n_136),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_354),
.A2(n_355),
.B1(n_188),
.B2(n_324),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_322),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_358),
.A2(n_366),
.B1(n_374),
.B2(n_381),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_335),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_343),
.A2(n_310),
.B(n_301),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_362),
.A2(n_368),
.B(n_369),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_336),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_378),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_345),
.B(n_320),
.Y(n_364)
);

NAND3xp33_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_370),
.C(n_372),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_365),
.A2(n_341),
.B1(n_355),
.B2(n_354),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_337),
.A2(n_303),
.B1(n_307),
.B2(n_312),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_343),
.A2(n_319),
.B(n_303),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_300),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_350),
.A2(n_303),
.B(n_323),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_373),
.A2(n_379),
.B(n_382),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_337),
.A2(n_299),
.B1(n_314),
.B2(n_313),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_308),
.C(n_321),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_352),
.C(n_353),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_351),
.B(n_311),
.Y(n_377)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_377),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_350),
.A2(n_323),
.B(n_308),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_330),
.B(n_325),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_383),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_329),
.A2(n_318),
.B1(n_309),
.B2(n_306),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_339),
.A2(n_324),
.B1(n_192),
.B2(n_187),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_336),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_344),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_388),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_386),
.B(n_397),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_387),
.A2(n_366),
.B1(n_358),
.B2(n_374),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_347),
.C(n_332),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_390),
.B(n_380),
.Y(n_422)
);

INVxp33_ASAP7_75t_SL g391 ( 
.A(n_377),
.Y(n_391)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_391),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_368),
.A2(n_333),
.B(n_346),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_392),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_362),
.A2(n_338),
.B(n_342),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_393),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_375),
.B(n_357),
.Y(n_394)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_394),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_369),
.A2(n_331),
.B(n_178),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_396),
.A2(n_404),
.B(n_383),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_236),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_359),
.B(n_151),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_401),
.B(n_386),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_236),
.C(n_119),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_405),
.C(n_360),
.Y(n_413)
);

O2A1O1Ixp33_ASAP7_75t_L g404 ( 
.A1(n_376),
.A2(n_236),
.B(n_161),
.C(n_154),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_361),
.B(n_236),
.C(n_154),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_406),
.A2(n_416),
.B1(n_399),
.B2(n_396),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_410),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_367),
.Y(n_411)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_411),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_371),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_413),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_379),
.C(n_373),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_414),
.B(n_421),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_365),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_418),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_400),
.A2(n_381),
.B1(n_367),
.B2(n_376),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_382),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_419),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_399),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_138),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_390),
.B(n_363),
.C(n_378),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_423),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_426),
.A2(n_156),
.B1(n_106),
.B2(n_141),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_424),
.A2(n_384),
.B(n_389),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_427),
.A2(n_437),
.B(n_439),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_389),
.C(n_384),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_429),
.B(n_430),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_395),
.C(n_402),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_402),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_433),
.B(n_435),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_423),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_395),
.C(n_387),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_SL g443 ( 
.A(n_436),
.B(n_422),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_404),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_417),
.B(n_151),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_16),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_425),
.A2(n_418),
.B(n_406),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_442),
.A2(n_452),
.B(n_438),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_444),
.Y(n_466)
);

INVx11_ASAP7_75t_L g444 ( 
.A(n_430),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_431),
.A2(n_419),
.B1(n_414),
.B2(n_420),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_445),
.B(n_449),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_441),
.A2(n_413),
.B(n_156),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_448),
.A2(n_16),
.B(n_20),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_10),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_451),
.B(n_453),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_429),
.A2(n_16),
.B(n_20),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_10),
.Y(n_453)
);

BUFx24_ASAP7_75t_SL g454 ( 
.A(n_434),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_454),
.B(n_440),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_455),
.B(n_438),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_458),
.Y(n_470)
);

AO21x1_ASAP7_75t_L g467 ( 
.A1(n_457),
.A2(n_460),
.B(n_461),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_434),
.C(n_436),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_459),
.B(n_462),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_16),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_8),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_442),
.A2(n_14),
.B(n_13),
.Y(n_465)
);

NAND3xp33_ASAP7_75t_SL g473 ( 
.A(n_465),
.B(n_11),
.C(n_3),
.Y(n_473)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_466),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_469),
.Y(n_476)
);

A2O1A1O1Ixp25_ASAP7_75t_L g471 ( 
.A1(n_458),
.A2(n_444),
.B(n_449),
.C(n_455),
.D(n_20),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_471),
.A2(n_472),
.B(n_463),
.Y(n_475)
);

A2O1A1Ixp33_ASAP7_75t_L g472 ( 
.A1(n_464),
.A2(n_13),
.B(n_11),
.C(n_20),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_473),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_470),
.A2(n_465),
.B(n_456),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_474),
.A2(n_475),
.B(n_11),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_477),
.B(n_468),
.C(n_467),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_478),
.B(n_479),
.C(n_480),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_476),
.A2(n_2),
.B(n_4),
.Y(n_480)
);

AOI221xp5_ASAP7_75t_L g482 ( 
.A1(n_481),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_469),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_482),
.B(n_5),
.Y(n_483)
);


endmodule