module fake_jpeg_16869_n_297 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_9),
.B(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_15),
.Y(n_107)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_0),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_24),
.B(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_32),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_56),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_23),
.B(n_9),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_62),
.Y(n_98)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_20),
.B(n_9),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_68),
.B(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_79),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_16),
.B(n_38),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_73),
.A2(n_100),
.B(n_66),
.C(n_106),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_77),
.B(n_78),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_27),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_41),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_89),
.B1(n_16),
.B2(n_50),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_88),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_22),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_97),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_19),
.B1(n_18),
.B2(n_28),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_12),
.B1(n_7),
.B2(n_10),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_37),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_19),
.B1(n_27),
.B2(n_36),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_36),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_92),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_25),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_20),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_1),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_98),
.B(n_66),
.C(n_97),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_104),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_25),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_103),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_23),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_26),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_26),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_16),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_108),
.A2(n_148),
.B(n_93),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_78),
.A2(n_45),
.B1(n_46),
.B2(n_44),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_109),
.A2(n_121),
.B1(n_142),
.B2(n_105),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_110),
.B(n_125),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_50),
.B1(n_2),
.B2(n_3),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_111),
.A2(n_134),
.B1(n_141),
.B2(n_105),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_122),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_70),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_115),
.A2(n_120),
.B1(n_124),
.B2(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_77),
.B(n_58),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_133),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_63),
.B1(n_17),
.B2(n_1),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_82),
.A2(n_17),
.B1(n_3),
.B2(n_5),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_69),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_131),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_70),
.A2(n_17),
.B1(n_6),
.B2(n_7),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_84),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_145),
.B(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_101),
.B(n_63),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_68),
.A2(n_1),
.B1(n_11),
.B2(n_14),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_75),
.B1(n_94),
.B2(n_99),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_82),
.A2(n_72),
.B1(n_67),
.B2(n_98),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_134),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_74),
.A2(n_65),
.B1(n_96),
.B2(n_76),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_146),
.B(n_107),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_114),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_153),
.B(n_161),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_83),
.C(n_93),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_151),
.C(n_171),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_164),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_83),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_167),
.Y(n_186)
);

NOR4xp25_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_110),
.C(n_120),
.D(n_128),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_114),
.B(n_74),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_176),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_126),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_138),
.B1(n_147),
.B2(n_123),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g166 ( 
.A(n_108),
.B(n_76),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_170),
.B(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_130),
.B(n_96),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_65),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_178),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_111),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_116),
.B(n_112),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_174),
.C(n_122),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_112),
.B(n_119),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_109),
.B(n_148),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_151),
.B(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_117),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_125),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_132),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_137),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_181),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_117),
.B(n_131),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_135),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_180),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_188),
.B(n_192),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_146),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_206),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_190),
.A2(n_208),
.B(n_197),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_198),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_147),
.B1(n_172),
.B2(n_165),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_150),
.A2(n_162),
.B1(n_177),
.B2(n_175),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_166),
.B1(n_155),
.B2(n_157),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_170),
.A2(n_158),
.B1(n_176),
.B2(n_159),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_200),
.B1(n_210),
.B2(n_214),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_159),
.A2(n_164),
.B1(n_183),
.B2(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_156),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_213),
.B1(n_211),
.B2(n_197),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_184),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_149),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_208),
.C(n_199),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_171),
.A2(n_180),
.B1(n_182),
.B2(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_175),
.B1(n_172),
.B2(n_165),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_152),
.A2(n_175),
.B1(n_172),
.B2(n_165),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_202),
.B1(n_196),
.B2(n_209),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_185),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_216),
.B(n_226),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_160),
.Y(n_218)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_193),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_227),
.C(n_238),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_207),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_215),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_SL g241 ( 
.A1(n_228),
.A2(n_194),
.B(n_200),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_188),
.B(n_206),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_210),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_191),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_220),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_232),
.B(n_235),
.Y(n_242)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_236),
.B1(n_202),
.B2(n_212),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_214),
.B(n_195),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_250),
.B1(n_252),
.B2(n_230),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_243),
.B(n_245),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_255),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_220),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_221),
.A2(n_192),
.B1(n_236),
.B2(n_232),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_221),
.A2(n_238),
.B1(n_235),
.B2(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_223),
.C(n_218),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_256),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_217),
.C(n_229),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_226),
.Y(n_259)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_259),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_230),
.Y(n_260)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_223),
.Y(n_262)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_239),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_239),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_258),
.A2(n_257),
.B1(n_252),
.B2(n_250),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_259),
.B1(n_269),
.B2(n_260),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_234),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_265),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_242),
.B(n_248),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_274),
.B(n_271),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_242),
.C(n_244),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_251),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_279),
.B(n_281),
.Y(n_290)
);

FAx1_ASAP7_75t_SL g280 ( 
.A(n_274),
.B(n_263),
.CI(n_267),
.CON(n_280),
.SN(n_280)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_265),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_256),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_266),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_272),
.C(n_275),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_277),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_288),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_289),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_280),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_279),
.B1(n_276),
.B2(n_282),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_288),
.C(n_286),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_295),
.C(n_292),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_287),
.Y(n_297)
);


endmodule