module fake_jpeg_7625_n_122 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_122);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx8_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_19),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_39),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_13),
.B1(n_19),
.B2(n_25),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_13),
.B1(n_25),
.B2(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_15),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_20),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_61),
.B(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_22),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_38),
.B1(n_25),
.B2(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_66),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_71),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_40),
.C(n_38),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_61),
.Y(n_77)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_0),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_57),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_80),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_84),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_36),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_84),
.C(n_85),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_65),
.B1(n_74),
.B2(n_62),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_95),
.B1(n_73),
.B2(n_18),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_52),
.B(n_62),
.C(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_94),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_47),
.B1(n_64),
.B2(n_66),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_12),
.B(n_17),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_102),
.B1(n_91),
.B2(n_14),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_22),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_18),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_106),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_101),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_87),
.B1(n_86),
.B2(n_17),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_98),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_14),
.C(n_12),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_12),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_9),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_114),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_105),
.B1(n_106),
.B2(n_109),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_117),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_9),
.B1(n_11),
.B2(n_3),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_2),
.B(n_3),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_4),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_4),
.Y(n_122)
);


endmodule