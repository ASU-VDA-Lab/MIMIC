module fake_jpeg_18157_n_255 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_255);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_6),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_11),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_19),
.B1(n_14),
.B2(n_18),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_33),
.B1(n_27),
.B2(n_22),
.Y(n_49)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_52),
.B1(n_59),
.B2(n_36),
.Y(n_75)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_31),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_25),
.C(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_50),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_41),
.B1(n_36),
.B2(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_56),
.Y(n_65)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_53),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_58),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_19),
.B1(n_27),
.B2(n_35),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_38),
.B1(n_36),
.B2(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_29),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_78),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_63),
.A2(n_67),
.B1(n_74),
.B2(n_45),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_66),
.B1(n_49),
.B2(n_45),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_19),
.B1(n_33),
.B2(n_43),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_25),
.B1(n_33),
.B2(n_19),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_53),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_74)
);

CKINVDCx10_ASAP7_75t_R g95 ( 
.A(n_75),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_28),
.C(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_87),
.Y(n_101)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_79),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_47),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_91),
.Y(n_104)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_48),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_57),
.C(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_58),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_67),
.B1(n_96),
.B2(n_83),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_63),
.B1(n_64),
.B2(n_88),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_99),
.B1(n_44),
.B2(n_61),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_79),
.B(n_74),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_106),
.B(n_111),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_81),
.B1(n_68),
.B2(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_16),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_55),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_37),
.Y(n_133)
);

NAND2x1_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_74),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_77),
.B(n_74),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_112),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_12),
.B(n_60),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_113),
.A2(n_86),
.B1(n_21),
.B2(n_72),
.Y(n_117)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_116),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g115 ( 
.A(n_80),
.B(n_28),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_34),
.Y(n_140)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_126),
.C(n_138),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_119),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_61),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_127),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_29),
.B(n_12),
.C(n_21),
.Y(n_123)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_139),
.Y(n_143)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

OAI211xp5_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_28),
.B(n_26),
.C(n_15),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_26),
.C(n_37),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_133),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_70),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_70),
.Y(n_132)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_133),
.B(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_20),
.Y(n_137)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_37),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_15),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_115),
.B(n_114),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_150),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_101),
.Y(n_145)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_138),
.B1(n_113),
.B2(n_140),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_146),
.A2(n_117),
.B1(n_22),
.B2(n_18),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_20),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_97),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_108),
.B(n_98),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_152),
.A2(n_22),
.B(n_59),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_140),
.B(n_118),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_97),
.B1(n_44),
.B2(n_52),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_161),
.B1(n_59),
.B2(n_14),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_120),
.Y(n_155)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_119),
.A2(n_44),
.B1(n_52),
.B2(n_18),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_15),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_15),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_15),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_121),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_125),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_160),
.B(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_165),
.B(n_175),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_123),
.C(n_126),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_162),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_171),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_148),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_174),
.A2(n_182),
.B(n_184),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_157),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_176),
.B(n_9),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_10),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_143),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_14),
.B1(n_10),
.B2(n_9),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_181),
.B1(n_161),
.B2(n_154),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_14),
.B1(n_15),
.B2(n_9),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_34),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_194),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_192),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_188),
.A2(n_195),
.B1(n_184),
.B2(n_13),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_150),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_197),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_146),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_151),
.B1(n_159),
.B2(n_142),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_178),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_153),
.C(n_156),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_170),
.C(n_182),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_200),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_185),
.C(n_34),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_191),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_204),
.B(n_208),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_169),
.B1(n_177),
.B2(n_180),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_211),
.B1(n_185),
.B2(n_1),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_182),
.C(n_156),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_168),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_213),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_7),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_7),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_205),
.A2(n_194),
.B(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_206),
.A2(n_208),
.B(n_201),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_223),
.B(n_203),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_216),
.B(n_0),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_221),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_17),
.C(n_23),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_203),
.B1(n_8),
.B2(n_2),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_1),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_20),
.Y(n_223)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_225),
.Y(n_234)
);

INVx11_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_231),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_228),
.B(n_229),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_221),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_219),
.B1(n_224),
.B2(n_223),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_233),
.B(n_3),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_238),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_16),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_240),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_229),
.C(n_230),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_16),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_237),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_236),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_246),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_245),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_243),
.A3(n_242),
.B1(n_234),
.B2(n_23),
.C1(n_17),
.C2(n_5),
.Y(n_249)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_250),
.B(n_3),
.Y(n_251)
);

AOI322xp5_ASAP7_75t_L g250 ( 
.A1(n_247),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_17),
.C1(n_23),
.C2(n_245),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_251),
.A2(n_3),
.B(n_4),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_252),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_4),
.B(n_5),
.C(n_17),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_254),
.A2(n_17),
.B(n_216),
.Y(n_255)
);


endmodule