module fake_jpeg_20379_n_255 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_42),
.B(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_21),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_53),
.C(n_42),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_30),
.B1(n_19),
.B2(n_23),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_58),
.B1(n_32),
.B2(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_21),
.Y(n_53)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_30),
.B1(n_25),
.B2(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_69),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_30),
.B1(n_28),
.B2(n_25),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_109)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_19),
.B1(n_23),
.B2(n_26),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_41),
.B1(n_42),
.B2(n_37),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_46),
.B1(n_55),
.B2(n_47),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_24),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_19),
.B1(n_23),
.B2(n_26),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_72),
.A2(n_79),
.B1(n_20),
.B2(n_1),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_22),
.B(n_20),
.C(n_37),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_42),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_40),
.B(n_39),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_24),
.B1(n_27),
.B2(n_18),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_18),
.B1(n_31),
.B2(n_21),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_82),
.B1(n_88),
.B2(n_37),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_46),
.B1(n_54),
.B2(n_21),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_86),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_18),
.B1(n_31),
.B2(n_21),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_22),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_31),
.B1(n_22),
.B2(n_20),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_107),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_102),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_64),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_113),
.B1(n_69),
.B2(n_75),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_67),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_61),
.A2(n_22),
.B1(n_20),
.B2(n_2),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_40),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_39),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_134),
.B(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_80),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_66),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_72),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_131),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_63),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_75),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_128),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_138),
.B1(n_115),
.B2(n_99),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_68),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_68),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_140),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_68),
.B1(n_67),
.B2(n_86),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_135),
.B1(n_102),
.B2(n_107),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_71),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_92),
.A2(n_67),
.B(n_81),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_81),
.B1(n_85),
.B2(n_65),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_90),
.B(n_16),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_137),
.B(n_14),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_85),
.B1(n_84),
.B2(n_2),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_87),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_142),
.B(n_0),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_163),
.B(n_166),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_147),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_103),
.B1(n_114),
.B2(n_90),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_146),
.A2(n_155),
.B(n_162),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_122),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_151),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_128),
.B1(n_120),
.B2(n_134),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_114),
.Y(n_152)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_101),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_127),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_108),
.B1(n_3),
.B2(n_4),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_101),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_97),
.B(n_99),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_165),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_135),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_118),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_177),
.B1(n_159),
.B2(n_167),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_142),
.C(n_116),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_153),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_116),
.C(n_117),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_186),
.C(n_161),
.Y(n_191)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_121),
.C(n_15),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_185),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_158),
.A2(n_141),
.B1(n_138),
.B2(n_130),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_178),
.B(n_184),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_141),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_108),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_115),
.B(n_1),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_108),
.C(n_15),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_188),
.A2(n_164),
.B1(n_153),
.B2(n_160),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_195),
.B1(n_203),
.B2(n_205),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_196),
.Y(n_218)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_151),
.C(n_162),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_198),
.C(n_178),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_156),
.B1(n_148),
.B2(n_158),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_149),
.C(n_162),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_150),
.C(n_146),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_182),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_189),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_160),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_166),
.B1(n_165),
.B2(n_164),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_180),
.B(n_145),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_206),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_194),
.B(n_170),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_186),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_209),
.B(n_213),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_175),
.B(n_183),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_211),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_184),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_215),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_199),
.A2(n_181),
.B(n_185),
.Y(n_213)
);

OAI21x1_ASAP7_75t_L g216 ( 
.A1(n_204),
.A2(n_172),
.B(n_171),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_197),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_219),
.B(n_200),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_201),
.B1(n_197),
.B2(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_224),
.C(n_229),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_226),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_200),
.C(n_3),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_0),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_227),
.A2(n_230),
.B(n_7),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_4),
.C(n_5),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_6),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_231),
.B(n_232),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_208),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_213),
.B(n_210),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_237),
.B(n_225),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_218),
.C(n_208),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_238),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_7),
.B(n_8),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_230),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_240),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_229),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_224),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_241),
.B(n_242),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_8),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_240),
.A2(n_238),
.B(n_10),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_10),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_9),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_244),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g252 ( 
.A(n_249),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_SL g253 ( 
.A(n_250),
.B(n_251),
.C(n_248),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_11),
.B(n_12),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_252),
.Y(n_255)
);


endmodule