module real_jpeg_18515_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_290;
wire n_239;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_0),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_0),
.A2(n_56),
.B1(n_430),
.B2(n_433),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_0),
.A2(n_56),
.B1(n_532),
.B2(n_535),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_2),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_3),
.A2(n_125),
.B1(n_129),
.B2(n_130),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_3),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_3),
.A2(n_129),
.B1(n_277),
.B2(n_283),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_3),
.A2(n_129),
.B1(n_340),
.B2(n_345),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_3),
.A2(n_63),
.B1(n_129),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_4),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_4),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_4),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_4),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_5),
.A2(n_192),
.B1(n_193),
.B2(n_197),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_5),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_5),
.A2(n_192),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_5),
.A2(n_192),
.B1(n_395),
.B2(n_400),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_5),
.A2(n_175),
.B1(n_192),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_6),
.B(n_152),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g245 ( 
.A1(n_6),
.A2(n_70),
.A3(n_99),
.B1(n_246),
.B2(n_249),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_6),
.B(n_123),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_6),
.A2(n_62),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_6),
.A2(n_28),
.B1(n_362),
.B2(n_369),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_7),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g374 ( 
.A(n_7),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_8),
.A2(n_423),
.B1(n_424),
.B2(n_425),
.Y(n_422)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_8),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_8),
.A2(n_236),
.B1(n_425),
.B2(n_440),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_L g181 ( 
.A1(n_9),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_9),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_9),
.A2(n_185),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_9),
.A2(n_185),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_9),
.A2(n_163),
.B1(n_185),
.B2(n_457),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_10),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_10),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_10),
.Y(n_214)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_10),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_10),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_10),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_11),
.A2(n_39),
.B1(n_413),
.B2(n_416),
.Y(n_412)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_11),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_SL g491 ( 
.A1(n_11),
.A2(n_416),
.B1(n_492),
.B2(n_495),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_12),
.Y(n_156)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_12),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_13),
.A2(n_115),
.B1(n_118),
.B2(n_122),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_13),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_13),
.A2(n_122),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_13),
.A2(n_122),
.B1(n_271),
.B2(n_275),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_13),
.A2(n_122),
.B1(n_359),
.B2(n_363),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_14),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g439 ( 
.A1(n_14),
.A2(n_43),
.B1(n_440),
.B2(n_441),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_14),
.A2(n_43),
.B1(n_509),
.B2(n_511),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_15),
.A2(n_140),
.B1(n_146),
.B2(n_147),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_15),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_15),
.A2(n_146),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_15),
.A2(n_146),
.B1(n_463),
.B2(n_466),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_15),
.A2(n_146),
.B1(n_551),
.B2(n_553),
.Y(n_550)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g208 ( 
.A(n_16),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_16),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

BUFx8_ASAP7_75t_L g164 ( 
.A(n_17),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_519),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_483),
.B(n_517),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_387),
.B(n_480),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_264),
.B(n_386),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_228),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_24),
.B(n_228),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_160),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_87),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_26),
.B(n_87),
.C(n_160),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_60),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_27),
.B(n_60),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_36),
.B1(n_48),
.B2(n_57),
.Y(n_27)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_28),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_28),
.A2(n_288),
.B1(n_291),
.B2(n_295),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_28),
.A2(n_339),
.B1(n_362),
.B2(n_372),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_28),
.A2(n_48),
.B1(n_412),
.B2(n_449),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_28),
.A2(n_422),
.B(n_499),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_29),
.A2(n_138),
.B1(n_139),
.B2(n_256),
.Y(n_255)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_32),
.Y(n_452)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_35),
.Y(n_205)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_35),
.Y(n_359)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_35),
.Y(n_415)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_37),
.A2(n_138),
.B1(n_139),
.B2(n_148),
.Y(n_137)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_38),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_41),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_42),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_54),
.Y(n_423)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_57),
.B(n_62),
.Y(n_360)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_58),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_59),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_67),
.B1(n_73),
.B2(n_80),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_61),
.A2(n_62),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_62),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_62),
.B(n_321),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_SL g331 ( 
.A1(n_62),
.A2(n_320),
.B(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_R g375 ( 
.A(n_62),
.B(n_227),
.Y(n_375)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_66),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_66),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_72),
.Y(n_308)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_72),
.Y(n_465)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_72),
.Y(n_539)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_77),
.Y(n_189)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_79),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OA21x2_ASAP7_75t_L g165 ( 
.A1(n_81),
.A2(n_153),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_83),
.Y(n_459)
);

INVx6_ASAP7_75t_L g552 ( 
.A(n_83),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_84),
.Y(n_178)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_137),
.C(n_151),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_88),
.B(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_113),
.B1(n_123),
.B2(n_124),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_89),
.A2(n_123),
.B1(n_124),
.B2(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_89),
.A2(n_123),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_90),
.A2(n_114),
.B1(n_304),
.B2(n_309),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_90),
.A2(n_309),
.B1(n_393),
.B2(n_394),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_90),
.A2(n_309),
.B1(n_394),
.B2(n_462),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_90),
.A2(n_309),
.B1(n_462),
.B2(n_508),
.Y(n_507)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_99),
.B(n_105),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22x1_ASAP7_75t_SL g153 ( 
.A1(n_97),
.A2(n_154),
.B1(n_157),
.B2(n_159),
.Y(n_153)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_106),
.B1(n_108),
.B2(n_110),
.Y(n_105)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_102),
.Y(n_534)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_103),
.Y(n_510)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_106),
.Y(n_221)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_106),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_107),
.Y(n_282)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_107),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_109),
.Y(n_248)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_109),
.Y(n_432)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_121),
.Y(n_184)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_123),
.Y(n_309)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_125),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_128),
.Y(n_514)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_137),
.B(n_151),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_138),
.A2(n_338),
.B1(n_348),
.B2(n_350),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_138),
.A2(n_411),
.B1(n_417),
.B2(n_421),
.Y(n_410)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_144),
.Y(n_289)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_145),
.Y(n_290)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_148),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_149),
.Y(n_349)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_150),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_152),
.A2(n_162),
.B1(n_165),
.B2(n_171),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_152),
.A2(n_165),
.B1(n_171),
.B2(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_152),
.Y(n_460)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_158),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_179),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_161),
.B(n_180),
.C(n_190),
.Y(n_474)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_164),
.Y(n_407)
);

INVx3_ASAP7_75t_SL g455 ( 
.A(n_165),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_178),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_178),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_190),
.Y(n_179)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_181),
.Y(n_393)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_200),
.B1(n_219),
.B2(n_226),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_195),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_196),
.Y(n_199)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_196),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_200),
.A2(n_226),
.B1(n_270),
.B2(n_276),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_200),
.A2(n_226),
.B1(n_235),
.B2(n_276),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_200),
.A2(n_226),
.B1(n_270),
.B2(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_200),
.B(n_438),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_200),
.A2(n_226),
.B1(n_541),
.B2(n_542),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_212),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_205),
.B1(n_206),
.B2(n_209),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_208),
.Y(n_347)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_214),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_217),
.Y(n_319)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_218),
.Y(n_440)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_220),
.A2(n_227),
.B1(n_233),
.B2(n_439),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_226),
.B(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_227),
.A2(n_233),
.B1(n_234),
.B2(n_242),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_227),
.A2(n_233),
.B1(n_429),
.B2(n_491),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.C(n_243),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_230),
.B(n_382),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_232),
.A2(n_243),
.B1(n_244),
.B2(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_232),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_254),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_245),
.A2(n_254),
.B1(n_255),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_256),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_380),
.B(n_385),
.Y(n_264)
);

AOI21x1_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_312),
.B(n_379),
.Y(n_265)
);

NAND2xp33_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_298),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_267),
.B(n_298),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_287),
.C(n_296),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_268),
.A2(n_269),
.B1(n_296),
.B2(n_297),
.Y(n_334)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_285),
.Y(n_332)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_287),
.B(n_334),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

OAI32xp33_ASAP7_75t_L g315 ( 
.A1(n_290),
.A2(n_316),
.A3(n_319),
.B1(n_320),
.B2(n_324),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_299),
.B(n_302),
.C(n_311),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_310),
.B2(n_311),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_335),
.B(n_378),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_333),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_314),
.B(n_333),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_329),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_315),
.A2(n_329),
.B1(n_330),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_318),
.Y(n_494)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx5_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_353),
.B(n_377),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_351),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_337),
.B(n_351),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_344),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_347),
.Y(n_424)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_370),
.B(n_376),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_361),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_360),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_375),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_371),
.B(n_375),
.Y(n_376)
);

INVx6_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx12f_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_384),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_389),
.A2(n_468),
.B(n_475),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_389),
.B(n_468),
.C(n_482),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_408),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_390),
.B(n_409),
.C(n_445),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_402),
.C(n_403),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_392),
.B(n_403),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_399),
.Y(n_401)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_402),
.B(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_405),
.A2(n_455),
.B1(n_456),
.B2(n_460),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_445),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_426),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_410),
.A2(n_427),
.B(n_437),
.Y(n_515)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_437),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_432),
.Y(n_436)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_453),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_446),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

XOR2x2_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_448),
.Y(n_472)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_451),
.Y(n_450)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_461),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_454),
.B(n_461),
.C(n_487),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_455),
.A2(n_456),
.B1(n_460),
.B2(n_504),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_455),
.A2(n_460),
.B1(n_504),
.B2(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx6_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_472),
.C(n_473),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_469),
.A2(n_470),
.B1(n_478),
.B2(n_479),
.Y(n_477)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_472),
.B(n_474),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_476),
.B(n_477),
.Y(n_482)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_478),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_485),
.B(n_516),
.Y(n_484)
);

NOR2xp67_ASAP7_75t_SL g518 ( 
.A(n_485),
.B(n_516),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_488),
.Y(n_485)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_486),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_501),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_489),
.B(n_522),
.C(n_523),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_490),
.A2(n_497),
.B1(n_498),
.B2(n_500),
.Y(n_489)
);

INVxp33_ASAP7_75t_SL g500 ( 
.A(n_490),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_490),
.B(n_498),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_491),
.Y(n_541)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_497),
.A2(n_498),
.B1(n_548),
.B2(n_549),
.Y(n_547)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_501),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_515),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_507),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_503),
.B(n_507),
.C(n_515),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_508),
.Y(n_529)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_556),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_524),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_521),
.B(n_524),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_526),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_544),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_528),
.A2(n_540),
.B(n_543),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_528),
.B(n_540),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_545),
.A2(n_546),
.B1(n_547),
.B2(n_555),
.Y(n_544)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_545),
.Y(n_555)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

INVx3_ASAP7_75t_SL g553 ( 
.A(n_554),
.Y(n_553)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);


endmodule