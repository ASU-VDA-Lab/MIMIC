module real_aes_2694_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_756;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_0), .B(n_128), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_1), .A2(n_31), .B1(n_104), .B2(n_105), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_1), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_2), .A2(n_122), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_3), .B(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_4), .B(n_128), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_5), .B(n_139), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_6), .B(n_139), .Y(n_214) );
INVx1_ASAP7_75t_L g127 ( .A(n_7), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_8), .B(n_139), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g740 ( .A(n_9), .Y(n_740) );
NAND2xp33_ASAP7_75t_L g190 ( .A(n_10), .B(n_137), .Y(n_190) );
AND2x2_ASAP7_75t_L g447 ( .A(n_11), .B(n_184), .Y(n_447) );
AND2x2_ASAP7_75t_L g455 ( .A(n_12), .B(n_151), .Y(n_455) );
INVx2_ASAP7_75t_L g119 ( .A(n_13), .Y(n_119) );
AOI221x1_ASAP7_75t_L g121 ( .A1(n_14), .A2(n_25), .B1(n_122), .B2(n_128), .C(n_135), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_15), .B(n_139), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g417 ( .A(n_16), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_17), .B(n_128), .Y(n_186) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_18), .A2(n_184), .B(n_185), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_19), .B(n_117), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_20), .B(n_139), .Y(n_198) );
AO21x1_ASAP7_75t_L g209 ( .A1(n_21), .A2(n_128), .B(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_22), .B(n_128), .Y(n_486) );
INVx1_ASAP7_75t_L g421 ( .A(n_23), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_24), .A2(n_89), .B1(n_128), .B2(n_516), .Y(n_515) );
NAND2x1_ASAP7_75t_L g147 ( .A(n_26), .B(n_139), .Y(n_147) );
NAND2x1_ASAP7_75t_L g177 ( .A(n_27), .B(n_137), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_28), .Y(n_755) );
OR2x2_ASAP7_75t_L g120 ( .A(n_29), .B(n_86), .Y(n_120) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_29), .A2(n_86), .B(n_119), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_30), .B(n_137), .Y(n_172) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_31), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_32), .B(n_139), .Y(n_189) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_33), .A2(n_151), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_34), .B(n_137), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_35), .A2(n_122), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_36), .B(n_139), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_37), .A2(n_122), .B(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g123 ( .A(n_38), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g134 ( .A(n_38), .B(n_127), .Y(n_134) );
INVx1_ASAP7_75t_L g524 ( .A(n_38), .Y(n_524) );
OR2x6_ASAP7_75t_L g419 ( .A(n_39), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_40), .B(n_128), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_41), .B(n_128), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_42), .B(n_139), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_43), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_44), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_45), .B(n_137), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_46), .B(n_128), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_47), .A2(n_122), .B(n_451), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_48), .A2(n_122), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_49), .B(n_137), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_50), .B(n_137), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_51), .B(n_128), .Y(n_460) );
INVx1_ASAP7_75t_L g126 ( .A(n_52), .Y(n_126) );
INVx1_ASAP7_75t_L g131 ( .A(n_52), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_53), .B(n_139), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_54), .A2(n_61), .B1(n_750), .B2(n_751), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_54), .Y(n_750) );
AND2x2_ASAP7_75t_L g477 ( .A(n_55), .B(n_117), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_56), .B(n_137), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_57), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_58), .B(n_137), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_59), .A2(n_122), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_60), .B(n_128), .Y(n_454) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_61), .A2(n_101), .B1(n_734), .B2(n_744), .C1(n_756), .C2(n_760), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_61), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_62), .B(n_128), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_63), .A2(n_122), .B(n_468), .Y(n_467) );
AO21x1_ASAP7_75t_L g211 ( .A1(n_64), .A2(n_122), .B(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g492 ( .A(n_65), .B(n_118), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_66), .B(n_128), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_67), .B(n_137), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_68), .B(n_128), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_69), .B(n_137), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_70), .A2(n_94), .B1(n_122), .B2(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g162 ( .A(n_71), .B(n_118), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_72), .B(n_139), .Y(n_489) );
INVx1_ASAP7_75t_L g124 ( .A(n_73), .Y(n_124) );
INVx1_ASAP7_75t_L g133 ( .A(n_73), .Y(n_133) );
AND2x2_ASAP7_75t_L g181 ( .A(n_74), .B(n_151), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_75), .B(n_137), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_76), .A2(n_122), .B(n_481), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_77), .A2(n_122), .B(n_434), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_78), .A2(n_122), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g472 ( .A(n_79), .B(n_118), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_80), .B(n_117), .Y(n_513) );
INVx1_ASAP7_75t_L g422 ( .A(n_81), .Y(n_422) );
AND2x2_ASAP7_75t_L g166 ( .A(n_82), .B(n_151), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_83), .B(n_128), .Y(n_200) );
AND2x2_ASAP7_75t_L g437 ( .A(n_84), .B(n_184), .Y(n_437) );
AND2x2_ASAP7_75t_L g210 ( .A(n_85), .B(n_191), .Y(n_210) );
AND2x2_ASAP7_75t_L g154 ( .A(n_87), .B(n_151), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_88), .B(n_137), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_90), .B(n_139), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_91), .B(n_137), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_92), .A2(n_122), .B(n_197), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_93), .A2(n_122), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_95), .B(n_139), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_96), .B(n_139), .Y(n_171) );
BUFx2_ASAP7_75t_L g491 ( .A(n_97), .Y(n_491) );
BUFx2_ASAP7_75t_L g741 ( .A(n_98), .Y(n_741) );
BUFx2_ASAP7_75t_SL g766 ( .A(n_98), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_99), .A2(n_122), .B(n_188), .Y(n_187) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AOI221xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_106), .B1(n_725), .B2(n_728), .C(n_729), .Y(n_102) );
INVx1_ASAP7_75t_L g728 ( .A(n_103), .Y(n_728) );
OAI22x1_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_414), .B1(n_423), .B2(n_723), .Y(n_106) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_108), .A2(n_416), .B1(n_424), .B2(n_726), .Y(n_725) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_326), .Y(n_108) );
AND4x1_ASAP7_75t_L g109 ( .A(n_110), .B(n_238), .C(n_265), .D(n_300), .Y(n_109) );
AOI221xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_163), .B1(n_203), .B2(n_218), .C(n_222), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_142), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_113), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OR2x2_ASAP7_75t_L g279 ( .A(n_114), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g334 ( .A(n_114), .B(n_289), .Y(n_334) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g237 ( .A(n_115), .B(n_155), .Y(n_237) );
AND2x4_ASAP7_75t_L g273 ( .A(n_115), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g287 ( .A(n_115), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g204 ( .A(n_116), .Y(n_204) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_116), .Y(n_376) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_141), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_117), .A2(n_168), .B(n_169), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_117), .Y(n_180) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_117), .A2(n_121), .B(n_141), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_117), .A2(n_432), .B(n_433), .Y(n_431) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_117), .A2(n_515), .B(n_521), .Y(n_514) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_SL g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x4_ASAP7_75t_L g191 ( .A(n_119), .B(n_120), .Y(n_191) );
AND2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
BUFx3_ASAP7_75t_L g520 ( .A(n_123), .Y(n_520) );
AND2x6_ASAP7_75t_L g137 ( .A(n_124), .B(n_130), .Y(n_137) );
INVx2_ASAP7_75t_L g526 ( .A(n_124), .Y(n_526) );
AND2x4_ASAP7_75t_L g522 ( .A(n_125), .B(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x4_ASAP7_75t_L g139 ( .A(n_126), .B(n_132), .Y(n_139) );
INVx2_ASAP7_75t_L g518 ( .A(n_126), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_127), .Y(n_519) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_134), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx5_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_138), .B(n_140), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_137), .B(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_140), .A2(n_147), .B(n_148), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_140), .A2(n_159), .B(n_160), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_140), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_140), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_140), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_140), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_140), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_140), .A2(n_435), .B(n_436), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_140), .A2(n_444), .B(n_445), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_140), .A2(n_452), .B(n_453), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_140), .A2(n_463), .B(n_464), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_140), .A2(n_469), .B(n_470), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_140), .A2(n_482), .B(n_483), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_140), .A2(n_489), .B(n_490), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_SL g231 ( .A1(n_142), .A2(n_204), .B(n_232), .C(n_236), .Y(n_231) );
AND2x2_ASAP7_75t_L g252 ( .A(n_142), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_142), .B(n_204), .Y(n_392) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_155), .Y(n_142) );
INVx2_ASAP7_75t_L g272 ( .A(n_143), .Y(n_272) );
BUFx3_ASAP7_75t_L g288 ( .A(n_143), .Y(n_288) );
INVxp67_ASAP7_75t_L g292 ( .A(n_143), .Y(n_292) );
AO21x2_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_150), .B(n_154), .Y(n_143) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_144), .A2(n_150), .B(n_154), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
AO21x2_ASAP7_75t_L g155 ( .A1(n_150), .A2(n_156), .B(n_162), .Y(n_155) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_150), .A2(n_156), .B(n_162), .Y(n_217) );
AO21x1_ASAP7_75t_SL g465 ( .A1(n_150), .A2(n_466), .B(n_472), .Y(n_465) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_150), .A2(n_466), .B(n_472), .Y(n_499) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_152), .A2(n_449), .B(n_455), .Y(n_448) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx4f_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
INVx2_ASAP7_75t_L g271 ( .A(n_155), .Y(n_271) );
AND2x2_ASAP7_75t_L g277 ( .A(n_155), .B(n_250), .Y(n_277) );
AND2x2_ASAP7_75t_L g303 ( .A(n_155), .B(n_272), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_157), .B(n_161), .Y(n_156) );
AOI211xp5_ASAP7_75t_L g300 ( .A1(n_163), .A2(n_301), .B(n_304), .C(n_314), .Y(n_300) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_164), .B(n_182), .Y(n_163) );
OAI321xp33_ASAP7_75t_L g275 ( .A1(n_164), .A2(n_223), .A3(n_276), .B1(n_278), .B2(n_279), .C(n_281), .Y(n_275) );
AND2x2_ASAP7_75t_L g396 ( .A(n_164), .B(n_371), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_164), .Y(n_399) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_173), .Y(n_164) );
INVx5_ASAP7_75t_L g221 ( .A(n_165), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_165), .B(n_235), .Y(n_234) );
NOR2x1_ASAP7_75t_SL g266 ( .A(n_165), .B(n_267), .Y(n_266) );
BUFx2_ASAP7_75t_L g311 ( .A(n_165), .Y(n_311) );
AND2x2_ASAP7_75t_L g413 ( .A(n_165), .B(n_183), .Y(n_413) );
OR2x6_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
AND2x2_ASAP7_75t_L g220 ( .A(n_173), .B(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_173), .Y(n_230) );
INVx4_ASAP7_75t_L g235 ( .A(n_173), .Y(n_235) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_180), .B(n_181), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_179), .Y(n_174) );
AOI21x1_ASAP7_75t_L g440 ( .A1(n_180), .A2(n_441), .B(n_447), .Y(n_440) );
INVx1_ASAP7_75t_L g278 ( .A(n_182), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_R g381 ( .A1(n_182), .A2(n_220), .B(n_252), .C(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g401 ( .A(n_182), .B(n_226), .Y(n_401) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_192), .Y(n_182) );
INVx1_ASAP7_75t_L g219 ( .A(n_183), .Y(n_219) );
INVx2_ASAP7_75t_L g225 ( .A(n_183), .Y(n_225) );
OR2x2_ASAP7_75t_L g244 ( .A(n_183), .B(n_235), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_183), .B(n_267), .Y(n_313) );
BUFx3_ASAP7_75t_L g320 ( .A(n_183), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_184), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_191), .Y(n_185) );
INVx1_ASAP7_75t_SL g194 ( .A(n_191), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_191), .B(n_216), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_191), .A2(n_460), .B(n_461), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_191), .A2(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g283 ( .A(n_192), .Y(n_283) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_192), .Y(n_296) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g229 ( .A(n_193), .Y(n_229) );
INVx1_ASAP7_75t_L g338 ( .A(n_193), .Y(n_338) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_201), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_194), .B(n_202), .Y(n_201) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_194), .A2(n_195), .B(n_201), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_200), .Y(n_195) );
AND2x2_ASAP7_75t_L g239 ( .A(n_203), .B(n_240), .Y(n_239) );
OAI31xp33_ASAP7_75t_L g390 ( .A1(n_203), .A2(n_391), .A3(n_393), .B(n_396), .Y(n_390) );
INVx1_ASAP7_75t_SL g408 ( .A(n_203), .Y(n_408) );
AND2x4_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
AOI21xp33_ASAP7_75t_L g222 ( .A1(n_204), .A2(n_223), .B(n_231), .Y(n_222) );
NAND2x1_ASAP7_75t_L g302 ( .A(n_204), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g331 ( .A(n_204), .Y(n_331) );
INVx2_ASAP7_75t_L g280 ( .A(n_205), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_205), .B(n_263), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_205), .B(n_262), .Y(n_372) );
NOR2xp33_ASAP7_75t_SL g380 ( .A(n_205), .B(n_331), .Y(n_380) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_217), .Y(n_205) );
AND2x2_ASAP7_75t_SL g249 ( .A(n_206), .B(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g260 ( .A(n_206), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g289 ( .A(n_206), .B(n_271), .Y(n_289) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
BUFx2_ASAP7_75t_L g253 ( .A(n_207), .Y(n_253) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
OAI21x1_ASAP7_75t_SL g208 ( .A1(n_209), .A2(n_211), .B(n_215), .Y(n_208) );
INVx1_ASAP7_75t_L g216 ( .A(n_210), .Y(n_216) );
INVx2_ASAP7_75t_L g261 ( .A(n_217), .Y(n_261) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_217), .Y(n_321) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
INVx1_ASAP7_75t_L g257 ( .A(n_219), .Y(n_257) );
AND2x2_ASAP7_75t_L g336 ( .A(n_219), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g247 ( .A(n_220), .B(n_241), .Y(n_247) );
INVx2_ASAP7_75t_SL g295 ( .A(n_220), .Y(n_295) );
INVx4_ASAP7_75t_L g226 ( .A(n_221), .Y(n_226) );
AND2x2_ASAP7_75t_L g324 ( .A(n_221), .B(n_267), .Y(n_324) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_221), .B(n_337), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g359 ( .A(n_221), .B(n_235), .Y(n_359) );
INVx1_ASAP7_75t_L g365 ( .A(n_223), .Y(n_365) );
OR2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_227), .Y(n_223) );
INVx1_ASAP7_75t_L g284 ( .A(n_224), .Y(n_284) );
OR2x2_ASAP7_75t_L g297 ( .A(n_224), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
OR2x2_ASAP7_75t_L g349 ( .A(n_225), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g379 ( .A(n_225), .B(n_267), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_226), .B(n_229), .Y(n_255) );
AND2x2_ASAP7_75t_L g347 ( .A(n_226), .B(n_337), .Y(n_347) );
AND2x4_ASAP7_75t_L g409 ( .A(n_226), .B(n_288), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
INVx2_ASAP7_75t_L g233 ( .A(n_228), .Y(n_233) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp67_ASAP7_75t_SL g232 ( .A(n_233), .B(n_234), .Y(n_232) );
OAI322xp33_ASAP7_75t_SL g245 ( .A1(n_233), .A2(n_246), .A3(n_248), .B1(n_251), .B2(n_254), .C1(n_256), .C2(n_258), .Y(n_245) );
INVx1_ASAP7_75t_L g403 ( .A(n_233), .Y(n_403) );
OR2x2_ASAP7_75t_L g256 ( .A(n_234), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g282 ( .A(n_235), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_235), .B(n_283), .Y(n_298) );
INVx2_ASAP7_75t_L g325 ( .A(n_235), .Y(n_325) );
AND2x4_ASAP7_75t_L g337 ( .A(n_235), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_SL g340 ( .A(n_237), .B(n_253), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_243), .B(n_245), .Y(n_238) );
AND2x2_ASAP7_75t_L g306 ( .A(n_240), .B(n_273), .Y(n_306) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_241), .B(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g264 ( .A(n_242), .Y(n_264) );
AND2x4_ASAP7_75t_SL g346 ( .A(n_242), .B(n_261), .Y(n_346) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g254 ( .A(n_244), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_247), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g382 ( .A(n_249), .B(n_346), .Y(n_382) );
NOR4xp25_ASAP7_75t_L g386 ( .A(n_249), .B(n_263), .C(n_303), .D(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g263 ( .A(n_250), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g299 ( .A(n_250), .B(n_274), .Y(n_299) );
AND2x4_ASAP7_75t_L g363 ( .A(n_250), .B(n_274), .Y(n_363) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_253), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
OR2x2_ASAP7_75t_L g352 ( .A(n_260), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g406 ( .A(n_260), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_261), .B(n_273), .Y(n_307) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AOI211xp5_ASAP7_75t_SL g265 ( .A1(n_266), .A2(n_268), .B(n_275), .C(n_290), .Y(n_265) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_273), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_271), .B(n_274), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_272), .B(n_277), .Y(n_276) );
BUFx2_ASAP7_75t_L g354 ( .A(n_272), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_273), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g369 ( .A(n_273), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_284), .B(n_285), .Y(n_281) );
AND2x4_ASAP7_75t_L g318 ( .A(n_282), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g412 ( .A(n_282), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_SL g316 ( .A(n_288), .Y(n_316) );
AND2x2_ASAP7_75t_L g375 ( .A(n_289), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g389 ( .A(n_289), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_293), .B(n_297), .C(n_299), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_291), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g367 ( .A(n_292), .B(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g388 ( .A(n_292), .B(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
OR2x2_ASAP7_75t_L g377 ( .A(n_295), .B(n_319), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_298), .A2(n_305), .B1(n_307), .B2(n_308), .Y(n_304) );
INVx1_ASAP7_75t_SL g395 ( .A(n_299), .Y(n_395) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_310), .B(n_319), .Y(n_361) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_313), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B1(n_321), .B2(n_322), .Y(n_314) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AOI21xp5_ASAP7_75t_SL g328 ( .A1(n_319), .A2(n_329), .B(n_332), .Y(n_328) );
AND2x2_ASAP7_75t_L g357 ( .A(n_319), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND3x2_ASAP7_75t_L g323 ( .A(n_320), .B(n_324), .C(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g385 ( .A(n_320), .B(n_342), .Y(n_385) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g370 ( .A(n_325), .B(n_371), .Y(n_370) );
NOR2xp67_ASAP7_75t_L g326 ( .A(n_327), .B(n_383), .Y(n_326) );
NAND4xp25_ASAP7_75t_L g327 ( .A(n_328), .B(n_343), .C(n_364), .D(n_381), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B1(n_339), .B2(n_341), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_335), .A2(n_349), .B1(n_369), .B2(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g350 ( .A(n_337), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_339), .A2(n_362), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx3_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .B1(n_348), .B2(n_351), .C(n_355), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_360), .B1(n_361), .B2(n_362), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_358), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_358), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B1(n_370), .B2(n_372), .C(n_373), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_367), .B(n_369), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .B1(n_378), .B2(n_380), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI211xp5_ASAP7_75t_SL g398 ( .A1(n_379), .A2(n_399), .B(n_400), .C(n_402), .Y(n_398) );
OAI211xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .B(n_390), .C(n_397), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_404), .B1(n_407), .B2(n_409), .C(n_410), .Y(n_397) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_415), .Y(n_414) );
CKINVDCx11_ASAP7_75t_R g415 ( .A(n_416), .Y(n_415) );
OR2x6_ASAP7_75t_SL g416 ( .A(n_417), .B(n_418), .Y(n_416) );
AND2x6_ASAP7_75t_SL g724 ( .A(n_417), .B(n_419), .Y(n_724) );
OR2x2_ASAP7_75t_L g733 ( .A(n_417), .B(n_419), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_417), .B(n_418), .Y(n_743) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_423), .B(n_753), .Y(n_752) );
INVx4_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2x1p5_ASAP7_75t_L g748 ( .A(n_424), .B(n_749), .Y(n_748) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_631), .Y(n_424) );
NOR3xp33_ASAP7_75t_SL g425 ( .A(n_426), .B(n_554), .C(n_589), .Y(n_425) );
OAI211xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_456), .B(n_506), .C(n_544), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_438), .Y(n_428) );
AND2x2_ASAP7_75t_L g537 ( .A(n_429), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_429), .B(n_543), .Y(n_577) );
AND2x2_ASAP7_75t_L g602 ( .A(n_429), .B(n_557), .Y(n_602) );
INVx4_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g509 ( .A(n_430), .Y(n_509) );
OR2x2_ASAP7_75t_L g540 ( .A(n_430), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g548 ( .A(n_430), .B(n_448), .Y(n_548) );
AND2x2_ASAP7_75t_L g556 ( .A(n_430), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g583 ( .A(n_430), .B(n_584), .Y(n_583) );
NOR2x1_ASAP7_75t_L g594 ( .A(n_430), .B(n_586), .Y(n_594) );
AND2x4_ASAP7_75t_L g611 ( .A(n_430), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g649 ( .A(n_430), .Y(n_649) );
AND2x4_ASAP7_75t_SL g654 ( .A(n_430), .B(n_439), .Y(n_654) );
OR2x6_ASAP7_75t_L g430 ( .A(n_431), .B(n_437), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_438), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_438), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_448), .Y(n_438) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_439), .Y(n_549) );
INVx2_ASAP7_75t_L g585 ( .A(n_439), .Y(n_585) );
INVx1_ASAP7_75t_L g612 ( .A(n_439), .Y(n_612) );
AND2x2_ASAP7_75t_L g711 ( .A(n_439), .B(n_621), .Y(n_711) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_440), .Y(n_543) );
AND2x2_ASAP7_75t_L g557 ( .A(n_440), .B(n_448), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_446), .Y(n_441) );
INVx2_ASAP7_75t_L g586 ( .A(n_448), .Y(n_586) );
INVx2_ASAP7_75t_L g621 ( .A(n_448), .Y(n_621) );
OR2x2_ASAP7_75t_L g706 ( .A(n_448), .B(n_538), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_454), .Y(n_449) );
AOI211xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_473), .B(n_493), .C(n_500), .Y(n_456) );
INVx2_ASAP7_75t_SL g595 ( .A(n_457), .Y(n_595) );
AND2x2_ASAP7_75t_L g601 ( .A(n_457), .B(n_474), .Y(n_601) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_465), .Y(n_457) );
INVx1_ASAP7_75t_L g497 ( .A(n_458), .Y(n_497) );
INVx1_ASAP7_75t_L g503 ( .A(n_458), .Y(n_503) );
INVx2_ASAP7_75t_L g528 ( .A(n_458), .Y(n_528) );
AND2x2_ASAP7_75t_L g552 ( .A(n_458), .B(n_476), .Y(n_552) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_458), .Y(n_581) );
OR2x2_ASAP7_75t_L g661 ( .A(n_458), .B(n_484), .Y(n_661) );
AND2x2_ASAP7_75t_L g527 ( .A(n_465), .B(n_528), .Y(n_527) );
NOR2x1_ASAP7_75t_SL g559 ( .A(n_465), .B(n_484), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .Y(n_466) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g573 ( .A(n_474), .B(n_496), .Y(n_573) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
OR2x2_ASAP7_75t_L g505 ( .A(n_475), .B(n_484), .Y(n_505) );
BUFx2_ASAP7_75t_L g529 ( .A(n_475), .Y(n_529) );
NOR2xp67_ASAP7_75t_L g580 ( .A(n_475), .B(n_581), .Y(n_580) );
INVx4_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_476), .Y(n_532) );
AND2x2_ASAP7_75t_L g558 ( .A(n_476), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g568 ( .A(n_476), .Y(n_568) );
NAND2x1_ASAP7_75t_L g606 ( .A(n_476), .B(n_484), .Y(n_606) );
OR2x2_ASAP7_75t_L g681 ( .A(n_476), .B(n_498), .Y(n_681) );
OR2x6_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx2_ASAP7_75t_SL g494 ( .A(n_484), .Y(n_494) );
AND2x2_ASAP7_75t_L g553 ( .A(n_484), .B(n_498), .Y(n_553) );
AND2x2_ASAP7_75t_L g624 ( .A(n_484), .B(n_625), .Y(n_624) );
BUFx2_ASAP7_75t_L g645 ( .A(n_484), .Y(n_645) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_492), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g567 ( .A(n_496), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
BUFx2_ASAP7_75t_L g562 ( .A(n_497), .Y(n_562) );
AND2x2_ASAP7_75t_L g534 ( .A(n_498), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g625 ( .A(n_498), .Y(n_625) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
OR2x2_ASAP7_75t_L g571 ( .A(n_502), .B(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_SL g613 ( .A(n_502), .B(n_614), .Y(n_613) );
AOI322xp5_ASAP7_75t_L g650 ( .A1(n_502), .A2(n_529), .A3(n_651), .B1(n_653), .B2(n_656), .C1(n_658), .C2(n_660), .Y(n_650) );
AND2x2_ASAP7_75t_L g715 ( .A(n_502), .B(n_716), .Y(n_715) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_503), .B(n_529), .Y(n_539) );
AOI322xp5_ASAP7_75t_L g590 ( .A1(n_504), .A2(n_591), .A3(n_595), .B1(n_596), .B2(n_599), .C1(n_601), .C2(n_602), .Y(n_590) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g642 ( .A(n_505), .B(n_595), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_505), .A2(n_702), .B1(n_704), .B2(n_707), .Y(n_701) );
OR2x2_ASAP7_75t_L g719 ( .A(n_505), .B(n_668), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_529), .B(n_530), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
AOI221xp5_ASAP7_75t_SL g569 ( .A1(n_508), .A2(n_545), .B1(n_570), .B2(n_573), .C(n_574), .Y(n_569) );
AND2x2_ASAP7_75t_L g596 ( .A(n_508), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_509), .B(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g638 ( .A(n_509), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g667 ( .A(n_510), .Y(n_667) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_527), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_511), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g609 ( .A(n_511), .Y(n_609) );
OR2x2_ASAP7_75t_L g616 ( .A(n_511), .B(n_617), .Y(n_616) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g659 ( .A(n_512), .B(n_621), .Y(n_659) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
AND2x4_ASAP7_75t_L g538 ( .A(n_513), .B(n_514), .Y(n_538) );
AND2x4_ASAP7_75t_L g516 ( .A(n_517), .B(n_520), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
NOR2x1p5_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_527), .B(n_588), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_527), .B(n_568), .Y(n_664) );
INVx1_ASAP7_75t_L g668 ( .A(n_527), .Y(n_668) );
INVx1_ASAP7_75t_L g535 ( .A(n_528), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_536), .B1(n_539), .B2(n_540), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_SL g646 ( .A(n_534), .Y(n_646) );
AND2x2_ASAP7_75t_L g703 ( .A(n_535), .B(n_559), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_537), .B(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_SL g575 ( .A(n_537), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_537), .B(n_696), .Y(n_695) );
BUFx3_ASAP7_75t_L g563 ( .A(n_538), .Y(n_563) );
INVx2_ASAP7_75t_L g593 ( .A(n_538), .Y(n_593) );
AND2x2_ASAP7_75t_L g636 ( .A(n_538), .B(n_620), .Y(n_636) );
INVx1_ASAP7_75t_L g550 ( .A(n_540), .Y(n_550) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OAI21xp5_ASAP7_75t_SL g544 ( .A1(n_545), .A2(n_550), .B(n_551), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g629 ( .A(n_548), .Y(n_629) );
INVx2_ASAP7_75t_L g617 ( .A(n_549), .Y(n_617) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_L g614 ( .A(n_553), .B(n_568), .Y(n_614) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_553), .A2(n_651), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_555), .B(n_569), .Y(n_554) );
AOI32xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_558), .A3(n_560), .B1(n_564), .B2(n_567), .Y(n_555) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_556), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_556), .A2(n_645), .B1(n_663), .B2(n_665), .C(n_671), .Y(n_662) );
AND2x2_ASAP7_75t_L g682 ( .A(n_556), .B(n_563), .Y(n_682) );
BUFx2_ASAP7_75t_L g566 ( .A(n_557), .Y(n_566) );
INVx1_ASAP7_75t_L g691 ( .A(n_557), .Y(n_691) );
INVx1_ASAP7_75t_L g696 ( .A(n_557), .Y(n_696) );
INVx1_ASAP7_75t_SL g689 ( .A(n_558), .Y(n_689) );
INVx2_ASAP7_75t_L g572 ( .A(n_559), .Y(n_572) );
AND2x2_ASAP7_75t_L g684 ( .A(n_560), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g656 ( .A(n_562), .B(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g628 ( .A(n_563), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_563), .B(n_654), .Y(n_676) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g588 ( .A(n_568), .Y(n_588) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g578 ( .A(n_572), .B(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g587 ( .A(n_572), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g692 ( .A(n_573), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_578), .B1(n_582), .B2(n_587), .Y(n_574) );
INVx2_ASAP7_75t_SL g666 ( .A(n_576), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_576), .B(n_705), .Y(n_707) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_578), .A2(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g623 ( .A(n_580), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g651 ( .A(n_583), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g598 ( .A(n_584), .Y(n_598) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g640 ( .A(n_586), .Y(n_640) );
INVx1_ASAP7_75t_L g685 ( .A(n_587), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_603), .C(n_626), .Y(n_589) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
INVx2_ASAP7_75t_L g652 ( .A(n_592), .Y(n_652) );
AND2x2_ASAP7_75t_L g670 ( .A(n_592), .B(n_611), .Y(n_670) );
OR2x2_ASAP7_75t_L g709 ( .A(n_592), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_593), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g605 ( .A(n_595), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g672 ( .A(n_598), .B(n_609), .Y(n_672) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_601), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g713 ( .A(n_601), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_607), .B1(n_611), .B2(n_613), .C(n_615), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g626 ( .A1(n_604), .A2(n_627), .B(n_630), .Y(n_626) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx3_ASAP7_75t_L g657 ( .A(n_606), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_606), .B(n_700), .Y(n_699) );
INVxp33_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g618 ( .A(n_614), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .B1(n_619), .B2(n_622), .Y(n_615) );
INVx2_ASAP7_75t_L g721 ( .A(n_617), .Y(n_721) );
BUFx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVxp67_ASAP7_75t_L g700 ( .A(n_625), .Y(n_700) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
NOR2x1_ASAP7_75t_L g631 ( .A(n_632), .B(n_677), .Y(n_631) );
NAND4xp25_ASAP7_75t_L g632 ( .A(n_633), .B(n_650), .C(n_662), .D(n_674), .Y(n_632) );
O2A1O1Ixp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_637), .B(n_641), .C(n_643), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g673 ( .A(n_636), .Y(n_673) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI21xp5_ASAP7_75t_L g643 ( .A1(n_638), .A2(n_644), .B(n_647), .Y(n_643) );
INVx2_ASAP7_75t_L g722 ( .A(n_639), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_640), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g655 ( .A(n_640), .Y(n_655) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
OR2x2_ASAP7_75t_L g717 ( .A(n_645), .B(n_681), .Y(n_717) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_652), .Y(n_688) );
AND2x2_ASAP7_75t_SL g653 ( .A(n_654), .B(n_655), .Y(n_653) );
AND2x2_ASAP7_75t_L g658 ( .A(n_654), .B(n_659), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_654), .A2(n_684), .B(n_686), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_654), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_SL g712 ( .A(n_654), .Y(n_712) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI22xp33_ASAP7_75t_SL g665 ( .A1(n_666), .A2(n_667), .B1(n_668), .B2(n_669), .Y(n_665) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NAND4xp25_ASAP7_75t_L g677 ( .A(n_678), .B(n_683), .C(n_693), .D(n_714), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_682), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B1(n_690), .B2(n_692), .Y(n_686) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI211xp5_ASAP7_75t_SL g693 ( .A1(n_694), .A2(n_697), .B(n_701), .C(n_708), .Y(n_693) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_712), .B(n_713), .Y(n_708) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
OAI21xp5_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_718), .B(n_720), .Y(n_714) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx3_ASAP7_75t_SL g727 ( .A(n_723), .Y(n_727) );
CKINVDCx5p33_ASAP7_75t_R g723 ( .A(n_724), .Y(n_723) );
CKINVDCx6p67_ASAP7_75t_R g726 ( .A(n_727), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx3_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_742), .Y(n_735) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_738), .B(n_741), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_SL g759 ( .A(n_739), .B(n_741), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_739), .A2(n_764), .B(n_767), .Y(n_763) );
BUFx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
BUFx2_ASAP7_75t_R g746 ( .A(n_743), .Y(n_746) );
BUFx2_ASAP7_75t_L g768 ( .A(n_743), .Y(n_768) );
INVxp67_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B(n_754), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_746), .B(n_755), .Y(n_754) );
NAND2x1_ASAP7_75t_L g747 ( .A(n_748), .B(n_752), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_749), .Y(n_753) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
CKINVDCx11_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
CKINVDCx8_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
endmodule