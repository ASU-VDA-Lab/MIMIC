module fake_jpeg_6536_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_33),
.B1(n_18),
.B2(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_33),
.B1(n_18),
.B2(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_57),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_59),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_24),
.B1(n_18),
.B2(n_33),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_18),
.B1(n_17),
.B2(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_74),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_69),
.B(n_76),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_42),
.B1(n_39),
.B2(n_38),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_61),
.B1(n_64),
.B2(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_78),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_86),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_81),
.Y(n_121)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_84),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_21),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_16),
.B1(n_20),
.B2(n_23),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_86),
.B(n_77),
.C(n_71),
.Y(n_117)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_96),
.Y(n_111)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_47),
.A2(n_23),
.B1(n_17),
.B2(n_32),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_38),
.C(n_19),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_116),
.B1(n_84),
.B2(n_72),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_63),
.C(n_62),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_67),
.C(n_91),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_114),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_55),
.B(n_53),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_115),
.B(n_32),
.Y(n_135)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_SL g115 ( 
.A(n_76),
.B(n_21),
.C(n_23),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_61),
.B1(n_63),
.B2(n_62),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_86),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_51),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_122),
.Y(n_131)
);

AO21x2_ASAP7_75t_L g119 ( 
.A1(n_70),
.A2(n_61),
.B(n_42),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_72),
.B1(n_64),
.B2(n_98),
.Y(n_141)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_95),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_51),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_128),
.A2(n_151),
.B1(n_158),
.B2(n_125),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_119),
.A2(n_79),
.B1(n_62),
.B2(n_63),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_141),
.B1(n_145),
.B2(n_119),
.Y(n_160)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_136),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_89),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_148),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_134),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_142),
.B(n_109),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_138),
.A2(n_34),
.B1(n_31),
.B2(n_22),
.Y(n_193)
);

OR2x2_ASAP7_75t_SL g139 ( 
.A(n_103),
.B(n_0),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_146),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_144),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_68),
.B(n_69),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_54),
.B1(n_92),
.B2(n_80),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_19),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_19),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_67),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_75),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_156),
.Y(n_179)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_152),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_108),
.A2(n_74),
.B1(n_42),
.B2(n_39),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_90),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_16),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_108),
.B(n_26),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_0),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_20),
.B1(n_26),
.B2(n_30),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_160),
.Y(n_200)
);

OAI32xp33_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_108),
.A3(n_105),
.B1(n_119),
.B2(n_115),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_164),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_162),
.A2(n_169),
.B(n_175),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_127),
.C(n_105),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_167),
.A2(n_183),
.B1(n_190),
.B2(n_141),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_109),
.B1(n_125),
.B2(n_106),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_168),
.A2(n_189),
.B1(n_151),
.B2(n_128),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_30),
.B(n_100),
.C(n_38),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_170),
.B(n_177),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_133),
.C(n_147),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_176),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_156),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_184),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_26),
.B(n_19),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_150),
.B(n_120),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_19),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_187),
.Y(n_195)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_138),
.A2(n_65),
.B1(n_99),
.B2(n_113),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_137),
.B(n_99),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_191),
.Y(n_207)
);

CKINVDCx10_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_186),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_1),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_147),
.A2(n_65),
.B1(n_29),
.B2(n_22),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_25),
.B(n_2),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_101),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_198),
.A2(n_216),
.B1(n_210),
.B2(n_206),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_147),
.B1(n_142),
.B2(n_139),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_214),
.B1(n_220),
.B2(n_193),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_139),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_208),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_211),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_215),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_155),
.B1(n_154),
.B2(n_132),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_1),
.Y(n_217)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

AOI22x1_ASAP7_75t_L g220 ( 
.A1(n_161),
.A2(n_29),
.B1(n_22),
.B2(n_31),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_132),
.Y(n_222)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_232),
.B1(n_246),
.B2(n_198),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_171),
.C(n_180),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_229),
.C(n_235),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_238),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_162),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_190),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_164),
.C(n_179),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_163),
.B(n_176),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_230),
.A2(n_241),
.B(n_243),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_200),
.A2(n_160),
.B1(n_163),
.B2(n_173),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_179),
.C(n_174),
.Y(n_235)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_221),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_174),
.C(n_175),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_174),
.C(n_166),
.Y(n_262)
);

AO22x1_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_199),
.B1(n_213),
.B2(n_207),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_220),
.A2(n_175),
.B(n_172),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_203),
.A2(n_169),
.B1(n_185),
.B2(n_166),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_248),
.A2(n_34),
.B1(n_25),
.B2(n_3),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_196),
.B1(n_201),
.B2(n_197),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_265),
.B1(n_236),
.B2(n_226),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_218),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_257),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_217),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_194),
.Y(n_255)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_256),
.B(n_258),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_204),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

FAx1_ASAP7_75t_SL g259 ( 
.A(n_239),
.B(n_241),
.CI(n_231),
.CON(n_259),
.SN(n_259)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_263),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_262),
.C(n_266),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_188),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_267),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_188),
.B1(n_132),
.B2(n_29),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_25),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_29),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_25),
.C(n_22),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_243),
.C(n_25),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_247),
.Y(n_271)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_275),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_230),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_279),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_251),
.A2(n_241),
.B1(n_236),
.B2(n_234),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_224),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_259),
.A2(n_234),
.B1(n_228),
.B2(n_247),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_9),
.B(n_15),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_25),
.C(n_34),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_34),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_250),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_284),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_260),
.B(n_248),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_288),
.A2(n_291),
.B(n_295),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_SL g291 ( 
.A1(n_274),
.A2(n_262),
.A3(n_253),
.B1(n_281),
.B2(n_261),
.C1(n_266),
.C2(n_280),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_268),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_292),
.B(n_294),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_260),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_253),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_299),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_281),
.C(n_277),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_14),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_279),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_309),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_303),
.B(n_306),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_310),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_272),
.C(n_282),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_278),
.C(n_2),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_289),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_311),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_11),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_296),
.A2(n_9),
.B(n_8),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_306),
.A2(n_290),
.B1(n_297),
.B2(n_298),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_316),
.B(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_290),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_8),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_4),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_303),
.B(n_5),
.Y(n_322)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_8),
.A3(n_9),
.B1(n_6),
.B2(n_7),
.C1(n_4),
.C2(n_5),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_4),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_323),
.B(n_326),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_300),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_324),
.A2(n_325),
.B(n_320),
.C(n_313),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

AOI321xp33_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_329),
.A3(n_328),
.B1(n_301),
.B2(n_6),
.C(n_7),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_321),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_4),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_5),
.C(n_7),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_7),
.Y(n_333)
);


endmodule