module fake_jpeg_232_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_5),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_40),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_34),
.Y(n_72)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

OR2x2_ASAP7_75t_SL g36 ( 
.A(n_12),
.B(n_0),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_15),
.C(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_39),
.B(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_4),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_14),
.B(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_24),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_13),
.B(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_13),
.B(n_2),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_23),
.B1(n_26),
.B2(n_18),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_50),
.B1(n_67),
.B2(n_57),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_26),
.B1(n_18),
.B2(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_52),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_63),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_30),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_27),
.B1(n_35),
.B2(n_31),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_69),
.B1(n_50),
.B2(n_48),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_75),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_29),
.CI(n_66),
.CON(n_76),
.SN(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_77),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_80),
.B1(n_85),
.B2(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_62),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_49),
.B1(n_64),
.B2(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_53),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_72),
.B1(n_71),
.B2(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_89),
.B1(n_49),
.B2(n_74),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_54),
.B(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_96),
.Y(n_109)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_78),
.B(n_80),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_103),
.B(n_76),
.C(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_85),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_76),
.B(n_77),
.Y(n_103)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_95),
.B(n_104),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_107),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_99),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_92),
.B(n_103),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_121),
.B(n_113),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_93),
.C(n_91),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_108),
.C(n_106),
.Y(n_122)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_123),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_126),
.Y(n_128)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_113),
.C(n_112),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_125),
.B(n_120),
.Y(n_129)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_112),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_127),
.A2(n_119),
.B(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g133 ( 
.A(n_132),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_127),
.B(n_128),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_133),
.B(n_130),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_130),
.Y(n_137)
);


endmodule