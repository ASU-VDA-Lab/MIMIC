module fake_jpeg_7615_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_47),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

INVx2_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_58),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_29),
.B1(n_26),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_51),
.A2(n_52),
.B1(n_68),
.B2(n_69),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_29),
.B1(n_26),
.B2(n_23),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_22),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_16),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_28),
.B1(n_18),
.B2(n_35),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_33),
.B(n_21),
.Y(n_87)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_37),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_71),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_28),
.B1(n_18),
.B2(n_35),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_35),
.B1(n_18),
.B2(n_32),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_20),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_73),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_48),
.B(n_55),
.C(n_65),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_74),
.A2(n_113),
.B(n_11),
.C(n_15),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_75),
.B(n_79),
.Y(n_137)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_38),
.B1(n_32),
.B2(n_47),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_82),
.A2(n_94),
.B1(n_96),
.B2(n_102),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_47),
.B1(n_38),
.B2(n_32),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_83),
.A2(n_85),
.B1(n_89),
.B2(n_111),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_24),
.B1(n_27),
.B2(n_21),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_87),
.A2(n_95),
.B(n_45),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_24),
.B1(n_21),
.B2(n_34),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_30),
.B1(n_34),
.B2(n_14),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_30),
.B(n_41),
.C(n_43),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_31),
.Y(n_97)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_31),
.Y(n_99)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_34),
.B1(n_24),
.B2(n_31),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_70),
.B1(n_56),
.B2(n_46),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_61),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_114),
.B1(n_56),
.B2(n_72),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_59),
.A2(n_34),
.B1(n_46),
.B2(n_40),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_43),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_72),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_69),
.A2(n_10),
.B1(n_8),
.B2(n_7),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_12),
.B(n_1),
.Y(n_138)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_68),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_0),
.B(n_1),
.Y(n_135)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_60),
.A2(n_45),
.B1(n_40),
.B2(n_37),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_64),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_54),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_115),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_120),
.B1(n_124),
.B2(n_128),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_121),
.B(n_136),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_46),
.B1(n_45),
.B2(n_40),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_122),
.A2(n_103),
.B1(n_93),
.B2(n_111),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_79),
.A2(n_11),
.B1(n_15),
.B2(n_12),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_125),
.B(n_130),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_141),
.B(n_142),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_77),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_107),
.B(n_87),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_77),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_76),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_0),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_81),
.B(n_0),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_145),
.B(n_1),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_148),
.A2(n_170),
.B(n_119),
.Y(n_201)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_153),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_150),
.B(n_119),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_76),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_171),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_88),
.B(n_84),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_152),
.A2(n_132),
.B(n_41),
.Y(n_210)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_92),
.B1(n_110),
.B2(n_96),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_81),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_157),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_139),
.B1(n_136),
.B2(n_121),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_158),
.A2(n_165),
.B1(n_166),
.B2(n_117),
.Y(n_204)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_160),
.Y(n_192)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_78),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_167),
.Y(n_189)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

CKINVDCx10_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_163),
.Y(n_194)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_98),
.B1(n_95),
.B2(n_84),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_88),
.B1(n_89),
.B2(n_78),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_78),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_169),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_74),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_138),
.A2(n_92),
.B1(n_113),
.B2(n_85),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_83),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_112),
.Y(n_172)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_1),
.B(n_2),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_108),
.C(n_114),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_104),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_175),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_118),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_176),
.B(n_118),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_115),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_177),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_91),
.B1(n_86),
.B2(n_126),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_144),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_181),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_128),
.B(n_122),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_182),
.A2(n_203),
.B(n_206),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_183),
.B(n_200),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_191),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_168),
.C(n_161),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_173),
.C(n_152),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_145),
.B(n_142),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_196),
.A2(n_201),
.B(n_202),
.Y(n_215)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_153),
.A2(n_156),
.B1(n_152),
.B2(n_148),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_147),
.A2(n_117),
.B(n_116),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_204),
.A2(n_207),
.B(n_210),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_205),
.B(n_2),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_131),
.B(n_43),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_151),
.B(n_166),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_54),
.B1(n_43),
.B2(n_41),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_165),
.A2(n_132),
.B1(n_126),
.B2(n_72),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_209),
.A2(n_163),
.B1(n_176),
.B2(n_160),
.Y(n_218)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_213),
.Y(n_250)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_229),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_149),
.C(n_174),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_226),
.C(n_238),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_218),
.A2(n_209),
.B1(n_184),
.B2(n_180),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_186),
.A2(n_171),
.B1(n_178),
.B2(n_159),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_220),
.A2(n_202),
.B1(n_188),
.B2(n_201),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_143),
.Y(n_221)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_230),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_164),
.C(n_43),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_228),
.C(n_236),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_225),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_43),
.C(n_41),
.Y(n_226)
);

BUFx8_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_227),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_41),
.C(n_54),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_237),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_2),
.Y(n_232)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_41),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_183),
.B(n_2),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_184),
.B(n_3),
.C(n_4),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_240),
.B(n_215),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_257),
.B1(n_258),
.B2(n_212),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_200),
.Y(n_247)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_219),
.A2(n_181),
.B1(n_208),
.B2(n_204),
.Y(n_251)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_220),
.A2(n_233),
.B1(n_224),
.B2(n_211),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_252),
.B(n_233),
.Y(n_261)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_216),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_254),
.Y(n_270)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_206),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_259),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_211),
.A2(n_203),
.B1(n_210),
.B2(n_198),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_224),
.A2(n_185),
.B1(n_197),
.B2(n_194),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_182),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_261),
.A2(n_245),
.B(n_191),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_253),
.B(n_185),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_262),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_217),
.C(n_223),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_267),
.C(n_269),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_265),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_215),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_235),
.Y(n_266)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_228),
.Y(n_267)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_226),
.C(n_236),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_222),
.C(n_213),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_239),
.C(n_252),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_194),
.C(n_197),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_276),
.B1(n_244),
.B2(n_250),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_238),
.B(n_229),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_279),
.B(n_276),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_227),
.C(n_191),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_227),
.Y(n_277)
);

NOR2x1_ASAP7_75t_R g293 ( 
.A(n_277),
.B(n_190),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_257),
.B(n_190),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_280),
.A2(n_254),
.B1(n_250),
.B2(n_251),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_293),
.C(n_4),
.Y(n_308)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_241),
.B1(n_246),
.B2(n_243),
.Y(n_288)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_272),
.A2(n_241),
.B1(n_244),
.B2(n_247),
.Y(n_289)
);

AOI221xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_292),
.B1(n_295),
.B2(n_296),
.C(n_3),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_264),
.A2(n_243),
.B1(n_248),
.B2(n_242),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_277),
.C(n_265),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_270),
.A2(n_248),
.B1(n_190),
.B2(n_245),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_275),
.Y(n_297)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_297),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_280),
.B(n_273),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_301),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_302),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_269),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_263),
.B(n_191),
.C(n_5),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_306),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_305),
.A2(n_308),
.B1(n_293),
.B2(n_283),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_3),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_287),
.B(n_4),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_307),
.B(n_297),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_6),
.C(n_286),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_296),
.C(n_295),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_311),
.B(n_312),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_301),
.C(n_281),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_309),
.B(n_289),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_318),
.A3(n_298),
.B1(n_286),
.B2(n_300),
.C1(n_283),
.C2(n_304),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_320),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_321),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_317),
.A2(n_306),
.B1(n_303),
.B2(n_288),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_316),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_285),
.C(n_6),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_285),
.C(n_6),
.Y(n_324)
);

AOI21x1_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_318),
.B(n_319),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_328),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_325),
.B(n_327),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_314),
.B(n_311),
.Y(n_333)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_333),
.Y(n_334)
);


endmodule