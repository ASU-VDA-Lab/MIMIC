module real_jpeg_22842_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_2),
.A2(n_25),
.B1(n_28),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_2),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_2),
.A2(n_35),
.B1(n_105),
.B2(n_150),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_2),
.A2(n_53),
.B1(n_54),
.B2(n_150),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_2),
.A2(n_70),
.B1(n_71),
.B2(n_150),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_4),
.A2(n_105),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_4),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_24),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_158),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_4),
.B(n_66),
.C(n_71),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_4),
.B(n_52),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_4),
.A2(n_90),
.B1(n_253),
.B2(n_256),
.Y(n_255)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_6),
.A2(n_25),
.B1(n_28),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_6),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_152),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_6),
.A2(n_70),
.B1(n_71),
.B2(n_152),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_6),
.A2(n_31),
.B1(n_114),
.B2(n_152),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_7),
.A2(n_35),
.B1(n_42),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_7),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_7),
.A2(n_25),
.B1(n_28),
.B2(n_161),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_7),
.A2(n_53),
.B1(n_54),
.B2(n_161),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_7),
.A2(n_70),
.B1(n_71),
.B2(n_161),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_8),
.A2(n_33),
.B1(n_57),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_8),
.A2(n_57),
.B1(n_70),
.B2(n_71),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_9),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_9),
.A2(n_25),
.B1(n_28),
.B2(n_34),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_9),
.A2(n_34),
.B1(n_53),
.B2(n_54),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_9),
.A2(n_34),
.B1(n_70),
.B2(n_71),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_11),
.A2(n_33),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_11),
.A2(n_25),
.B1(n_28),
.B2(n_39),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_11),
.A2(n_39),
.B1(n_53),
.B2(n_54),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_11),
.A2(n_39),
.B1(n_70),
.B2(n_71),
.Y(n_140)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_14),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_14),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_14),
.A2(n_35),
.B1(n_74),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_14),
.A2(n_25),
.B1(n_28),
.B2(n_74),
.Y(n_119)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_15),
.Y(n_93)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_15),
.Y(n_144)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_15),
.Y(n_239)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_15),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_123),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_108),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_19),
.B(n_108),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_75),
.C(n_86),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g332 ( 
.A(n_20),
.B(n_75),
.CI(n_86),
.CON(n_332),
.SN(n_332)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_44),
.B2(n_45),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_21),
.A2(n_22),
.B1(n_110),
.B2(n_121),
.Y(n_109)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_22),
.B(n_47),
.C(n_61),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_30),
.B(n_36),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_23),
.B(n_38),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_23),
.A2(n_154),
.B1(n_155),
.B2(n_159),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_23),
.B(n_104),
.Y(n_309)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_24),
.A2(n_40),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_24),
.A2(n_40),
.B1(n_160),
.B2(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_24),
.A2(n_40),
.B1(n_168),
.B2(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_25),
.A2(n_28),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_25),
.A2(n_29),
.B(n_157),
.C(n_173),
.Y(n_172)
);

HAxp5_ASAP7_75t_SL g201 ( 
.A(n_25),
.B(n_158),
.CON(n_201),
.SN(n_201)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_29),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_27),
.B(n_28),
.C(n_32),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g200 ( 
.A1(n_28),
.A2(n_51),
.A3(n_54),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_30),
.Y(n_112)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_32),
.B(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_40),
.A2(n_103),
.B(n_107),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_40),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_40),
.A2(n_290),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_61),
.B2(n_62),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_55),
.B(n_58),
.Y(n_47)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_48),
.B(n_60),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_48),
.A2(n_52),
.B1(n_192),
.B2(n_201),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

AO22x1_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_50),
.B(n_53),
.Y(n_202)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_52),
.B(n_119),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_54),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_54),
.B(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_59),
.A2(n_77),
.B(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_61),
.A2(n_62),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_69),
.B(n_72),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_64),
.A2(n_73),
.B(n_100),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_64),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_64),
.A2(n_82),
.B(n_208),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_64),
.A2(n_207),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_64),
.A2(n_206),
.B1(n_207),
.B2(n_226),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_64),
.A2(n_99),
.B1(n_207),
.B2(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_66),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_85),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_69),
.A2(n_83),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_69),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_69),
.B(n_158),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_70),
.B(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_75),
.A2(n_76),
.B(n_80),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_77),
.A2(n_79),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_77),
.A2(n_118),
.B(n_151),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_77),
.A2(n_79),
.B1(n_149),
.B2(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_78),
.A2(n_79),
.B(n_120),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B(n_101),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_87),
.B(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_98),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_88),
.A2(n_89),
.B1(n_98),
.B2(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_88),
.A2(n_89),
.B1(n_101),
.B2(n_102),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_94),
.B(n_96),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_90),
.A2(n_137),
.B(n_139),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_90),
.A2(n_96),
.B(n_139),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_90),
.A2(n_236),
.B(n_237),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_90),
.A2(n_94),
.B1(n_244),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_91),
.A2(n_138),
.B1(n_143),
.B2(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_91),
.B(n_140),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_91),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_92),
.Y(n_186)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_97),
.B(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_98),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_122),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_119),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_329),
.B(n_333),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_316),
.B(n_328),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_298),
.B(n_315),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_193),
.B(n_275),
.C(n_297),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_178),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_131),
.B(n_178),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_164),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_145),
.B1(n_162),
.B2(n_163),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_133),
.B(n_163),
.C(n_164),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_134),
.B(n_136),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_135),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_144),
.Y(n_260)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_153),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_181),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_153),
.B(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_158),
.B(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_167),
.B(n_169),
.C(n_171),
.Y(n_295)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_186),
.B(n_187),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.C(n_184),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_179),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_182),
.B(n_184),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_188),
.B1(n_189),
.B2(n_213),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_185),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_187),
.B(n_237),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_270),
.B(n_274),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_220),
.B(n_269),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_209),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_198),
.B(n_209),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.C(n_205),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_199),
.B(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_203),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_204),
.B(n_205),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_214),
.B2(n_215),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_210),
.B(n_217),
.C(n_219),
.Y(n_271)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_216),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_264),
.B(n_268),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_240),
.B(n_263),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_223),
.B(n_229),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_227),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_234),
.C(n_235),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_249),
.B(n_262),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_248),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_254),
.B(n_261),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_251),
.B(n_252),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_265),
.B(n_266),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_277),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_295),
.B2(n_296),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_286),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_286),
.C(n_296),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_285),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_285),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_283),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_294),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_291),
.C(n_294),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_299),
.B(n_300),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_314),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_304),
.B1(n_312),
.B2(n_313),
.Y(n_301)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_313),
.C(n_314),
.Y(n_317)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_308),
.C(n_310),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_310),
.B2(n_311),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_317),
.B(n_318),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_326),
.B2(n_327),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_321),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_325),
.C(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_331),
.B(n_332),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_332),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);


endmodule