module fake_jpeg_7774_n_83 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_24),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_44),
.Y(n_54)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_46),
.Y(n_56)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_5),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_0),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_4),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

AO22x1_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_64)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_58),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_61),
.B(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_35),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_34),
.B1(n_7),
.B2(n_9),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_21),
.C(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_68),
.B1(n_64),
.B2(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_74),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_54),
.C(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_72),
.B(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_67),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_68),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_69),
.Y(n_81)
);

A2O1A1O1Ixp25_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_23),
.B(n_25),
.C(n_26),
.D(n_27),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_29),
.Y(n_83)
);


endmodule