module fake_netlist_5_1705_n_4408 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_111, n_483, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_355, n_486, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_479, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_213, n_129, n_342, n_482, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_85, n_463, n_239, n_466, n_420, n_55, n_49, n_310, n_54, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_441, n_450, n_312, n_476, n_429, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_4408);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_111;
input n_483;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_213;
input n_129;
input n_342;
input n_482;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_85;
input n_463;
input n_239;
input n_466;
input n_420;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_4408;

wire n_924;
wire n_1263;
wire n_3304;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_3912;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_3241;
wire n_4129;
wire n_549;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_532;
wire n_1161;
wire n_3795;
wire n_3863;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_3732;
wire n_1488;
wire n_4250;
wire n_667;
wire n_2955;
wire n_2899;
wire n_790;
wire n_3619;
wire n_1055;
wire n_3541;
wire n_3622;
wire n_4112;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_4337;
wire n_2395;
wire n_3906;
wire n_4127;
wire n_880;
wire n_4138;
wire n_3086;
wire n_3297;
wire n_544;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_552;
wire n_1528;
wire n_4217;
wire n_4395;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_4292;
wire n_2568;
wire n_3641;
wire n_956;
wire n_564;
wire n_4240;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_4236;
wire n_3088;
wire n_4202;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_551;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_1466;
wire n_1695;
wire n_688;
wire n_2487;
wire n_3766;
wire n_1353;
wire n_800;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_3813;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_671;
wire n_4238;
wire n_819;
wire n_1451;
wire n_1022;
wire n_4109;
wire n_2302;
wire n_915;
wire n_4038;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3599;
wire n_3571;
wire n_3785;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_3621;
wire n_4211;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_3039;
wire n_3019;
wire n_2011;
wire n_2096;
wire n_4013;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_877;
wire n_2105;
wire n_2538;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_4242;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_3710;
wire n_4243;
wire n_3851;
wire n_1860;
wire n_2543;
wire n_4155;
wire n_1359;
wire n_530;
wire n_1728;
wire n_2031;
wire n_556;
wire n_2076;
wire n_1107;
wire n_2482;
wire n_3036;
wire n_3891;
wire n_4145;
wire n_2677;
wire n_1230;
wire n_4144;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3832;
wire n_4374;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_3987;
wire n_4131;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_659;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_4021;
wire n_579;
wire n_1698;
wire n_3880;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_3624;
wire n_3834;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_3796;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_3937;
wire n_3696;
wire n_519;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_4315;
wire n_546;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_3782;
wire n_1845;
wire n_2193;
wire n_2052;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_3810;
wire n_2466;
wire n_1517;
wire n_2091;
wire n_2652;
wire n_2635;
wire n_4311;
wire n_1289;
wire n_4264;
wire n_3631;
wire n_2715;
wire n_3806;
wire n_3087;
wire n_4197;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1946;
wire n_1449;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_3060;
wire n_4276;
wire n_2651;
wire n_3947;
wire n_4358;
wire n_3490;
wire n_3656;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2643;
wire n_1374;
wire n_1328;
wire n_2561;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_3868;
wire n_4369;
wire n_2099;
wire n_2408;
wire n_4168;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_4203;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_4394;
wire n_1723;
wire n_955;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_4350;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_3156;
wire n_550;
wire n_696;
wire n_3101;
wire n_3669;
wire n_897;
wire n_798;
wire n_3376;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_3798;
wire n_3702;
wire n_1040;
wire n_4065;
wire n_3836;
wire n_2202;
wire n_2648;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_578;
wire n_2976;
wire n_3876;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_4135;
wire n_2439;
wire n_1931;
wire n_1218;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_4187;
wire n_1547;
wire n_777;
wire n_1070;
wire n_4166;
wire n_2089;
wire n_3420;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1561;
wire n_1165;
wire n_1267;
wire n_1071;
wire n_496;
wire n_1801;
wire n_3985;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_3361;
wire n_2970;
wire n_2908;
wire n_1600;
wire n_521;
wire n_3744;
wire n_663;
wire n_845;
wire n_2235;
wire n_4263;
wire n_1862;
wire n_673;
wire n_837;
wire n_3980;
wire n_1239;
wire n_2915;
wire n_528;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_4255;
wire n_1587;
wire n_1473;
wire n_680;
wire n_2682;
wire n_553;
wire n_901;
wire n_3755;
wire n_2432;
wire n_3668;
wire n_813;
wire n_4258;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_4237;
wire n_2506;
wire n_675;
wire n_2699;
wire n_4064;
wire n_888;
wire n_1880;
wire n_2769;
wire n_3550;
wire n_2337;
wire n_3436;
wire n_1167;
wire n_1626;
wire n_3542;
wire n_637;
wire n_2615;
wire n_3940;
wire n_1556;
wire n_1384;
wire n_3907;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_3841;
wire n_2238;
wire n_923;
wire n_2118;
wire n_2985;
wire n_691;
wire n_1151;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_4080;
wire n_4006;
wire n_3141;
wire n_4226;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_3986;
wire n_4376;
wire n_3716;
wire n_4025;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_3191;
wire n_1585;
wire n_571;
wire n_2684;
wire n_2712;
wire n_3593;
wire n_3193;
wire n_3837;
wire n_3885;
wire n_1971;
wire n_1599;
wire n_3936;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3507;
wire n_3273;
wire n_3821;
wire n_2713;
wire n_3544;
wire n_2700;
wire n_2644;
wire n_4310;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_4020;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_1447;
wire n_907;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_3915;
wire n_2370;
wire n_3496;
wire n_3954;
wire n_4114;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_3735;
wire n_4067;
wire n_2248;
wire n_4042;
wire n_4176;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_4385;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_3899;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_4159;
wire n_3714;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_4089;
wire n_3651;
wire n_3310;
wire n_3487;
wire n_593;
wire n_4333;
wire n_2258;
wire n_4069;
wire n_748;
wire n_1058;
wire n_586;
wire n_1667;
wire n_3359;
wire n_838;
wire n_2784;
wire n_3718;
wire n_3983;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_3470;
wire n_1224;
wire n_2865;
wire n_4327;
wire n_4405;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_4195;
wire n_953;
wire n_1014;
wire n_4218;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_4375;
wire n_2241;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_3781;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_4246;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_4353;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_534;
wire n_3106;
wire n_1882;
wire n_4164;
wire n_884;
wire n_3328;
wire n_944;
wire n_4130;
wire n_1754;
wire n_4234;
wire n_3889;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_4256;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_4088;
wire n_4224;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_4161;
wire n_647;
wire n_3433;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_3392;
wire n_832;
wire n_857;
wire n_2305;
wire n_3430;
wire n_1072;
wire n_3975;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_1319;
wire n_561;
wire n_2379;
wire n_3447;
wire n_3331;
wire n_2616;
wire n_2911;
wire n_3992;
wire n_3305;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_4148;
wire n_4151;
wire n_1906;
wire n_1883;
wire n_4103;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_3528;
wire n_3649;
wire n_2262;
wire n_4302;
wire n_2462;
wire n_2514;
wire n_4373;
wire n_1532;
wire n_4252;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_4331;
wire n_4160;
wire n_2945;
wire n_2331;
wire n_2798;
wire n_2293;
wire n_686;
wire n_3989;
wire n_2837;
wire n_847;
wire n_3804;
wire n_4051;
wire n_4344;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_4097;
wire n_558;
wire n_3655;
wire n_3009;
wire n_702;
wire n_1276;
wire n_2808;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_3981;
wire n_2108;
wire n_3640;
wire n_728;
wire n_4388;
wire n_2930;
wire n_1162;
wire n_1538;
wire n_4206;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_3602;
wire n_1038;
wire n_2967;
wire n_520;
wire n_1369;
wire n_3909;
wire n_2611;
wire n_4261;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_3944;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_4090;
wire n_809;
wire n_3923;
wire n_931;
wire n_870;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_4001;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_4219;
wire n_868;
wire n_2454;
wire n_4371;
wire n_639;
wire n_2804;
wire n_914;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_3120;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_4007;
wire n_3790;
wire n_4011;
wire n_4268;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_3643;
wire n_3895;
wire n_4194;
wire n_2222;
wire n_1892;
wire n_4120;
wire n_3510;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_4278;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_2690;
wire n_4028;
wire n_4082;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_4085;
wire n_1259;
wire n_4073;
wire n_1690;
wire n_4260;
wire n_3819;
wire n_706;
wire n_746;
wire n_1649;
wire n_3150;
wire n_4163;
wire n_747;
wire n_2064;
wire n_784;
wire n_3978;
wire n_4325;
wire n_2449;
wire n_3867;
wire n_1733;
wire n_4372;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_4186;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_3747;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_3833;
wire n_865;
wire n_2227;
wire n_3775;
wire n_4133;
wire n_678;
wire n_2671;
wire n_697;
wire n_4262;
wire n_4184;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_1798;
wire n_2022;
wire n_776;
wire n_3814;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_4099;
wire n_2592;
wire n_3416;
wire n_4379;
wire n_525;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_4340;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_4295;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_4030;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_4334;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_4397;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_744;
wire n_629;
wire n_590;
wire n_3770;
wire n_4014;
wire n_2631;
wire n_1308;
wire n_3068;
wire n_2178;
wire n_2871;
wire n_1767;
wire n_3144;
wire n_4244;
wire n_2943;
wire n_2913;
wire n_4254;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_4179;
wire n_3469;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_1615;
wire n_4175;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_3317;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_604;
wire n_2007;
wire n_3220;
wire n_4391;
wire n_949;
wire n_2539;
wire n_3917;
wire n_3942;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_3855;
wire n_1539;
wire n_946;
wire n_2736;
wire n_4157;
wire n_4283;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_3765;
wire n_498;
wire n_1468;
wire n_1559;
wire n_3823;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_4173;
wire n_689;
wire n_3158;
wire n_738;
wire n_1624;
wire n_3000;
wire n_640;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_624;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_3113;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_2577;
wire n_3760;
wire n_4108;
wire n_4078;
wire n_1760;
wire n_2875;
wire n_936;
wire n_568;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_757;
wire n_3844;
wire n_3280;
wire n_2342;
wire n_633;
wire n_2856;
wire n_4054;
wire n_3471;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_3205;
wire n_4156;
wire n_2046;
wire n_4146;
wire n_2848;
wire n_2741;
wire n_4360;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3828;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_4404;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_3988;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_1145;
wire n_878;
wire n_524;
wire n_3843;
wire n_3457;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_3856;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_4324;
wire n_1068;
wire n_3030;
wire n_3558;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_4249;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_906;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_4086;
wire n_2412;
wire n_4356;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_724;
wire n_3753;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_658;
wire n_2061;
wire n_3773;
wire n_3555;
wire n_3579;
wire n_3918;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_4317;
wire n_3969;
wire n_2857;
wire n_3932;
wire n_1586;
wire n_4291;
wire n_959;
wire n_2459;
wire n_3031;
wire n_4154;
wire n_535;
wire n_3396;
wire n_3701;
wire n_940;
wire n_4386;
wire n_1445;
wire n_3516;
wire n_4023;
wire n_4149;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1923;
wire n_1773;
wire n_592;
wire n_3243;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_978;
wire n_2768;
wire n_4299;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_4019;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_514;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2473;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_603;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_3767;
wire n_4279;
wire n_4396;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_3820;
wire n_636;
wire n_4367;
wire n_3741;
wire n_660;
wire n_3410;
wire n_2087;
wire n_1640;
wire n_4294;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_750;
wire n_2029;
wire n_742;
wire n_995;
wire n_3221;
wire n_4125;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3629;
wire n_3021;
wire n_4232;
wire n_1989;
wire n_3818;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_4387;
wire n_662;
wire n_2312;
wire n_3990;
wire n_962;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_4170;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_4147;
wire n_4308;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_4365;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_3830;
wire n_1043;
wire n_2585;
wire n_3505;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_3730;
wire n_3883;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_974;
wire n_2565;
wire n_4152;
wire n_727;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_957;
wire n_3787;
wire n_773;
wire n_2124;
wire n_743;
wire n_3001;
wire n_2081;
wire n_3945;
wire n_4392;
wire n_3149;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_4296;
wire n_2418;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_4281;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_4200;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_3614;
wire n_4198;
wire n_2909;
wire n_2111;
wire n_1724;
wire n_2521;
wire n_3301;
wire n_4285;
wire n_3466;
wire n_3458;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_1366;
wire n_1300;
wire n_3960;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2477;
wire n_761;
wire n_2277;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_3905;
wire n_4329;
wire n_1006;
wire n_3411;
wire n_3887;
wire n_4087;
wire n_2110;
wire n_3811;
wire n_4093;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_4271;
wire n_1486;
wire n_582;
wire n_3586;
wire n_1332;
wire n_3519;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_4174;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_512;
wire n_2367;
wire n_2033;
wire n_1591;
wire n_4071;
wire n_4330;
wire n_4341;
wire n_4257;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_3399;
wire n_4312;
wire n_2896;
wire n_652;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_4074;
wire n_1927;
wire n_3065;
wire n_4361;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_3645;
wire n_609;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3838;
wire n_3077;
wire n_3929;
wire n_4277;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_834;
wire n_3474;
wire n_765;
wire n_4140;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_3984;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_3938;
wire n_1913;
wire n_988;
wire n_2878;
wire n_504;
wire n_1823;
wire n_511;
wire n_3679;
wire n_3779;
wire n_874;
wire n_2464;
wire n_3422;
wire n_3888;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_4326;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_4189;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_4110;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_987;
wire n_4207;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_4305;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_3849;
wire n_3946;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_545;
wire n_860;
wire n_3229;
wire n_4213;
wire n_2849;
wire n_1805;
wire n_3925;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_948;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4059;
wire n_2455;
wire n_4349;
wire n_628;
wire n_1849;
wire n_3788;
wire n_4084;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_4313;
wire n_970;
wire n_4037;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_513;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_3421;
wire n_4139;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_4063;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_3242;
wire n_1552;
wire n_2508;
wire n_3592;
wire n_3618;
wire n_4031;
wire n_495;
wire n_602;
wire n_3525;
wire n_574;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_879;
wire n_3394;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_623;
wire n_3995;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_3808;
wire n_824;
wire n_4036;
wire n_1645;
wire n_3881;
wire n_4339;
wire n_4041;
wire n_2461;
wire n_490;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_4060;
wire n_1684;
wire n_921;
wire n_2658;
wire n_3590;
wire n_996;
wire n_1717;
wire n_572;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_4210;
wire n_2578;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_1381;
wire n_2555;
wire n_3751;
wire n_2662;
wire n_2740;
wire n_3824;
wire n_3890;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_4076;
wire n_2554;
wire n_3465;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_1438;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_589;
wire n_3961;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_716;
wire n_3589;
wire n_4102;
wire n_562;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_3658;
wire n_3449;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_3993;
wire n_2216;
wire n_531;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_4230;
wire n_2308;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_3860;
wire n_1382;
wire n_1029;
wire n_925;
wire n_3546;
wire n_1206;
wire n_4248;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_3941;
wire n_3195;
wire n_1519;
wire n_3190;
wire n_950;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_3847;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3893;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_968;
wire n_912;
wire n_3548;
wire n_4348;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_3334;
wire n_967;
wire n_1442;
wire n_2923;
wire n_4162;
wire n_3665;
wire n_4355;
wire n_3494;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_515;
wire n_2333;
wire n_3953;
wire n_885;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_3875;
wire n_3976;
wire n_4122;
wire n_1357;
wire n_2125;
wire n_3771;
wire n_3979;
wire n_4297;
wire n_683;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_4003;
wire n_3800;
wire n_721;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_4301;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_4048;
wire n_4026;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_983;
wire n_1844;
wire n_4104;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_4377;
wire n_1305;
wire n_3749;
wire n_3178;
wire n_873;
wire n_1826;
wire n_3962;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1283;
wire n_1644;
wire n_762;
wire n_4172;
wire n_2334;
wire n_2637;
wire n_4384;
wire n_3695;
wire n_690;
wire n_4046;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_3537;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_4096;
wire n_4199;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_821;
wire n_3816;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_4286;
wire n_3864;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_507;
wire n_2269;
wire n_2732;
wire n_3569;
wire n_2415;
wire n_2309;
wire n_2948;
wire n_3274;
wire n_3041;
wire n_3299;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_4362;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_972;
wire n_3504;
wire n_692;
wire n_2037;
wire n_2685;
wire n_3920;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_3737;
wire n_3913;
wire n_1185;
wire n_991;
wire n_2903;
wire n_3417;
wire n_3482;
wire n_3866;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_3717;
wire n_4106;
wire n_4034;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_945;
wire n_2997;
wire n_492;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_4400;
wire n_943;
wire n_3326;
wire n_3956;
wire n_3572;
wire n_992;
wire n_3067;
wire n_4215;
wire n_1932;
wire n_4280;
wire n_3375;
wire n_2755;
wire n_4047;
wire n_543;
wire n_842;
wire n_3734;
wire n_650;
wire n_984;
wire n_694;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_4402;
wire n_3167;
wire n_4239;
wire n_4029;
wire n_3400;
wire n_1594;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_3423;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_3870;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_4352;
wire n_918;
wire n_3529;
wire n_3854;
wire n_2169;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_4201;
wire n_1610;
wire n_4347;
wire n_1077;
wire n_1422;
wire n_3196;
wire n_4095;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_4338;
wire n_540;
wire n_3492;
wire n_618;
wire n_3094;
wire n_896;
wire n_2310;
wire n_2780;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_4043;
wire n_3704;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_4027;
wire n_831;
wire n_2280;
wire n_4123;
wire n_2192;
wire n_964;
wire n_3633;
wire n_3363;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1735;
wire n_1575;
wire n_1697;
wire n_833;
wire n_2393;
wire n_2318;
wire n_3689;
wire n_2020;
wire n_3831;
wire n_1646;
wire n_2502;
wire n_3801;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_2749;
wire n_3372;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2751;
wire n_2707;
wire n_2793;
wire n_3451;
wire n_2971;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3950;
wire n_4000;
wire n_655;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_4121;
wire n_3998;
wire n_1446;
wire n_2285;
wire n_4406;
wire n_3147;
wire n_2758;
wire n_4141;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_3869;
wire n_4307;
wire n_1149;
wire n_2618;
wire n_4359;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_3230;
wire n_1020;
wire n_1062;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_3931;
wire n_3708;
wire n_1204;
wire n_4010;
wire n_4107;
wire n_2840;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_3861;
wire n_3780;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_4117;
wire n_2893;
wire n_3636;
wire n_1188;
wire n_2962;
wire n_2588;
wire n_4004;
wire n_4118;
wire n_1722;
wire n_3957;
wire n_661;
wire n_2441;
wire n_3848;
wire n_1802;
wire n_3083;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_4079;
wire n_3898;
wire n_849;
wire n_2795;
wire n_4091;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_510;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3829;
wire n_3380;
wire n_3177;
wire n_4053;
wire n_830;
wire n_4274;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3409;
wire n_3460;
wire n_2352;
wire n_3538;
wire n_1413;
wire n_801;
wire n_4040;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_749;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_4316;
wire n_939;
wire n_3697;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_3393;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_4247;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_4018;
wire n_4044;
wire n_3900;
wire n_4062;
wire n_4113;
wire n_3520;
wire n_3971;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_3759;
wire n_1338;
wire n_577;
wire n_4005;
wire n_2016;
wire n_1522;
wire n_4321;
wire n_4342;
wire n_3872;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_4336;
wire n_3933;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_3578;
wire n_3966;
wire n_836;
wire n_990;
wire n_2867;
wire n_3812;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_3145;
wire n_4183;
wire n_3124;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4253;
wire n_4290;
wire n_4233;
wire n_3192;
wire n_2608;
wire n_3877;
wire n_3764;
wire n_2657;
wire n_770;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_3547;
wire n_2649;
wire n_3977;
wire n_1102;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_4052;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_711;
wire n_1499;
wire n_3061;
wire n_4398;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1834;
wire n_2097;
wire n_1659;
wire n_2313;
wire n_2542;
wire n_489;
wire n_1174;
wire n_2431;
wire n_3324;
wire n_3356;
wire n_3758;
wire n_2835;
wire n_3914;
wire n_4304;
wire n_3911;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3803;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_4192;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_3736;
wire n_1190;
wire n_3506;
wire n_3896;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_3958;
wire n_2409;
wire n_601;
wire n_917;
wire n_3450;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_4115;
wire n_726;
wire n_3174;
wire n_982;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_3746;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_3817;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_3408;
wire n_1904;
wire n_4167;
wire n_2640;
wire n_1993;
wire n_774;
wire n_3835;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1514;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_1345;
wire n_1059;
wire n_3967;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_3090;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_3762;
wire n_3902;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_4070;
wire n_2148;
wire n_4282;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_4180;
wire n_1584;
wire n_1726;
wire n_665;
wire n_1835;
wire n_3035;
wire n_3654;
wire n_1440;
wire n_3839;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_4143;
wire n_4323;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_3972;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_3639;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4105;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_3791;
wire n_4204;
wire n_3308;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_2224;
wire n_1979;
wire n_791;
wire n_1991;
wire n_1533;
wire n_732;
wire n_3368;
wire n_2924;
wire n_3467;
wire n_808;
wire n_2484;
wire n_4111;
wire n_797;
wire n_3530;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_4322;
wire n_500;
wire n_2994;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_4354;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_766;
wire n_3928;
wire n_541;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_3534;
wire n_715;
wire n_3901;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3757;
wire n_536;
wire n_3438;
wire n_4098;
wire n_872;
wire n_2012;
wire n_594;
wire n_3792;
wire n_4272;
wire n_1291;
wire n_3974;
wire n_3381;
wire n_3871;
wire n_4094;
wire n_3503;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_4269;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_2965;
wire n_3536;
wire n_3661;
wire n_3635;
wire n_4150;
wire n_827;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_1703;
wire n_3312;
wire n_4055;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_1144;
wire n_3973;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_3882;
wire n_3934;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_3826;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_3922;
wire n_3846;
wire n_676;
wire n_2103;
wire n_653;
wire n_3968;
wire n_2160;
wire n_642;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_4017;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_3943;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_4072;
wire n_916;
wire n_1081;
wire n_2549;
wire n_493;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_4380;
wire n_980;
wire n_1115;
wire n_698;
wire n_703;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_4022;
wire n_998;
wire n_3802;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_3600;
wire n_501;
wire n_823;
wire n_2686;
wire n_2528;
wire n_4134;
wire n_725;
wire n_2344;
wire n_3892;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_4035;
wire n_2316;
wire n_672;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_3315;
wire n_581;
wire n_2906;
wire n_554;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_3172;
wire n_3139;
wire n_2773;
wire n_3292;
wire n_3239;
wire n_2598;
wire n_3878;
wire n_1762;
wire n_1013;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_718;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_2850;
wire n_1747;
wire n_714;
wire n_4220;
wire n_4251;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_4075;
wire n_4193;
wire n_3982;
wire n_2654;
wire n_997;
wire n_3431;
wire n_3104;
wire n_932;
wire n_3169;
wire n_3151;
wire n_612;
wire n_3822;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_3850;
wire n_788;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_4066;
wire n_3647;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_559;
wire n_825;
wire n_4351;
wire n_2819;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_4368;
wire n_737;
wire n_1718;
wire n_4050;
wire n_3700;
wire n_3609;
wire n_4136;
wire n_986;
wire n_2315;
wire n_509;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_4077;
wire n_4223;
wire n_4393;
wire n_1192;
wire n_2221;
wire n_3576;
wire n_1024;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_733;
wire n_1922;
wire n_2966;
wire n_4049;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_3862;
wire n_1569;
wire n_2188;
wire n_3495;
wire n_3879;
wire n_867;
wire n_2348;
wire n_2422;
wire n_3959;
wire n_2239;
wire n_587;
wire n_2950;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_4346;
wire n_3852;
wire n_548;
wire n_3170;
wire n_3724;
wire n_812;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_518;
wire n_505;
wire n_2057;
wire n_3272;
wire n_4008;
wire n_3011;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_4196;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_862;
wire n_3584;
wire n_1425;
wire n_760;
wire n_3858;
wire n_1901;
wire n_3069;
wire n_3756;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_2889;
wire n_3691;
wire n_4235;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_4382;
wire n_2939;
wire n_1745;
wire n_3924;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_3999;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_3807;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2447;
wire n_1813;
wire n_2343;
wire n_3761;
wire n_886;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_654;
wire n_1172;
wire n_2535;
wire n_4205;
wire n_1341;
wire n_2774;
wire n_570;
wire n_2726;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_853;
wire n_4178;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_751;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_4229;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_704;
wire n_787;
wire n_4399;
wire n_1770;
wire n_2781;
wire n_4100;
wire n_4228;
wire n_2456;
wire n_4401;
wire n_3904;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_522;
wire n_3364;
wire n_1287;
wire n_4363;
wire n_1262;
wire n_2691;
wire n_930;
wire n_4092;
wire n_3908;
wire n_1873;
wire n_1411;
wire n_3926;
wire n_3201;
wire n_3054;
wire n_4335;
wire n_1962;
wire n_622;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_4181;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_4225;
wire n_3391;
wire n_682;
wire n_1567;
wire n_4259;
wire n_2567;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_922;
wire n_3122;
wire n_816;
wire n_1648;
wire n_4015;
wire n_591;
wire n_3842;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_4056;
wire n_4153;
wire n_1344;
wire n_2041;
wire n_631;
wire n_3627;
wire n_1246;
wire n_3840;
wire n_4300;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_2957;
wire n_839;
wire n_3551;
wire n_3903;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_4267;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_3865;
wire n_3722;
wire n_3859;
wire n_4171;
wire n_1842;
wire n_871;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_4045;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_772;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_499;
wire n_2531;
wire n_1589;
wire n_4116;
wire n_517;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_3754;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_3115;
wire n_4287;
wire n_3509;
wire n_3352;
wire n_4390;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_4182;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_3251;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_3955;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_3794;
wire n_2050;
wire n_2809;
wire n_4270;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_1277;
wire n_722;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_844;
wire n_3384;
wire n_852;
wire n_3497;
wire n_1487;
wire n_1864;
wire n_3644;
wire n_1028;
wire n_1601;
wire n_4016;
wire n_3336;
wire n_3935;
wire n_781;
wire n_2940;
wire n_542;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_595;
wire n_502;
wire n_3562;
wire n_3948;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_4231;
wire n_979;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3322;
wire n_3232;
wire n_3652;
wire n_1245;
wire n_846;
wire n_2505;
wire n_2438;
wire n_2427;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_4061;
wire n_2296;
wire n_2070;
wire n_3250;
wire n_1937;
wire n_585;
wire n_2112;
wire n_4083;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_616;
wire n_2278;
wire n_2594;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3234;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_4328;
wire n_3004;
wire n_3323;
wire n_3916;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_3921;
wire n_4081;
wire n_3132;
wire n_3556;
wire n_648;
wire n_1379;
wire n_2734;
wire n_3874;
wire n_4101;
wire n_4407;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3951;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_494;
wire n_1761;
wire n_641;
wire n_3238;
wire n_3210;
wire n_4389;
wire n_3930;
wire n_730;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_575;
wire n_795;
wire n_2404;
wire n_4345;
wire n_2083;
wire n_695;
wire n_3281;
wire n_656;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3964;
wire n_3266;
wire n_2485;
wire n_4318;
wire n_3772;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_3884;
wire n_4185;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_3726;
wire n_2210;
wire n_4169;
wire n_805;
wire n_3247;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_4032;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_4319;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_657;
wire n_4320;
wire n_644;
wire n_1741;
wire n_2229;
wire n_4124;
wire n_1160;
wire n_1397;
wire n_4057;
wire n_4332;
wire n_491;
wire n_1258;
wire n_4314;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_3809;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_3694;
wire n_1448;
wire n_4288;
wire n_4245;
wire n_4364;
wire n_2225;
wire n_3567;
wire n_3613;
wire n_1507;
wire n_4378;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_597;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_3853;
wire n_1181;
wire n_1505;
wire n_4222;
wire n_4216;
wire n_1634;
wire n_3939;
wire n_1196;
wire n_4012;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_811;
wire n_1558;
wire n_3225;
wire n_4241;
wire n_807;
wire n_3321;
wire n_2166;
wire n_3910;
wire n_2938;
wire n_3212;
wire n_835;
wire n_666;
wire n_3319;
wire n_3594;
wire n_1433;
wire n_4309;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_1254;
wire n_3799;
wire n_4119;
wire n_4298;
wire n_1026;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_2044;
wire n_927;
wire n_1089;
wire n_2013;
wire n_2689;
wire n_1990;
wire n_2920;
wire n_3259;
wire n_4265;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_4191;
wire n_2511;
wire n_4293;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_3016;
wire n_2894;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_4188;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_4214;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1180;
wire n_1827;
wire n_3360;
wire n_4209;
wire n_2524;
wire n_3873;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_533;
wire n_1542;
wire n_1251;
wire n_3693;
wire n_4366;
wire n_4009;
wire n_3159;
wire n_2728;
wire n_3857;
wire n_2268;
wire n_3778;

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_313),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_388),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_431),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_201),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_305),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_387),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_57),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_465),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_182),
.Y(n_496)
);

BUFx2_ASAP7_75t_SL g497 ( 
.A(n_243),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_175),
.Y(n_498)
);

BUFx10_ASAP7_75t_L g499 ( 
.A(n_38),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_333),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_55),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_188),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_285),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_296),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_305),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_402),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_31),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_142),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_348),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_75),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_386),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_146),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_463),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_26),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_179),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_95),
.Y(n_516)
);

BUFx10_ASAP7_75t_L g517 ( 
.A(n_78),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_404),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_423),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_234),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_454),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_365),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_287),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_41),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_269),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_66),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_6),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_470),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_168),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_107),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_153),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_158),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_240),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_228),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_419),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_479),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_134),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_168),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_201),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_212),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_450),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_6),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_0),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_214),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_257),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_35),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_442),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_173),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_331),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_197),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_333),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_247),
.Y(n_552)
);

BUFx10_ASAP7_75t_L g553 ( 
.A(n_426),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_109),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_58),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_260),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_477),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_427),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_466),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_164),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_279),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_360),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_143),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_252),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_9),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_25),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_160),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_420),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_374),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_29),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_137),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_435),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_344),
.Y(n_573)
);

CKINVDCx14_ASAP7_75t_R g574 ( 
.A(n_298),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_169),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_31),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_379),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_249),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_365),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_57),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_190),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_152),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_405),
.Y(n_583)
);

BUFx10_ASAP7_75t_L g584 ( 
.A(n_248),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_392),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_224),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_396),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_395),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_203),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_27),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_29),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_283),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_336),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_421),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_416),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_403),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_215),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_87),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_156),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_82),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_481),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_115),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_66),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_363),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_343),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_171),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_26),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_474),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_89),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_90),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_255),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_249),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_85),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_101),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_385),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_476),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_200),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_480),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_5),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_92),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_456),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_81),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_282),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_334),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_376),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_349),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_182),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_452),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_145),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_432),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_32),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_177),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_309),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_180),
.Y(n_634)
);

CKINVDCx16_ASAP7_75t_R g635 ( 
.A(n_233),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_181),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_223),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_227),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_246),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_13),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_151),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_118),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_214),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_358),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_243),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_225),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_206),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_213),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_337),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_457),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_225),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_106),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_281),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_319),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_218),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_334),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_487),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_384),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_162),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_455),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_78),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_297),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_446),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_441),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_282),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_49),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_272),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_215),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_371),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_98),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_122),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_235),
.Y(n_672)
);

INVxp67_ASAP7_75t_SL g673 ( 
.A(n_80),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_202),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_406),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_352),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_257),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_169),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_153),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_245),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_180),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_67),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_335),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_82),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_253),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_336),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_331),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_253),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_332),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_398),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_106),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_445),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_461),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_358),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_323),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_429),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_323),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_317),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_280),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_459),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_472),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_458),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_107),
.Y(n_703)
);

BUFx10_ASAP7_75t_L g704 ( 
.A(n_129),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_96),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_399),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_219),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_204),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_81),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_352),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_71),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_251),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_341),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_231),
.Y(n_714)
);

BUFx5_ASAP7_75t_L g715 ( 
.A(n_179),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_307),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_138),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_102),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_200),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_284),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_15),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_255),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_104),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_252),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_103),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_30),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_350),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_156),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_368),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_90),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_413),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_283),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_17),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_324),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_47),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_237),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_400),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_32),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_145),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_335),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_60),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_165),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_22),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_451),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_438),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_343),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_23),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_94),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_380),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_326),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_484),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_486),
.Y(n_752)
);

BUFx10_ASAP7_75t_L g753 ( 
.A(n_286),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_259),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_202),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_16),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_322),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_341),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_482),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_121),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_195),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_30),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_3),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_475),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_241),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_112),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_210),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_293),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_275),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_22),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_97),
.Y(n_771)
);

HB1xp67_ASAP7_75t_SL g772 ( 
.A(n_49),
.Y(n_772)
);

BUFx2_ASAP7_75t_R g773 ( 
.A(n_372),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_197),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_473),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_370),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_393),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_232),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_27),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_270),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_2),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_322),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_91),
.Y(n_783)
);

CKINVDCx14_ASAP7_75t_R g784 ( 
.A(n_389),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_183),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_375),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_79),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_428),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_209),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_150),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_4),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_284),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_167),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_84),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_55),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_715),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_574),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_715),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_715),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_545),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_541),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_503),
.Y(n_802)
);

INVxp33_ASAP7_75t_L g803 ( 
.A(n_503),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_715),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_715),
.Y(n_805)
);

INVxp67_ASAP7_75t_SL g806 ( 
.A(n_596),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_596),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_715),
.Y(n_808)
);

INVxp33_ASAP7_75t_SL g809 ( 
.A(n_694),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_694),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_715),
.Y(n_811)
);

INVxp33_ASAP7_75t_SL g812 ( 
.A(n_497),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_715),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_715),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_545),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_542),
.Y(n_816)
);

INVxp67_ASAP7_75t_SL g817 ( 
.A(n_669),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_542),
.Y(n_818)
);

NOR2xp67_ASAP7_75t_L g819 ( 
.A(n_491),
.B(n_0),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_542),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_669),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_542),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_542),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_569),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_542),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_552),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_552),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_650),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_635),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_518),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_552),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_552),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_675),
.Y(n_833)
);

CKINVDCx16_ASAP7_75t_R g834 ( 
.A(n_635),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_552),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_540),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_552),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_570),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_669),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_570),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_570),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_570),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_570),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_570),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_670),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_670),
.Y(n_846)
);

INVxp33_ASAP7_75t_L g847 ( 
.A(n_772),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_670),
.Y(n_848)
);

INVxp67_ASAP7_75t_SL g849 ( 
.A(n_670),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_670),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_497),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_494),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_711),
.Y(n_853)
);

BUFx5_ASAP7_75t_L g854 ( 
.A(n_495),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_495),
.Y(n_855)
);

INVxp67_ASAP7_75t_SL g856 ( 
.A(n_670),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_513),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_513),
.Y(n_858)
);

CKINVDCx16_ASAP7_75t_R g859 ( 
.A(n_711),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_777),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_488),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_494),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_536),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_734),
.Y(n_864)
);

INVxp33_ASAP7_75t_SL g865 ( 
.A(n_492),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_536),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_568),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_568),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_572),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_572),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_511),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_496),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_585),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_585),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_498),
.Y(n_875)
);

CKINVDCx14_ASAP7_75t_R g876 ( 
.A(n_784),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_511),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_587),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_587),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_588),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_588),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_608),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_608),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_489),
.Y(n_884)
);

CKINVDCx16_ASAP7_75t_R g885 ( 
.A(n_499),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_504),
.Y(n_886)
);

INVxp67_ASAP7_75t_SL g887 ( 
.A(n_734),
.Y(n_887)
);

CKINVDCx16_ASAP7_75t_R g888 ( 
.A(n_499),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_490),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_493),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_615),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_615),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_616),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_616),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_663),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_505),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_507),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_663),
.Y(n_898)
);

CKINVDCx16_ASAP7_75t_R g899 ( 
.A(n_499),
.Y(n_899)
);

CKINVDCx16_ASAP7_75t_R g900 ( 
.A(n_499),
.Y(n_900)
);

INVxp33_ASAP7_75t_SL g901 ( 
.A(n_508),
.Y(n_901)
);

INVxp33_ASAP7_75t_L g902 ( 
.A(n_500),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_664),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_734),
.Y(n_904)
);

CKINVDCx16_ASAP7_75t_R g905 ( 
.A(n_517),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_664),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_692),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_692),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_540),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_509),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_701),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_701),
.Y(n_912)
);

CKINVDCx14_ASAP7_75t_R g913 ( 
.A(n_517),
.Y(n_913)
);

NOR2xp67_ASAP7_75t_L g914 ( 
.A(n_491),
.B(n_1),
.Y(n_914)
);

INVxp33_ASAP7_75t_L g915 ( 
.A(n_500),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_506),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_702),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_502),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_702),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_521),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_749),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_749),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_734),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_734),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_734),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_771),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_528),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_514),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_771),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_751),
.B(n_1),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_518),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_771),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_553),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_515),
.Y(n_934)
);

INVxp33_ASAP7_75t_SL g935 ( 
.A(n_520),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_771),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_771),
.Y(n_937)
);

INVxp67_ASAP7_75t_SL g938 ( 
.A(n_771),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_512),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_512),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_535),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_539),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_539),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_631),
.Y(n_944)
);

INVxp33_ASAP7_75t_L g945 ( 
.A(n_510),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_631),
.Y(n_946)
);

BUFx2_ASAP7_75t_SL g947 ( 
.A(n_556),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_830),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_830),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_800),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_818),
.Y(n_951)
);

OAI22x1_ASAP7_75t_SL g952 ( 
.A1(n_809),
.A2(n_543),
.B1(n_554),
.B2(n_529),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_821),
.Y(n_953)
);

INVx5_ASAP7_75t_L g954 ( 
.A(n_830),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_830),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_816),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_830),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_816),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_800),
.Y(n_959)
);

BUFx8_ASAP7_75t_SL g960 ( 
.A(n_871),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_818),
.Y(n_961)
);

OAI22x1_ASAP7_75t_R g962 ( 
.A1(n_877),
.A2(n_613),
.B1(n_629),
.B2(n_610),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_808),
.A2(n_621),
.B(n_751),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_817),
.B(n_540),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_931),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_841),
.B(n_621),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_864),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_815),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_849),
.B(n_759),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_931),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_SL g971 ( 
.A1(n_809),
.A2(n_666),
.B1(n_680),
.B2(n_634),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_820),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_931),
.Y(n_973)
);

CKINVDCx16_ASAP7_75t_R g974 ( 
.A(n_834),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_806),
.B(n_807),
.Y(n_975)
);

BUFx12f_ASAP7_75t_L g976 ( 
.A(n_797),
.Y(n_976)
);

BUFx8_ASAP7_75t_L g977 ( 
.A(n_836),
.Y(n_977)
);

INVx6_ASAP7_75t_L g978 ( 
.A(n_931),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_931),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_808),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_821),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_815),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_829),
.Y(n_983)
);

AOI22x1_ASAP7_75t_SL g984 ( 
.A1(n_801),
.A2(n_720),
.B1(n_727),
.B2(n_686),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_820),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_864),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_856),
.B(n_759),
.Y(n_987)
);

INVx5_ASAP7_75t_L g988 ( 
.A(n_904),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_933),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_822),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_853),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_904),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_839),
.B(n_547),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_876),
.B(n_557),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_822),
.Y(n_995)
);

INVx6_ASAP7_75t_L g996 ( 
.A(n_854),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_933),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_823),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_887),
.B(n_764),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_823),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_825),
.Y(n_1001)
);

AOI22x1_ASAP7_75t_SL g1002 ( 
.A1(n_824),
.A2(n_756),
.B1(n_782),
.B2(n_735),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_853),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_825),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_861),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_859),
.A2(n_791),
.B1(n_789),
.B2(n_555),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_826),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_826),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_827),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_827),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_831),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_831),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_798),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_832),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_861),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_832),
.Y(n_1016)
);

OA21x2_ASAP7_75t_L g1017 ( 
.A1(n_835),
.A2(n_788),
.B(n_764),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_835),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_837),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_836),
.B(n_682),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_837),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_838),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_909),
.B(n_682),
.Y(n_1023)
);

INVx6_ASAP7_75t_L g1024 ( 
.A(n_854),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_838),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_SL g1026 ( 
.A1(n_918),
.A2(n_614),
.B1(n_668),
.B2(n_501),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_840),
.Y(n_1027)
);

OAI22x1_ASAP7_75t_SL g1028 ( 
.A1(n_812),
.A2(n_523),
.B1(n_533),
.B2(n_527),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_840),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_938),
.B(n_788),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_842),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_797),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_842),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_843),
.Y(n_1034)
);

INVxp67_ASAP7_75t_L g1035 ( 
.A(n_872),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_843),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_844),
.Y(n_1037)
);

BUFx12f_ASAP7_75t_L g1038 ( 
.A(n_875),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_844),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_854),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_845),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_854),
.Y(n_1042)
);

OA21x2_ASAP7_75t_L g1043 ( 
.A1(n_845),
.A2(n_787),
.B(n_783),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_865),
.B(n_752),
.Y(n_1044)
);

AOI22x1_ASAP7_75t_SL g1045 ( 
.A1(n_828),
.A2(n_730),
.B1(n_781),
.B2(n_689),
.Y(n_1045)
);

BUFx12f_ASAP7_75t_L g1046 ( 
.A(n_875),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_909),
.B(n_682),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_855),
.B(n_519),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_857),
.B(n_518),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_846),
.Y(n_1050)
);

BUFx12f_ASAP7_75t_L g1051 ( 
.A(n_886),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_846),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_848),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_884),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_848),
.Y(n_1055)
);

AND2x6_ASAP7_75t_L g1056 ( 
.A(n_798),
.B(n_518),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_897),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_854),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_850),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_886),
.Y(n_1060)
);

BUFx8_ASAP7_75t_L g1061 ( 
.A(n_913),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_850),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_SL g1063 ( 
.A1(n_833),
.A2(n_523),
.B1(n_527),
.B2(n_510),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_851),
.B(n_558),
.Y(n_1064)
);

OAI22x1_ASAP7_75t_R g1065 ( 
.A1(n_860),
.A2(n_524),
.B1(n_525),
.B2(n_522),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_923),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_858),
.B(n_775),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_928),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_863),
.B(n_775),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_923),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_924),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_924),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1013),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_965),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_953),
.B(n_925),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1018),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_960),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1018),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1018),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1013),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1013),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_1043),
.B(n_518),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_953),
.B(n_925),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_965),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_993),
.B(n_975),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_964),
.B(n_947),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_1054),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_1038),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_974),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_964),
.B(n_1020),
.Y(n_1090)
);

BUFx8_ASAP7_75t_L g1091 ( 
.A(n_976),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1013),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_951),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_965),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_951),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1020),
.B(n_947),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_974),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_R g1098 ( 
.A(n_1061),
.B(n_889),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_966),
.B(n_926),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1038),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_956),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_966),
.B(n_926),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_1046),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_961),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_1046),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_956),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_965),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_1051),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_965),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_973),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_1051),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_961),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_973),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_976),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_1061),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_972),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_973),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1061),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_973),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_966),
.B(n_929),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_966),
.B(n_929),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_973),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_981),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1061),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_972),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_958),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_981),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_985),
.Y(n_1128)
);

NOR2xp67_ASAP7_75t_L g1129 ( 
.A(n_1005),
.B(n_896),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_958),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_985),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_967),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_990),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_977),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_SL g1135 ( 
.A1(n_971),
.A2(n_888),
.B1(n_899),
.B2(n_885),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_977),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_967),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1023),
.B(n_847),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_963),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_977),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_981),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_963),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_990),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_977),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_948),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_948),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_992),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1032),
.Y(n_1148)
);

OA21x2_ASAP7_75t_L g1149 ( 
.A1(n_1004),
.A2(n_804),
.B(n_796),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1004),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_1023),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_1032),
.Y(n_1152)
);

NAND2x1p5_ASAP7_75t_L g1153 ( 
.A(n_1043),
.B(n_518),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_984),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_992),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1007),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_969),
.B(n_866),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1007),
.Y(n_1158)
);

INVxp67_ASAP7_75t_SL g1159 ( 
.A(n_970),
.Y(n_1159)
);

CKINVDCx16_ASAP7_75t_R g1160 ( 
.A(n_962),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1008),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1047),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_984),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1008),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_1015),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1002),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1019),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1002),
.Y(n_1168)
);

NAND2xp33_ASAP7_75t_R g1169 ( 
.A(n_950),
.B(n_896),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_950),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_982),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_982),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_1060),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1019),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1022),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1022),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1044),
.B(n_865),
.Y(n_1177)
);

OA21x2_ASAP7_75t_L g1178 ( 
.A1(n_1027),
.A2(n_805),
.B(n_799),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1047),
.Y(n_1179)
);

CKINVDCx16_ASAP7_75t_R g1180 ( 
.A(n_962),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1017),
.A2(n_811),
.B(n_799),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_991),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_991),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_952),
.Y(n_1184)
);

CKINVDCx16_ASAP7_75t_R g1185 ( 
.A(n_1065),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1027),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_983),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_969),
.B(n_932),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_959),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1029),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1029),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_952),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1031),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1068),
.B(n_900),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_995),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_968),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_995),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_969),
.B(n_867),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_948),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1031),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_948),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_948),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1048),
.B(n_868),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_948),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1034),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1003),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_998),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_998),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_971),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_1045),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1034),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1000),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1000),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1045),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1036),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1006),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1006),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_949),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1036),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1035),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1017),
.A2(n_813),
.B(n_811),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1048),
.B(n_869),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1057),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_1065),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1037),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1037),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_949),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1064),
.B(n_901),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1041),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1010),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1041),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1026),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1026),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1068),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_989),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_969),
.B(n_932),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1010),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_989),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1050),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1050),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_997),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_994),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_987),
.B(n_870),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_997),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1063),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1052),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1011),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_949),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1048),
.B(n_873),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1011),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1052),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_987),
.B(n_936),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_R g1253 ( 
.A(n_987),
.B(n_890),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1063),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_949),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1066),
.Y(n_1256)
);

NOR2xp67_ASAP7_75t_L g1257 ( 
.A(n_980),
.B(n_910),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1012),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_987),
.B(n_936),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1066),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1001),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1001),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1001),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_999),
.B(n_937),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1028),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1028),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_R g1267 ( 
.A(n_999),
.B(n_916),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1048),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1001),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_999),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_949),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_999),
.B(n_874),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1030),
.B(n_937),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1012),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1001),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1016),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1014),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1016),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_SL g1279 ( 
.A(n_1030),
.B(n_773),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1030),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1030),
.B(n_878),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1049),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_980),
.B(n_854),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1049),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1043),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1014),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1021),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1016),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_949),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_SL g1290 ( 
.A(n_1049),
.B(n_920),
.Y(n_1290)
);

NAND3xp33_ASAP7_75t_L g1291 ( 
.A(n_1043),
.B(n_934),
.C(n_910),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1016),
.Y(n_1292)
);

INVxp67_ASAP7_75t_L g1293 ( 
.A(n_1049),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1067),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1067),
.B(n_879),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1067),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1021),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1025),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1025),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1225),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1284),
.B(n_1067),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1085),
.B(n_1069),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1187),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1225),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1178),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1178),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1178),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1177),
.B(n_1234),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1073),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1228),
.B(n_1238),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1073),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1285),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1074),
.Y(n_1313)
);

NAND2xp33_ASAP7_75t_L g1314 ( 
.A(n_1270),
.B(n_775),
.Y(n_1314)
);

CKINVDCx6p67_ASAP7_75t_R g1315 ( 
.A(n_1115),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1086),
.B(n_1069),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1270),
.A2(n_1280),
.B1(n_1294),
.B2(n_1282),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1285),
.Y(n_1318)
);

NOR2x1_ASAP7_75t_L g1319 ( 
.A(n_1291),
.B(n_927),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1195),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_1086),
.B(n_905),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1178),
.Y(n_1322)
);

OR2x6_ASAP7_75t_L g1323 ( 
.A(n_1090),
.B(n_556),
.Y(n_1323)
);

INVx2_ASAP7_75t_SL g1324 ( 
.A(n_1096),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1096),
.B(n_1280),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1149),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1090),
.B(n_1069),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1138),
.B(n_803),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1238),
.B(n_941),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1149),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1157),
.B(n_1069),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1149),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1187),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1149),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1157),
.B(n_980),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1195),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1299),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1299),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1197),
.Y(n_1339)
);

INVx4_ASAP7_75t_L g1340 ( 
.A(n_1074),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1139),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1101),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1290),
.A2(n_934),
.B1(n_812),
.B2(n_810),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1298),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1241),
.B(n_901),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1138),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1197),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1203),
.B(n_802),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1157),
.A2(n_930),
.B1(n_1017),
.B2(n_854),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1162),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1162),
.Y(n_1351)
);

INVx4_ASAP7_75t_L g1352 ( 
.A(n_1074),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1203),
.B(n_902),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1198),
.A2(n_1017),
.B1(n_854),
.B2(n_1056),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1241),
.B(n_1244),
.Y(n_1355)
);

OR2x6_ASAP7_75t_L g1356 ( 
.A(n_1179),
.B(n_640),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1222),
.B(n_915),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1198),
.B(n_980),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1101),
.Y(n_1359)
);

INVx5_ASAP7_75t_L g1360 ( 
.A(n_1146),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1106),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1106),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1244),
.B(n_935),
.Y(n_1363)
);

INVxp67_ASAP7_75t_SL g1364 ( 
.A(n_1127),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1126),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1179),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1223),
.B(n_935),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1123),
.B(n_945),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1126),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1198),
.A2(n_1056),
.B1(n_819),
.B2(n_914),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1139),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1279),
.A2(n_673),
.B1(n_640),
.B2(n_671),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1243),
.B(n_1040),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1151),
.B(n_852),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1123),
.B(n_526),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1141),
.B(n_530),
.Y(n_1376)
);

INVx4_ASAP7_75t_L g1377 ( 
.A(n_1074),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1268),
.B(n_559),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1298),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_1089),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1130),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1222),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1130),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1243),
.B(n_1040),
.Y(n_1384)
);

INVx4_ASAP7_75t_L g1385 ( 
.A(n_1074),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1142),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1146),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1243),
.B(n_1040),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1132),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1132),
.Y(n_1390)
);

NAND2xp33_ASAP7_75t_SL g1391 ( 
.A(n_1253),
.B(n_544),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1141),
.B(n_531),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1137),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1137),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1235),
.B(n_1194),
.Y(n_1395)
);

INVx4_ASAP7_75t_L g1396 ( 
.A(n_1084),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1249),
.Y(n_1397)
);

INVx5_ASAP7_75t_L g1398 ( 
.A(n_1146),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_SL g1399 ( 
.A1(n_1216),
.A2(n_553),
.B1(n_517),
.B2(n_550),
.Y(n_1399)
);

INVx6_ASAP7_75t_L g1400 ( 
.A(n_1272),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1249),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1207),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1268),
.B(n_532),
.Y(n_1403)
);

BUFx4f_ASAP7_75t_L g1404 ( 
.A(n_1272),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1297),
.Y(n_1405)
);

AOI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1142),
.A2(n_814),
.B(n_813),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1272),
.A2(n_1281),
.B1(n_1295),
.B2(n_1236),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1147),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1257),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1147),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1216),
.A2(n_553),
.B1(n_517),
.B2(n_550),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1297),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1155),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1242),
.B(n_537),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1207),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1155),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1208),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1267),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1208),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1282),
.A2(n_577),
.B1(n_594),
.B2(n_583),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1077),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1281),
.B(n_862),
.Y(n_1422)
);

INVxp67_ASAP7_75t_SL g1423 ( 
.A(n_1099),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1281),
.B(n_595),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1295),
.A2(n_1056),
.B1(n_775),
.B2(n_814),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1212),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1212),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1213),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1213),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1188),
.A2(n_1056),
.B1(n_775),
.B2(n_671),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1146),
.Y(n_1431)
);

INVx4_ASAP7_75t_L g1432 ( 
.A(n_1084),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1169),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1077),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1230),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1230),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1237),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1293),
.B(n_880),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1237),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1247),
.Y(n_1440)
);

OR2x6_ASAP7_75t_L g1441 ( 
.A(n_1129),
.B(n_644),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1076),
.B(n_1040),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1098),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1078),
.B(n_1042),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1079),
.B(n_1042),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1247),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1250),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1252),
.A2(n_1056),
.B1(n_775),
.B2(n_709),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1259),
.A2(n_1056),
.B1(n_709),
.B2(n_736),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1097),
.Y(n_1450)
);

INVxp67_ASAP7_75t_SL g1451 ( 
.A(n_1102),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1294),
.A2(n_618),
.B1(n_625),
.B2(n_601),
.Y(n_1452)
);

AND2x6_ASAP7_75t_L g1453 ( 
.A(n_1080),
.B(n_533),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1250),
.Y(n_1454)
);

INVx5_ASAP7_75t_L g1455 ( 
.A(n_1146),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1258),
.Y(n_1456)
);

INVx4_ASAP7_75t_L g1457 ( 
.A(n_1084),
.Y(n_1457)
);

AND3x2_ASAP7_75t_L g1458 ( 
.A(n_1093),
.B(n_736),
.C(n_644),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1152),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1258),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1296),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1274),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1296),
.A2(n_630),
.B1(n_657),
.B2(n_628),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1084),
.Y(n_1464)
);

BUFx4f_ASAP7_75t_L g1465 ( 
.A(n_1095),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1199),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1075),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1274),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1199),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1277),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_1196),
.B(n_658),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1277),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1286),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1286),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1287),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1232),
.A2(n_795),
.B1(n_534),
.B2(n_576),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1264),
.A2(n_690),
.B1(n_693),
.B2(n_660),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1087),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1287),
.Y(n_1479)
);

INVxp33_ASAP7_75t_L g1480 ( 
.A(n_1135),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1081),
.Y(n_1481)
);

INVx8_ASAP7_75t_L g1482 ( 
.A(n_1118),
.Y(n_1482)
);

NAND3xp33_ASAP7_75t_L g1483 ( 
.A(n_1217),
.B(n_546),
.C(n_538),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1217),
.B(n_516),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1092),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1181),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1104),
.B(n_881),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1181),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1170),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1196),
.B(n_696),
.Y(n_1490)
);

INVx5_ASAP7_75t_L g1491 ( 
.A(n_1199),
.Y(n_1491)
);

OR2x6_ASAP7_75t_L g1492 ( 
.A(n_1273),
.B(n_795),
.Y(n_1492)
);

INVx5_ASAP7_75t_L g1493 ( 
.A(n_1199),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1120),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1206),
.B(n_700),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1112),
.B(n_882),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1206),
.B(n_706),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1145),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1221),
.Y(n_1499)
);

AND2x6_ASAP7_75t_L g1500 ( 
.A(n_1116),
.B(n_1125),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1121),
.Y(n_1501)
);

AO21x2_ASAP7_75t_L g1502 ( 
.A1(n_1261),
.A2(n_891),
.B(n_883),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1083),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1128),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1170),
.B(n_516),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1220),
.B(n_548),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1131),
.B(n_1058),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1171),
.B(n_549),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1171),
.B(n_731),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1133),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1143),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1221),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1150),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1156),
.Y(n_1514)
);

INVx5_ASAP7_75t_L g1515 ( 
.A(n_1199),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1172),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1172),
.B(n_560),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1182),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1158),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1161),
.A2(n_1056),
.B1(n_1053),
.B2(n_1039),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1182),
.B(n_737),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1164),
.B(n_892),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1167),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1174),
.Y(n_1524)
);

NAND2xp33_ASAP7_75t_L g1525 ( 
.A(n_1082),
.B(n_955),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1175),
.B(n_1042),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_SL g1527 ( 
.A1(n_1232),
.A2(n_562),
.B1(n_576),
.B2(n_534),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1082),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1176),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1183),
.B(n_563),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1186),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1183),
.B(n_744),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1190),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1191),
.B(n_1042),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1148),
.B(n_551),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1193),
.B(n_745),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1200),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1205),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1211),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1215),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1082),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1219),
.Y(n_1542)
);

NOR2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1118),
.B(n_551),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1226),
.B(n_564),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1229),
.B(n_1058),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1087),
.Y(n_1546)
);

INVx4_ASAP7_75t_L g1547 ( 
.A(n_1400),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1309),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1309),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1324),
.B(n_1231),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1312),
.B(n_1148),
.Y(n_1551)
);

INVxp33_ASAP7_75t_L g1552 ( 
.A(n_1368),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1324),
.A2(n_1239),
.B1(n_1246),
.B2(n_1240),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1302),
.B(n_1251),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1478),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1311),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1325),
.A2(n_1256),
.B1(n_1260),
.B2(n_1159),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1467),
.B(n_1262),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1308),
.B(n_1233),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1311),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1342),
.Y(n_1561)
);

AOI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1382),
.A2(n_1233),
.B1(n_1269),
.B2(n_1263),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1353),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1300),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1300),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1304),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1382),
.B(n_1124),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1304),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1342),
.Y(n_1569)
);

INVx2_ASAP7_75t_SL g1570 ( 
.A(n_1328),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1397),
.B(n_1124),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1350),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1481),
.Y(n_1573)
);

NAND2x1p5_ASAP7_75t_L g1574 ( 
.A(n_1312),
.B(n_1094),
.Y(n_1574)
);

OAI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1310),
.A2(n_1254),
.B1(n_1209),
.B2(n_1185),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1359),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1481),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1485),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1467),
.B(n_1275),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1312),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1312),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1353),
.Y(n_1582)
);

NAND2xp33_ASAP7_75t_L g1583 ( 
.A(n_1312),
.B(n_1134),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1400),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1350),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1397),
.B(n_1134),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1357),
.B(n_1254),
.Y(n_1587)
);

AO22x2_ASAP7_75t_L g1588 ( 
.A1(n_1351),
.A2(n_579),
.B1(n_586),
.B2(n_562),
.Y(n_1588)
);

NAND3x1_ASAP7_75t_L g1589 ( 
.A(n_1329),
.B(n_1180),
.C(n_1160),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1503),
.B(n_1276),
.Y(n_1590)
);

AND2x6_ASAP7_75t_L g1591 ( 
.A(n_1305),
.B(n_1278),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1328),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1421),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1401),
.B(n_1136),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1359),
.Y(n_1595)
);

AND2x6_ASAP7_75t_L g1596 ( 
.A(n_1305),
.B(n_1288),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1346),
.B(n_1209),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1361),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1478),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1361),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1318),
.A2(n_1245),
.B1(n_586),
.B2(n_589),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1485),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1301),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1480),
.A2(n_1224),
.B1(n_1266),
.B2(n_1265),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1301),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1362),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1318),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1362),
.Y(n_1608)
);

INVx4_ASAP7_75t_L g1609 ( 
.A(n_1400),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1301),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_SL g1611 ( 
.A(n_1421),
.B(n_1088),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1320),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1318),
.B(n_1153),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1365),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1318),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1320),
.Y(n_1616)
);

BUFx4f_ASAP7_75t_L g1617 ( 
.A(n_1482),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1357),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1407),
.A2(n_1153),
.B1(n_1140),
.B2(n_1144),
.Y(n_1619)
);

OR2x6_ASAP7_75t_L g1620 ( 
.A(n_1482),
.B(n_1091),
.Y(n_1620)
);

NAND3x1_ASAP7_75t_L g1621 ( 
.A(n_1319),
.B(n_1192),
.C(n_1184),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1459),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1318),
.B(n_1153),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1387),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1336),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1365),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1336),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1348),
.B(n_1136),
.Y(n_1628)
);

INVx4_ASAP7_75t_L g1629 ( 
.A(n_1400),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1404),
.B(n_1140),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1369),
.Y(n_1631)
);

AND2x6_ASAP7_75t_L g1632 ( 
.A(n_1306),
.B(n_1292),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_L g1633 ( 
.A(n_1387),
.Y(n_1633)
);

NAND3xp33_ASAP7_75t_L g1634 ( 
.A(n_1508),
.B(n_1266),
.C(n_1265),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1348),
.B(n_1144),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1401),
.A2(n_1189),
.B1(n_1173),
.B2(n_1165),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1387),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1337),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1461),
.B(n_1114),
.Y(n_1639)
);

INVx6_ASAP7_75t_L g1640 ( 
.A(n_1482),
.Y(n_1640)
);

INVx2_ASAP7_75t_SL g1641 ( 
.A(n_1374),
.Y(n_1641)
);

AND2x6_ASAP7_75t_L g1642 ( 
.A(n_1306),
.B(n_1145),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1346),
.B(n_1088),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1422),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1337),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1351),
.B(n_1100),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1459),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1366),
.B(n_1100),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1369),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_1341),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1546),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1381),
.Y(n_1652)
);

BUFx2_ASAP7_75t_L g1653 ( 
.A(n_1303),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1503),
.B(n_1094),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1381),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1338),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1338),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1333),
.Y(n_1658)
);

BUFx4_ASAP7_75t_L g1659 ( 
.A(n_1315),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1374),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1339),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1383),
.Y(n_1662)
);

INVx4_ASAP7_75t_L g1663 ( 
.A(n_1404),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1494),
.B(n_1094),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1433),
.B(n_1103),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1339),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1383),
.Y(n_1667)
);

NAND2x1p5_ASAP7_75t_L g1668 ( 
.A(n_1404),
.B(n_1109),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1461),
.B(n_1114),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1389),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1518),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1344),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1344),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1366),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1389),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1422),
.B(n_1103),
.Y(n_1676)
);

NAND2x1p5_ASAP7_75t_L g1677 ( 
.A(n_1465),
.B(n_1109),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1505),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1494),
.B(n_1109),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1498),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1390),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1387),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1519),
.B(n_1105),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1347),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1501),
.B(n_1423),
.Y(n_1685)
);

INVx8_ASAP7_75t_L g1686 ( 
.A(n_1482),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1498),
.Y(n_1687)
);

AND2x6_ASAP7_75t_L g1688 ( 
.A(n_1307),
.B(n_1145),
.Y(n_1688)
);

BUFx10_ASAP7_75t_L g1689 ( 
.A(n_1506),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1347),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1390),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1501),
.B(n_1451),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1379),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1355),
.B(n_1105),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1387),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1363),
.B(n_1108),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1498),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1393),
.Y(n_1698)
);

NAND2x1p5_ASAP7_75t_L g1699 ( 
.A(n_1465),
.B(n_1113),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1379),
.Y(n_1700)
);

AO22x2_ASAP7_75t_L g1701 ( 
.A1(n_1317),
.A2(n_589),
.B1(n_592),
.B2(n_579),
.Y(n_1701)
);

INVx8_ASAP7_75t_L g1702 ( 
.A(n_1500),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1465),
.B(n_1202),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1519),
.B(n_1108),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1402),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1316),
.B(n_1327),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1402),
.Y(n_1707)
);

INVxp67_ASAP7_75t_L g1708 ( 
.A(n_1375),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1405),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1434),
.Y(n_1710)
);

NAND2x1p5_ASAP7_75t_L g1711 ( 
.A(n_1313),
.B(n_1113),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1546),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1321),
.B(n_1111),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1523),
.B(n_1111),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1405),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1504),
.B(n_1113),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1484),
.B(n_1227),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1412),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1450),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1331),
.A2(n_1283),
.B1(n_1204),
.B2(n_1201),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1450),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1412),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1484),
.B(n_1227),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1431),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1376),
.B(n_550),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1393),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1415),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1415),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1392),
.B(n_550),
.Y(n_1729)
);

AND2x6_ASAP7_75t_L g1730 ( 
.A(n_1307),
.B(n_1201),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1417),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1505),
.B(n_1535),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1504),
.B(n_1510),
.Y(n_1733)
);

INVx8_ASAP7_75t_L g1734 ( 
.A(n_1500),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1516),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_1431),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1394),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1367),
.B(n_584),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1510),
.B(n_1227),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1523),
.B(n_592),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1417),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1403),
.B(n_584),
.Y(n_1742)
);

BUFx6f_ASAP7_75t_L g1743 ( 
.A(n_1431),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1380),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1431),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1323),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1323),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1394),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1419),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1419),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1431),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1524),
.B(n_600),
.Y(n_1752)
);

AO22x2_ASAP7_75t_L g1753 ( 
.A1(n_1483),
.A2(n_600),
.B1(n_612),
.B2(n_605),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1380),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1535),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1426),
.Y(n_1756)
);

AND2x6_ASAP7_75t_L g1757 ( 
.A(n_1322),
.B(n_1201),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1395),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1426),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1517),
.B(n_584),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1511),
.B(n_1255),
.Y(n_1761)
);

AO21x2_ASAP7_75t_L g1762 ( 
.A1(n_1525),
.A2(n_894),
.B(n_893),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1427),
.Y(n_1763)
);

O2A1O1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1527),
.A2(n_898),
.B(n_903),
.C(n_895),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1466),
.Y(n_1765)
);

INVx2_ASAP7_75t_SL g1766 ( 
.A(n_1516),
.Y(n_1766)
);

NOR3xp33_ASAP7_75t_L g1767 ( 
.A(n_1343),
.B(n_1163),
.C(n_1154),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1524),
.B(n_605),
.Y(n_1768)
);

INVx4_ASAP7_75t_L g1769 ( 
.A(n_1466),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1466),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1531),
.B(n_612),
.Y(n_1771)
);

AOI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1528),
.A2(n_1248),
.B1(n_1255),
.B2(n_1204),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1410),
.Y(n_1773)
);

BUFx6f_ASAP7_75t_L g1774 ( 
.A(n_1466),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1345),
.B(n_1204),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1427),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1372),
.B(n_1248),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1429),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1511),
.B(n_1248),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1531),
.B(n_619),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1429),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1513),
.B(n_1255),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1435),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1513),
.B(n_1271),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1530),
.B(n_584),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1410),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1428),
.Y(n_1787)
);

NAND2xp33_ASAP7_75t_L g1788 ( 
.A(n_1528),
.B(n_1202),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1435),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1489),
.B(n_1184),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1514),
.B(n_1271),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1364),
.B(n_1271),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1436),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1439),
.Y(n_1794)
);

INVxp67_ASAP7_75t_L g1795 ( 
.A(n_1438),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1552),
.B(n_1414),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1555),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1559),
.A2(n_1492),
.B1(n_1323),
.B2(n_1533),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1708),
.B(n_1418),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1549),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1549),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1559),
.A2(n_1492),
.B1(n_1323),
.B2(n_1533),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1548),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1556),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1708),
.A2(n_1409),
.B1(n_1441),
.B2(n_1424),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1585),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_SL g1807 ( 
.A1(n_1597),
.A2(n_1192),
.B1(n_1163),
.B2(n_1166),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1795),
.B(n_1438),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1758),
.B(n_1418),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1552),
.B(n_1509),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1758),
.B(n_1538),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1561),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1685),
.B(n_1542),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1560),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1692),
.B(n_1542),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1795),
.B(n_1514),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1597),
.B(n_1521),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1563),
.B(n_1529),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1563),
.B(n_1529),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1644),
.B(n_1538),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1755),
.B(n_1532),
.Y(n_1821)
);

INVx3_ASAP7_75t_L g1822 ( 
.A(n_1580),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1585),
.Y(n_1823)
);

NOR2x1p5_ASAP7_75t_L g1824 ( 
.A(n_1555),
.B(n_1443),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1561),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1582),
.B(n_1537),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1644),
.B(n_1539),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1755),
.B(n_1471),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1580),
.B(n_1539),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1706),
.A2(n_1349),
.B(n_1373),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1663),
.B(n_1540),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1580),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1580),
.B(n_1540),
.Y(n_1833)
);

INVx2_ASAP7_75t_SL g1834 ( 
.A(n_1581),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1581),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1569),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1581),
.B(n_1607),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1569),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_SL g1839 ( 
.A(n_1593),
.B(n_1434),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1582),
.B(n_1537),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1710),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1581),
.B(n_1420),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1607),
.B(n_1544),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1618),
.B(n_1487),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1607),
.B(n_1443),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1618),
.B(n_1487),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1607),
.B(n_1496),
.Y(n_1847)
);

AND2x4_ASAP7_75t_SL g1848 ( 
.A(n_1615),
.B(n_1441),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1733),
.B(n_1496),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1587),
.B(n_1441),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1576),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1564),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1565),
.Y(n_1853)
);

OAI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1641),
.A2(n_1441),
.B1(n_1356),
.B2(n_1492),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1554),
.B(n_1522),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1576),
.Y(n_1856)
);

INVxp67_ASAP7_75t_SL g1857 ( 
.A(n_1615),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1599),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1615),
.B(n_1522),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1601),
.B(n_1492),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1595),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1601),
.B(n_1356),
.Y(n_1862)
);

AND2x6_ASAP7_75t_SL g1863 ( 
.A(n_1696),
.B(n_1356),
.Y(n_1863)
);

AOI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1570),
.A2(n_1378),
.B1(n_1536),
.B2(n_1477),
.Y(n_1864)
);

BUFx6f_ASAP7_75t_L g1865 ( 
.A(n_1615),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1717),
.B(n_1723),
.Y(n_1866)
);

INVxp67_ASAP7_75t_L g1867 ( 
.A(n_1572),
.Y(n_1867)
);

BUFx12f_ASAP7_75t_L g1868 ( 
.A(n_1620),
.Y(n_1868)
);

OR2x6_ASAP7_75t_L g1869 ( 
.A(n_1686),
.B(n_1541),
.Y(n_1869)
);

NOR2x1p5_ASAP7_75t_L g1870 ( 
.A(n_1599),
.B(n_1315),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1595),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1650),
.A2(n_1541),
.B1(n_1354),
.B2(n_1388),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1598),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1592),
.A2(n_1391),
.B1(n_1500),
.B2(n_1495),
.Y(n_1874)
);

NAND2x1_ASAP7_75t_L g1875 ( 
.A(n_1769),
.B(n_1313),
.Y(n_1875)
);

INVx3_ASAP7_75t_L g1876 ( 
.A(n_1642),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1717),
.B(n_1436),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1566),
.B(n_1356),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1696),
.B(n_1490),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1660),
.B(n_1384),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1723),
.B(n_1437),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1598),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1568),
.B(n_1437),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1603),
.A2(n_1453),
.B1(n_1500),
.B2(n_1358),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_R g1885 ( 
.A(n_1617),
.B(n_1091),
.Y(n_1885)
);

BUFx2_ASAP7_75t_L g1886 ( 
.A(n_1735),
.Y(n_1886)
);

NOR2x1p5_ASAP7_75t_L g1887 ( 
.A(n_1651),
.B(n_1154),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1725),
.B(n_1456),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1729),
.B(n_1456),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1732),
.B(n_1497),
.Y(n_1890)
);

INVxp67_ASAP7_75t_L g1891 ( 
.A(n_1653),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1573),
.B(n_1470),
.Y(n_1892)
);

AND3x1_ASAP7_75t_L g1893 ( 
.A(n_1767),
.B(n_1636),
.C(n_1635),
.Y(n_1893)
);

NAND2x1p5_ASAP7_75t_L g1894 ( 
.A(n_1663),
.B(n_1341),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1605),
.A2(n_1453),
.B1(n_1500),
.B2(n_1335),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1577),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1578),
.B(n_1470),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1600),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1586),
.B(n_1370),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1551),
.A2(n_1500),
.B1(n_1452),
.B2(n_1463),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1586),
.B(n_1466),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1602),
.B(n_1472),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1610),
.A2(n_1777),
.B1(n_1746),
.B2(n_1747),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1694),
.B(n_1399),
.Y(n_1904)
);

INVx4_ASAP7_75t_L g1905 ( 
.A(n_1624),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1600),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1606),
.Y(n_1907)
);

INVx3_ASAP7_75t_L g1908 ( 
.A(n_1642),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1694),
.B(n_1411),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1651),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1547),
.B(n_1543),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1658),
.B(n_1476),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1606),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1594),
.B(n_1567),
.Y(n_1914)
);

NOR3xp33_ASAP7_75t_L g1915 ( 
.A(n_1713),
.B(n_1168),
.C(n_1166),
.Y(n_1915)
);

AOI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1777),
.A2(n_1453),
.B1(n_1314),
.B2(n_1502),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1547),
.B(n_1472),
.Y(n_1917)
);

NOR2x2_ASAP7_75t_L g1918 ( 
.A(n_1620),
.B(n_1322),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1674),
.B(n_1671),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1550),
.B(n_1473),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1594),
.B(n_1469),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1612),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1740),
.B(n_1502),
.Y(n_1923)
);

CKINVDCx11_ASAP7_75t_R g1924 ( 
.A(n_1620),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1567),
.B(n_1469),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1742),
.B(n_1473),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1746),
.A2(n_1453),
.B1(n_1314),
.B2(n_1502),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1608),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1608),
.Y(n_1929)
);

INVxp67_ASAP7_75t_SL g1930 ( 
.A(n_1624),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1747),
.A2(n_1453),
.B1(n_1475),
.B2(n_1474),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1614),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1674),
.B(n_1507),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1614),
.Y(n_1934)
);

INVxp67_ASAP7_75t_L g1935 ( 
.A(n_1622),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1571),
.B(n_1469),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1760),
.B(n_1474),
.Y(n_1937)
);

INVx2_ASAP7_75t_SL g1938 ( 
.A(n_1766),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1785),
.B(n_1475),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1740),
.A2(n_1453),
.B1(n_1479),
.B2(n_1460),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1775),
.B(n_1479),
.Y(n_1941)
);

NAND2x1p5_ASAP7_75t_L g1942 ( 
.A(n_1624),
.B(n_1637),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1626),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1626),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1571),
.B(n_1469),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1647),
.B(n_1326),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1631),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1631),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1665),
.B(n_1526),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1775),
.B(n_1428),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1558),
.B(n_1440),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1579),
.B(n_1440),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1628),
.B(n_1683),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1649),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1590),
.B(n_1738),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1752),
.B(n_1446),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1551),
.A2(n_1525),
.B1(n_1545),
.B2(n_1534),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1584),
.B(n_1446),
.Y(n_1958)
);

AOI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1613),
.A2(n_1488),
.B(n_1486),
.Y(n_1959)
);

INVx2_ASAP7_75t_SL g1960 ( 
.A(n_1678),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1649),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1652),
.Y(n_1962)
);

INVx3_ASAP7_75t_L g1963 ( 
.A(n_1642),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1752),
.B(n_1768),
.Y(n_1964)
);

A2O1A1Ixp33_ASAP7_75t_SL g1965 ( 
.A1(n_1792),
.A2(n_1371),
.B(n_1386),
.C(n_1341),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1768),
.B(n_1447),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1652),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1771),
.B(n_1447),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1665),
.B(n_1210),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1771),
.B(n_1454),
.Y(n_1970)
);

O2A1O1Ixp33_ASAP7_75t_L g1971 ( 
.A1(n_1764),
.A2(n_1462),
.B(n_1454),
.C(n_633),
.Y(n_1971)
);

INVx2_ASAP7_75t_SL g1972 ( 
.A(n_1574),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1780),
.A2(n_1753),
.B1(n_1619),
.B2(n_1584),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1683),
.B(n_1469),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1650),
.A2(n_1386),
.B1(n_1371),
.B2(n_1499),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1704),
.B(n_1313),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1642),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1780),
.B(n_1462),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1753),
.B(n_1326),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1704),
.B(n_1340),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1655),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1655),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1553),
.B(n_1439),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1792),
.B(n_1439),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1662),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1753),
.A2(n_1468),
.B1(n_1460),
.B2(n_1413),
.Y(n_1986)
);

BUFx3_ASAP7_75t_L g1987 ( 
.A(n_1712),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1714),
.B(n_1340),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1557),
.B(n_1460),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_L g1990 ( 
.A(n_1689),
.B(n_1210),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1616),
.B(n_1468),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1662),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1625),
.B(n_1468),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1712),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1627),
.B(n_1408),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1667),
.B(n_1670),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1714),
.B(n_1340),
.Y(n_1997)
);

BUFx3_ASAP7_75t_L g1998 ( 
.A(n_1719),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1638),
.B(n_1408),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1645),
.B(n_1408),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1656),
.B(n_1413),
.Y(n_2001)
);

NAND3xp33_ASAP7_75t_SL g2002 ( 
.A(n_1767),
.B(n_1168),
.C(n_1214),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1667),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1609),
.B(n_1330),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1670),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1675),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1657),
.B(n_1661),
.Y(n_2007)
);

NAND2xp33_ASAP7_75t_L g2008 ( 
.A(n_1702),
.B(n_1330),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1646),
.B(n_1648),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1675),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1666),
.B(n_1413),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1796),
.B(n_1689),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1855),
.B(n_1849),
.Y(n_2013)
);

BUFx2_ASAP7_75t_L g2014 ( 
.A(n_1886),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1813),
.B(n_1672),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1804),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1817),
.B(n_1643),
.Y(n_2017)
);

A2O1A1Ixp33_ASAP7_75t_L g2018 ( 
.A1(n_1904),
.A2(n_1713),
.B(n_1562),
.C(n_1617),
.Y(n_2018)
);

INVxp67_ASAP7_75t_SL g2019 ( 
.A(n_2004),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1815),
.B(n_1673),
.Y(n_2020)
);

INVx3_ASAP7_75t_L g2021 ( 
.A(n_2004),
.Y(n_2021)
);

BUFx3_ASAP7_75t_L g2022 ( 
.A(n_1998),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1808),
.B(n_1684),
.Y(n_2023)
);

OAI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_1909),
.A2(n_1611),
.B1(n_1634),
.B2(n_1790),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1865),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1804),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1801),
.Y(n_2027)
);

AND2x4_ASAP7_75t_L g2028 ( 
.A(n_1911),
.B(n_1719),
.Y(n_2028)
);

AND2x6_ASAP7_75t_SL g2029 ( 
.A(n_1990),
.B(n_1676),
.Y(n_2029)
);

NAND2x1p5_ASAP7_75t_L g2030 ( 
.A(n_1905),
.B(n_1609),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1801),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1862),
.B(n_1850),
.Y(n_2032)
);

NOR3xp33_ASAP7_75t_SL g2033 ( 
.A(n_2002),
.B(n_1214),
.C(n_1630),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_L g2034 ( 
.A(n_1879),
.B(n_1575),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_R g2035 ( 
.A(n_1841),
.B(n_1686),
.Y(n_2035)
);

BUFx4f_ASAP7_75t_L g2036 ( 
.A(n_1868),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_R g2037 ( 
.A(n_1841),
.B(n_1686),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1896),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1808),
.B(n_1690),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1812),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1803),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1949),
.B(n_1693),
.Y(n_2042)
);

BUFx6f_ASAP7_75t_L g2043 ( 
.A(n_1865),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1814),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_R g2045 ( 
.A(n_1839),
.B(n_1583),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1852),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1853),
.Y(n_2047)
);

BUFx2_ASAP7_75t_L g2048 ( 
.A(n_1886),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_1998),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1862),
.B(n_1676),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1955),
.B(n_1700),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1866),
.B(n_1705),
.Y(n_2052)
);

NOR2x1p5_ASAP7_75t_L g2053 ( 
.A(n_1868),
.B(n_1744),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1800),
.B(n_1707),
.Y(n_2054)
);

BUFx3_ASAP7_75t_L g2055 ( 
.A(n_1797),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_2004),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1800),
.B(n_1709),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_SL g2058 ( 
.A(n_1969),
.B(n_1091),
.Y(n_2058)
);

INVx2_ASAP7_75t_SL g2059 ( 
.A(n_1797),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1812),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1838),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1933),
.B(n_1715),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1996),
.B(n_1718),
.Y(n_2063)
);

NOR3xp33_ASAP7_75t_SL g2064 ( 
.A(n_1854),
.B(n_1630),
.C(n_566),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1922),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_R g2066 ( 
.A(n_1858),
.B(n_1744),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1996),
.B(n_1722),
.Y(n_2067)
);

OR2x6_ASAP7_75t_L g2068 ( 
.A(n_1870),
.B(n_1640),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1850),
.B(n_1721),
.Y(n_2069)
);

NAND2xp33_ASAP7_75t_SL g2070 ( 
.A(n_1885),
.B(n_1824),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1838),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1919),
.B(n_1639),
.Y(n_2072)
);

BUFx3_ASAP7_75t_L g2073 ( 
.A(n_1858),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_1924),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_1891),
.B(n_1754),
.Y(n_2075)
);

AND2x4_ASAP7_75t_L g2076 ( 
.A(n_1911),
.B(n_1721),
.Y(n_2076)
);

NAND2xp33_ASAP7_75t_SL g2077 ( 
.A(n_1887),
.B(n_1639),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_1806),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1851),
.Y(n_2079)
);

BUFx2_ASAP7_75t_L g2080 ( 
.A(n_1823),
.Y(n_2080)
);

BUFx6f_ASAP7_75t_L g2081 ( 
.A(n_1865),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1810),
.B(n_1669),
.Y(n_2082)
);

NOR3xp33_ASAP7_75t_SL g2083 ( 
.A(n_1799),
.B(n_567),
.C(n_565),
.Y(n_2083)
);

NOR2xp33_ASAP7_75t_L g2084 ( 
.A(n_1867),
.B(n_1754),
.Y(n_2084)
);

BUFx8_ASAP7_75t_L g2085 ( 
.A(n_1910),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1865),
.Y(n_2086)
);

OR2x6_ASAP7_75t_L g2087 ( 
.A(n_1914),
.B(n_1640),
.Y(n_2087)
);

NOR3xp33_ASAP7_75t_SL g2088 ( 
.A(n_1809),
.B(n_573),
.C(n_571),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1946),
.Y(n_2089)
);

BUFx2_ASAP7_75t_L g2090 ( 
.A(n_1910),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1946),
.Y(n_2091)
);

CKINVDCx8_ASAP7_75t_R g2092 ( 
.A(n_1863),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1920),
.B(n_1727),
.Y(n_2093)
);

INVx3_ASAP7_75t_L g2094 ( 
.A(n_1831),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1851),
.Y(n_2095)
);

AND2x4_ASAP7_75t_L g2096 ( 
.A(n_1911),
.B(n_1629),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1860),
.B(n_1669),
.Y(n_2097)
);

OR2x6_ASAP7_75t_L g2098 ( 
.A(n_1964),
.B(n_1640),
.Y(n_2098)
);

NOR3xp33_ASAP7_75t_SL g2099 ( 
.A(n_1890),
.B(n_578),
.C(n_575),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_1860),
.A2(n_1701),
.B1(n_1629),
.B2(n_553),
.Y(n_2100)
);

BUFx6f_ASAP7_75t_L g2101 ( 
.A(n_1865),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1825),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_1935),
.B(n_1604),
.Y(n_2103)
);

INVx1_ASAP7_75t_SL g2104 ( 
.A(n_1938),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_1987),
.B(n_1728),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1825),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1830),
.B(n_1731),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_1912),
.B(n_1654),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_R g2109 ( 
.A(n_1987),
.B(n_1702),
.Y(n_2109)
);

NOR3xp33_ASAP7_75t_SL g2110 ( 
.A(n_1953),
.B(n_581),
.C(n_580),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_1878),
.B(n_1994),
.Y(n_2111)
);

BUFx6f_ASAP7_75t_L g2112 ( 
.A(n_1938),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_1878),
.B(n_1741),
.Y(n_2113)
);

NOR2x1_ASAP7_75t_L g2114 ( 
.A(n_1869),
.B(n_1769),
.Y(n_2114)
);

BUFx3_ASAP7_75t_L g2115 ( 
.A(n_1960),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1836),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1836),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_L g2118 ( 
.A(n_1828),
.B(n_1750),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1856),
.Y(n_2119)
);

BUFx2_ASAP7_75t_L g2120 ( 
.A(n_1960),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1888),
.B(n_1749),
.Y(n_2121)
);

CKINVDCx14_ASAP7_75t_R g2122 ( 
.A(n_1924),
.Y(n_2122)
);

BUFx2_ASAP7_75t_L g2123 ( 
.A(n_1893),
.Y(n_2123)
);

AND2x4_ASAP7_75t_L g2124 ( 
.A(n_1974),
.B(n_1756),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1861),
.Y(n_2125)
);

CKINVDCx20_ASAP7_75t_R g2126 ( 
.A(n_2009),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1889),
.B(n_1759),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1861),
.Y(n_2128)
);

BUFx12f_ASAP7_75t_L g2129 ( 
.A(n_1834),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1856),
.Y(n_2130)
);

CKINVDCx5p33_ASAP7_75t_R g2131 ( 
.A(n_1807),
.Y(n_2131)
);

INVxp67_ASAP7_75t_SL g2132 ( 
.A(n_2008),
.Y(n_2132)
);

AND2x6_ASAP7_75t_L g2133 ( 
.A(n_1876),
.B(n_1332),
.Y(n_2133)
);

AOI22xp33_ASAP7_75t_L g2134 ( 
.A1(n_1903),
.A2(n_1899),
.B1(n_1821),
.B2(n_1923),
.Y(n_2134)
);

NAND2x1p5_ASAP7_75t_L g2135 ( 
.A(n_1905),
.B(n_1624),
.Y(n_2135)
);

HB1xp67_ASAP7_75t_L g2136 ( 
.A(n_1942),
.Y(n_2136)
);

BUFx2_ASAP7_75t_L g2137 ( 
.A(n_1822),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1882),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_1923),
.A2(n_1701),
.B1(n_1776),
.B2(n_1763),
.Y(n_2139)
);

NAND2xp33_ASAP7_75t_R g2140 ( 
.A(n_1831),
.B(n_1680),
.Y(n_2140)
);

INVx5_ASAP7_75t_L g2141 ( 
.A(n_1869),
.Y(n_2141)
);

BUFx6f_ASAP7_75t_L g2142 ( 
.A(n_1834),
.Y(n_2142)
);

AND2x4_ASAP7_75t_L g2143 ( 
.A(n_1831),
.B(n_1778),
.Y(n_2143)
);

AOI211xp5_ASAP7_75t_L g2144 ( 
.A1(n_1915),
.A2(n_1764),
.B(n_619),
.C(n_636),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1871),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1816),
.B(n_1781),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1882),
.Y(n_2147)
);

AND3x2_ASAP7_75t_SL g2148 ( 
.A(n_1918),
.B(n_1588),
.C(n_1701),
.Y(n_2148)
);

NOR2xp67_ASAP7_75t_L g2149 ( 
.A(n_1805),
.B(n_1845),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1818),
.B(n_1783),
.Y(n_2150)
);

INVxp33_ASAP7_75t_L g2151 ( 
.A(n_1844),
.Y(n_2151)
);

OR2x6_ASAP7_75t_L g2152 ( 
.A(n_1869),
.B(n_1702),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1898),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1898),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1819),
.B(n_1789),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1826),
.B(n_1793),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1906),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1840),
.B(n_1664),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1871),
.Y(n_2159)
);

BUFx8_ASAP7_75t_L g2160 ( 
.A(n_1979),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1846),
.B(n_1679),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1906),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_1811),
.B(n_1703),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1873),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1869),
.Y(n_2165)
);

BUFx8_ASAP7_75t_SL g2166 ( 
.A(n_1822),
.Y(n_2166)
);

AND2x4_ASAP7_75t_L g2167 ( 
.A(n_1848),
.B(n_1680),
.Y(n_2167)
);

INVx6_ASAP7_75t_L g2168 ( 
.A(n_1905),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1926),
.B(n_1681),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_SL g2170 ( 
.A(n_1937),
.B(n_1774),
.Y(n_2170)
);

CKINVDCx20_ASAP7_75t_R g2171 ( 
.A(n_1848),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_R g2172 ( 
.A(n_1822),
.B(n_1734),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1907),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_1832),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1939),
.B(n_1681),
.Y(n_2175)
);

OR2x6_ASAP7_75t_L g2176 ( 
.A(n_1976),
.B(n_1734),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1907),
.Y(n_2177)
);

NOR3xp33_ASAP7_75t_SL g2178 ( 
.A(n_1842),
.B(n_590),
.C(n_582),
.Y(n_2178)
);

BUFx2_ASAP7_75t_L g2179 ( 
.A(n_1832),
.Y(n_2179)
);

NOR3xp33_ASAP7_75t_SL g2180 ( 
.A(n_1901),
.B(n_593),
.C(n_591),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_R g2181 ( 
.A(n_1832),
.B(n_1734),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1913),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1913),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_R g2184 ( 
.A(n_1835),
.B(n_1687),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_L g2185 ( 
.A(n_1880),
.B(n_1703),
.Y(n_2185)
);

CKINVDCx5p33_ASAP7_75t_R g2186 ( 
.A(n_1864),
.Y(n_2186)
);

BUFx2_ASAP7_75t_L g2187 ( 
.A(n_1918),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_R g2188 ( 
.A(n_1835),
.B(n_1687),
.Y(n_2188)
);

BUFx10_ASAP7_75t_L g2189 ( 
.A(n_1917),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1873),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1934),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1979),
.B(n_1691),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1798),
.B(n_1633),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_1980),
.B(n_1697),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1802),
.B(n_1633),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1934),
.Y(n_2196)
);

BUFx6f_ASAP7_75t_L g2197 ( 
.A(n_1942),
.Y(n_2197)
);

AND2x4_ASAP7_75t_L g2198 ( 
.A(n_1988),
.B(n_1697),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1943),
.Y(n_2199)
);

BUFx3_ASAP7_75t_L g2200 ( 
.A(n_1942),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1928),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1928),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1877),
.B(n_1691),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1929),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1929),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_1820),
.B(n_1613),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1932),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1932),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1944),
.Y(n_2209)
);

INVx4_ASAP7_75t_L g2210 ( 
.A(n_1917),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1881),
.B(n_1698),
.Y(n_2211)
);

INVx3_ASAP7_75t_L g2212 ( 
.A(n_1958),
.Y(n_2212)
);

NOR3xp33_ASAP7_75t_SL g2213 ( 
.A(n_1921),
.B(n_598),
.C(n_597),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2007),
.B(n_1698),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1944),
.Y(n_2215)
);

NOR3xp33_ASAP7_75t_SL g2216 ( 
.A(n_1925),
.B(n_602),
.C(n_599),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1943),
.Y(n_2217)
);

BUFx10_ASAP7_75t_L g2218 ( 
.A(n_1917),
.Y(n_2218)
);

BUFx4f_ASAP7_75t_L g2219 ( 
.A(n_1972),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1947),
.Y(n_2220)
);

INVxp67_ASAP7_75t_L g2221 ( 
.A(n_1827),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1948),
.Y(n_2222)
);

AOI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_1997),
.A2(n_1589),
.B1(n_1621),
.B2(n_1623),
.Y(n_2223)
);

NAND3xp33_ASAP7_75t_SL g2224 ( 
.A(n_1874),
.B(n_1699),
.C(n_1677),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1941),
.B(n_1726),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1947),
.Y(n_2226)
);

AND2x4_ASAP7_75t_L g2227 ( 
.A(n_1936),
.B(n_1794),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1954),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1954),
.Y(n_2229)
);

OR2x6_ASAP7_75t_L g2230 ( 
.A(n_1945),
.B(n_1574),
.Y(n_2230)
);

OA22x2_ASAP7_75t_L g2231 ( 
.A1(n_1900),
.A2(n_1458),
.B1(n_604),
.B2(n_606),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1962),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1962),
.B(n_1726),
.Y(n_2233)
);

INVx3_ASAP7_75t_L g2234 ( 
.A(n_1958),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_SL g2235 ( 
.A(n_1973),
.B(n_1958),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_1948),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1981),
.B(n_1982),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1981),
.Y(n_2238)
);

HB1xp67_ASAP7_75t_L g2239 ( 
.A(n_1847),
.Y(n_2239)
);

AO21x2_ASAP7_75t_L g2240 ( 
.A1(n_1965),
.A2(n_1623),
.B(n_1762),
.Y(n_2240)
);

BUFx3_ASAP7_75t_L g2241 ( 
.A(n_1972),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1982),
.B(n_1737),
.Y(n_2242)
);

INVx3_ASAP7_75t_SL g2243 ( 
.A(n_1837),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2005),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_2005),
.Y(n_2245)
);

BUFx6f_ASAP7_75t_L g2246 ( 
.A(n_1876),
.Y(n_2246)
);

AND2x6_ASAP7_75t_L g2247 ( 
.A(n_2094),
.B(n_1876),
.Y(n_2247)
);

OAI21x1_ASAP7_75t_L g2248 ( 
.A1(n_2224),
.A2(n_1959),
.B(n_1975),
.Y(n_2248)
);

AO31x2_ASAP7_75t_L g2249 ( 
.A1(n_2107),
.A2(n_1872),
.A3(n_1950),
.B(n_1989),
.Y(n_2249)
);

BUFx2_ASAP7_75t_L g2250 ( 
.A(n_2014),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2013),
.B(n_1984),
.Y(n_2251)
);

OAI21xp5_ASAP7_75t_L g2252 ( 
.A1(n_2107),
.A2(n_1957),
.B(n_1916),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_2028),
.B(n_1857),
.Y(n_2253)
);

OAI21x1_ASAP7_75t_L g2254 ( 
.A1(n_2224),
.A2(n_1894),
.B(n_1908),
.Y(n_2254)
);

OAI21x1_ASAP7_75t_L g2255 ( 
.A1(n_2132),
.A2(n_1894),
.B(n_1908),
.Y(n_2255)
);

AOI21x1_ASAP7_75t_L g2256 ( 
.A1(n_2149),
.A2(n_1843),
.B(n_1833),
.Y(n_2256)
);

CKINVDCx20_ASAP7_75t_R g2257 ( 
.A(n_2126),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2016),
.Y(n_2258)
);

BUFx2_ASAP7_75t_L g2259 ( 
.A(n_2048),
.Y(n_2259)
);

AOI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_2132),
.A2(n_2008),
.B(n_1788),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2013),
.B(n_2010),
.Y(n_2261)
);

AND2x4_ASAP7_75t_L g2262 ( 
.A(n_2028),
.B(n_1859),
.Y(n_2262)
);

AOI21xp5_ASAP7_75t_L g2263 ( 
.A1(n_2019),
.A2(n_1788),
.B(n_1875),
.Y(n_2263)
);

INVx6_ASAP7_75t_L g2264 ( 
.A(n_2085),
.Y(n_2264)
);

A2O1A1Ixp33_ASAP7_75t_L g2265 ( 
.A1(n_2034),
.A2(n_1971),
.B(n_1983),
.C(n_1927),
.Y(n_2265)
);

NAND2x1p5_ASAP7_75t_L g2266 ( 
.A(n_2141),
.B(n_1908),
.Y(n_2266)
);

AO31x2_ASAP7_75t_L g2267 ( 
.A1(n_2206),
.A2(n_2010),
.A3(n_1951),
.B(n_1952),
.Y(n_2267)
);

AOI21x1_ASAP7_75t_L g2268 ( 
.A1(n_2193),
.A2(n_1829),
.B(n_1875),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_2186),
.B(n_1956),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_L g2270 ( 
.A(n_2017),
.B(n_2108),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_2066),
.Y(n_2271)
);

OAI21x1_ASAP7_75t_L g2272 ( 
.A1(n_2225),
.A2(n_1894),
.B(n_1963),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2032),
.B(n_1588),
.Y(n_2273)
);

OAI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2118),
.A2(n_1940),
.B1(n_1931),
.B2(n_1588),
.Y(n_2274)
);

AOI21xp33_ASAP7_75t_L g2275 ( 
.A1(n_2231),
.A2(n_1968),
.B(n_1966),
.Y(n_2275)
);

AOI21xp5_ASAP7_75t_L g2276 ( 
.A1(n_2019),
.A2(n_1895),
.B(n_1884),
.Y(n_2276)
);

OAI21x1_ASAP7_75t_L g2277 ( 
.A1(n_2225),
.A2(n_1977),
.B(n_1963),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2052),
.B(n_2003),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2026),
.Y(n_2279)
);

OAI21x1_ASAP7_75t_L g2280 ( 
.A1(n_2233),
.A2(n_1977),
.B(n_1963),
.Y(n_2280)
);

A2O1A1Ixp33_ASAP7_75t_L g2281 ( 
.A1(n_2018),
.A2(n_1978),
.B(n_1970),
.C(n_1892),
.Y(n_2281)
);

AOI21xp5_ASAP7_75t_L g2282 ( 
.A1(n_2042),
.A2(n_1377),
.B(n_1352),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2052),
.B(n_2003),
.Y(n_2283)
);

BUFx6f_ASAP7_75t_L g2284 ( 
.A(n_2022),
.Y(n_2284)
);

AO31x2_ASAP7_75t_L g2285 ( 
.A1(n_2185),
.A2(n_1961),
.A3(n_1985),
.B(n_1967),
.Y(n_2285)
);

OAI21x1_ASAP7_75t_L g2286 ( 
.A1(n_2233),
.A2(n_2242),
.B(n_2114),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2038),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2042),
.B(n_2015),
.Y(n_2288)
);

INVx6_ASAP7_75t_L g2289 ( 
.A(n_2085),
.Y(n_2289)
);

O2A1O1Ixp5_ASAP7_75t_L g2290 ( 
.A1(n_2195),
.A2(n_1977),
.B(n_1883),
.C(n_1902),
.Y(n_2290)
);

AOI21xp5_ASAP7_75t_L g2291 ( 
.A1(n_2015),
.A2(n_1377),
.B(n_1352),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2097),
.B(n_1961),
.Y(n_2292)
);

AO21x2_ASAP7_75t_L g2293 ( 
.A1(n_2240),
.A2(n_1762),
.B(n_1897),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2020),
.B(n_1967),
.Y(n_2294)
);

OR2x2_ASAP7_75t_L g2295 ( 
.A(n_2089),
.B(n_1985),
.Y(n_2295)
);

INVx3_ASAP7_75t_L g2296 ( 
.A(n_2168),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2041),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2069),
.B(n_1992),
.Y(n_2298)
);

AOI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2020),
.A2(n_1377),
.B(n_1352),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2158),
.B(n_1992),
.Y(n_2300)
);

OAI21x1_ASAP7_75t_L g2301 ( 
.A1(n_2242),
.A2(n_2211),
.B(n_2203),
.Y(n_2301)
);

OAI21xp5_ASAP7_75t_L g2302 ( 
.A1(n_2163),
.A2(n_1986),
.B(n_1716),
.Y(n_2302)
);

HB1xp67_ASAP7_75t_L g2303 ( 
.A(n_2080),
.Y(n_2303)
);

OAI21x1_ASAP7_75t_L g2304 ( 
.A1(n_2203),
.A2(n_1406),
.B(n_1668),
.Y(n_2304)
);

AOI21xp5_ASAP7_75t_L g2305 ( 
.A1(n_2093),
.A2(n_1396),
.B(n_1385),
.Y(n_2305)
);

NAND2x1p5_ASAP7_75t_L g2306 ( 
.A(n_2141),
.B(n_1633),
.Y(n_2306)
);

AOI21xp5_ASAP7_75t_L g2307 ( 
.A1(n_2093),
.A2(n_1396),
.B(n_1385),
.Y(n_2307)
);

A2O1A1Ixp33_ASAP7_75t_L g2308 ( 
.A1(n_2178),
.A2(n_1993),
.B(n_1995),
.C(n_1991),
.Y(n_2308)
);

OAI21x1_ASAP7_75t_L g2309 ( 
.A1(n_2211),
.A2(n_1406),
.B(n_1668),
.Y(n_2309)
);

OAI21x1_ASAP7_75t_L g2310 ( 
.A1(n_2192),
.A2(n_1386),
.B(n_1371),
.Y(n_2310)
);

AOI21xp5_ASAP7_75t_L g2311 ( 
.A1(n_2158),
.A2(n_1396),
.B(n_1385),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2161),
.B(n_2006),
.Y(n_2312)
);

AOI21xp5_ASAP7_75t_L g2313 ( 
.A1(n_2051),
.A2(n_1457),
.B(n_1432),
.Y(n_2313)
);

AOI21xp5_ASAP7_75t_L g2314 ( 
.A1(n_2051),
.A2(n_1457),
.B(n_1432),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2027),
.Y(n_2315)
);

AND3x4_ASAP7_75t_L g2316 ( 
.A(n_2033),
.B(n_1659),
.C(n_648),
.Y(n_2316)
);

NAND2x1_ASAP7_75t_L g2317 ( 
.A(n_2152),
.B(n_1682),
.Y(n_2317)
);

AOI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2062),
.A2(n_1457),
.B(n_1432),
.Y(n_2318)
);

A2O1A1Ixp33_ASAP7_75t_L g2319 ( 
.A1(n_2178),
.A2(n_2000),
.B(n_2001),
.C(n_1999),
.Y(n_2319)
);

AOI21xp5_ASAP7_75t_L g2320 ( 
.A1(n_2062),
.A2(n_1464),
.B(n_1398),
.Y(n_2320)
);

INVx3_ASAP7_75t_L g2321 ( 
.A(n_2168),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2161),
.B(n_2006),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2031),
.Y(n_2323)
);

AOI21x1_ASAP7_75t_SL g2324 ( 
.A1(n_2121),
.A2(n_2011),
.B(n_1791),
.Y(n_2324)
);

OAI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_2134),
.A2(n_2231),
.B(n_2192),
.Y(n_2325)
);

AOI21x1_ASAP7_75t_L g2326 ( 
.A1(n_2170),
.A2(n_1761),
.B(n_1739),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_2121),
.A2(n_1464),
.B(n_1398),
.Y(n_2327)
);

OAI21x1_ASAP7_75t_L g2328 ( 
.A1(n_2237),
.A2(n_1699),
.B(n_1677),
.Y(n_2328)
);

A2O1A1Ixp33_ASAP7_75t_L g2329 ( 
.A1(n_2064),
.A2(n_1930),
.B(n_1772),
.C(n_1782),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2040),
.Y(n_2330)
);

AOI21xp5_ASAP7_75t_L g2331 ( 
.A1(n_2127),
.A2(n_1464),
.B(n_1398),
.Y(n_2331)
);

AOI21xp33_ASAP7_75t_L g2332 ( 
.A1(n_2024),
.A2(n_1784),
.B(n_1779),
.Y(n_2332)
);

OAI21x1_ASAP7_75t_L g2333 ( 
.A1(n_2237),
.A2(n_1711),
.B(n_1737),
.Y(n_2333)
);

AND2x2_ASAP7_75t_SL g2334 ( 
.A(n_2058),
.B(n_633),
.Y(n_2334)
);

AO31x2_ASAP7_75t_L g2335 ( 
.A1(n_2102),
.A2(n_1488),
.A3(n_1499),
.B(n_1486),
.Y(n_2335)
);

BUFx3_ASAP7_75t_L g2336 ( 
.A(n_2055),
.Y(n_2336)
);

OAI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2169),
.A2(n_1720),
.B(n_1596),
.Y(n_2337)
);

OR2x2_ASAP7_75t_L g2338 ( 
.A(n_2091),
.B(n_1748),
.Y(n_2338)
);

OAI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_2169),
.A2(n_1596),
.B(n_1591),
.Y(n_2339)
);

OAI21xp5_ASAP7_75t_L g2340 ( 
.A1(n_2175),
.A2(n_1596),
.B(n_1591),
.Y(n_2340)
);

OA21x2_ASAP7_75t_L g2341 ( 
.A1(n_2235),
.A2(n_1512),
.B(n_1748),
.Y(n_2341)
);

OAI21x1_ASAP7_75t_L g2342 ( 
.A1(n_2054),
.A2(n_1711),
.B(n_1773),
.Y(n_2342)
);

BUFx2_ASAP7_75t_L g2343 ( 
.A(n_2111),
.Y(n_2343)
);

OAI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_2175),
.A2(n_1596),
.B(n_1591),
.Y(n_2344)
);

OAI21x1_ASAP7_75t_L g2345 ( 
.A1(n_2054),
.A2(n_1786),
.B(n_1773),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2060),
.Y(n_2346)
);

A2O1A1Ixp33_ASAP7_75t_L g2347 ( 
.A1(n_2064),
.A2(n_907),
.B(n_908),
.C(n_906),
.Y(n_2347)
);

OR2x2_ASAP7_75t_L g2348 ( 
.A(n_2078),
.B(n_1786),
.Y(n_2348)
);

A2O1A1Ixp33_ASAP7_75t_L g2349 ( 
.A1(n_2144),
.A2(n_912),
.B(n_917),
.C(n_911),
.Y(n_2349)
);

A2O1A1Ixp33_ASAP7_75t_L g2350 ( 
.A1(n_2099),
.A2(n_921),
.B(n_922),
.C(n_919),
.Y(n_2350)
);

AOI21xp5_ASAP7_75t_L g2351 ( 
.A1(n_2127),
.A2(n_1398),
.B(n_1360),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2146),
.B(n_1787),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2061),
.Y(n_2353)
);

AOI21xp5_ASAP7_75t_L g2354 ( 
.A1(n_2146),
.A2(n_1398),
.B(n_1360),
.Y(n_2354)
);

AOI21x1_ASAP7_75t_L g2355 ( 
.A1(n_2187),
.A2(n_1787),
.B(n_1512),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2123),
.B(n_1724),
.Y(n_2356)
);

AOI21xp33_ASAP7_75t_L g2357 ( 
.A1(n_2140),
.A2(n_1794),
.B(n_637),
.Y(n_2357)
);

NAND2x1p5_ASAP7_75t_L g2358 ( 
.A(n_2141),
.B(n_1633),
.Y(n_2358)
);

OAI21xp5_ASAP7_75t_L g2359 ( 
.A1(n_2023),
.A2(n_1596),
.B(n_1591),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_2073),
.Y(n_2360)
);

OR2x2_ASAP7_75t_L g2361 ( 
.A(n_2111),
.B(n_1332),
.Y(n_2361)
);

NAND3xp33_ASAP7_75t_L g2362 ( 
.A(n_2099),
.B(n_607),
.C(n_603),
.Y(n_2362)
);

OR2x2_ASAP7_75t_L g2363 ( 
.A(n_2050),
.B(n_1334),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2044),
.Y(n_2364)
);

OAI21xp5_ASAP7_75t_L g2365 ( 
.A1(n_2023),
.A2(n_2039),
.B(n_2214),
.Y(n_2365)
);

OAI21x1_ASAP7_75t_L g2366 ( 
.A1(n_2057),
.A2(n_1416),
.B(n_1334),
.Y(n_2366)
);

OAI21x1_ASAP7_75t_L g2367 ( 
.A1(n_2057),
.A2(n_1416),
.B(n_1442),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2151),
.B(n_704),
.Y(n_2368)
);

OAI21x1_ASAP7_75t_L g2369 ( 
.A1(n_2214),
.A2(n_1416),
.B(n_1444),
.Y(n_2369)
);

OAI21x1_ASAP7_75t_L g2370 ( 
.A1(n_2106),
.A2(n_2117),
.B(n_2116),
.Y(n_2370)
);

INVx3_ASAP7_75t_L g2371 ( 
.A(n_2168),
.Y(n_2371)
);

CKINVDCx8_ASAP7_75t_R g2372 ( 
.A(n_2029),
.Y(n_2372)
);

BUFx2_ASAP7_75t_SL g2373 ( 
.A(n_2171),
.Y(n_2373)
);

AOI221xp5_ASAP7_75t_SL g2374 ( 
.A1(n_2100),
.A2(n_639),
.B1(n_647),
.B2(n_637),
.C(n_636),
.Y(n_2374)
);

AOI21xp5_ASAP7_75t_L g2375 ( 
.A1(n_2150),
.A2(n_1455),
.B(n_1360),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2150),
.B(n_1591),
.Y(n_2376)
);

O2A1O1Ixp5_ASAP7_75t_L g2377 ( 
.A1(n_2012),
.A2(n_639),
.B(n_654),
.C(n_647),
.Y(n_2377)
);

OAI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_2155),
.A2(n_1682),
.B1(n_1695),
.B2(n_1637),
.Y(n_2378)
);

BUFx2_ASAP7_75t_L g2379 ( 
.A(n_2090),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2155),
.B(n_1632),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2046),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2082),
.A2(n_786),
.B1(n_776),
.B2(n_609),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_2076),
.B(n_1637),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_2072),
.B(n_1774),
.Y(n_2384)
);

OAI21x1_ASAP7_75t_L g2385 ( 
.A1(n_2125),
.A2(n_1445),
.B(n_1520),
.Y(n_2385)
);

HB1xp67_ASAP7_75t_L g2386 ( 
.A(n_2120),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2156),
.B(n_2063),
.Y(n_2387)
);

OR2x2_ASAP7_75t_L g2388 ( 
.A(n_2113),
.B(n_939),
.Y(n_2388)
);

AOI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2156),
.A2(n_1455),
.B(n_1360),
.Y(n_2389)
);

BUFx2_ASAP7_75t_L g2390 ( 
.A(n_2115),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2063),
.B(n_1632),
.Y(n_2391)
);

INVx4_ASAP7_75t_L g2392 ( 
.A(n_2112),
.Y(n_2392)
);

OR2x2_ASAP7_75t_L g2393 ( 
.A(n_2113),
.B(n_939),
.Y(n_2393)
);

AOI21xp5_ASAP7_75t_L g2394 ( 
.A1(n_2067),
.A2(n_1455),
.B(n_1360),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2076),
.B(n_2221),
.Y(n_2395)
);

OAI22x1_ASAP7_75t_L g2396 ( 
.A1(n_2223),
.A2(n_655),
.B1(n_661),
.B2(n_654),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2067),
.B(n_1632),
.Y(n_2397)
);

OAI21x1_ASAP7_75t_L g2398 ( 
.A1(n_2128),
.A2(n_1449),
.B(n_1448),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2071),
.Y(n_2399)
);

BUFx4f_ASAP7_75t_SL g2400 ( 
.A(n_2129),
.Y(n_2400)
);

CKINVDCx5p33_ASAP7_75t_R g2401 ( 
.A(n_2074),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2047),
.Y(n_2402)
);

OAI21x1_ASAP7_75t_L g2403 ( 
.A1(n_2138),
.A2(n_1430),
.B(n_1053),
.Y(n_2403)
);

AOI21xp5_ASAP7_75t_L g2404 ( 
.A1(n_2240),
.A2(n_1491),
.B(n_1455),
.Y(n_2404)
);

OAI21x1_ASAP7_75t_L g2405 ( 
.A1(n_2147),
.A2(n_1039),
.B(n_1425),
.Y(n_2405)
);

CKINVDCx5p33_ASAP7_75t_R g2406 ( 
.A(n_2122),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2079),
.Y(n_2407)
);

OAI21x1_ASAP7_75t_L g2408 ( 
.A1(n_2153),
.A2(n_970),
.B(n_942),
.Y(n_2408)
);

NOR2x1_ASAP7_75t_L g2409 ( 
.A(n_2068),
.B(n_1745),
.Y(n_2409)
);

BUFx8_ASAP7_75t_L g2410 ( 
.A(n_2112),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2065),
.Y(n_2411)
);

NAND2x1_ASAP7_75t_L g2412 ( 
.A(n_2152),
.B(n_1745),
.Y(n_2412)
);

NAND2x1_ASAP7_75t_L g2413 ( 
.A(n_2152),
.B(n_1745),
.Y(n_2413)
);

OAI21x1_ASAP7_75t_L g2414 ( 
.A1(n_2154),
.A2(n_970),
.B(n_942),
.Y(n_2414)
);

OAI21x1_ASAP7_75t_L g2415 ( 
.A1(n_2157),
.A2(n_970),
.B(n_943),
.Y(n_2415)
);

INVx6_ASAP7_75t_L g2416 ( 
.A(n_2189),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_SL g2417 ( 
.A(n_2045),
.B(n_1637),
.Y(n_2417)
);

AOI22xp33_ASAP7_75t_SL g2418 ( 
.A1(n_2131),
.A2(n_648),
.B1(n_561),
.B2(n_704),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2162),
.Y(n_2419)
);

OAI21xp5_ASAP7_75t_L g2420 ( 
.A1(n_2039),
.A2(n_1632),
.B(n_1642),
.Y(n_2420)
);

BUFx8_ASAP7_75t_L g2421 ( 
.A(n_2112),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2139),
.B(n_1632),
.Y(n_2422)
);

OAI21x1_ASAP7_75t_L g2423 ( 
.A1(n_2173),
.A2(n_943),
.B(n_940),
.Y(n_2423)
);

AOI21xp5_ASAP7_75t_L g2424 ( 
.A1(n_2176),
.A2(n_1491),
.B(n_1455),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2177),
.Y(n_2425)
);

AND2x4_ASAP7_75t_L g2426 ( 
.A(n_2096),
.B(n_1682),
.Y(n_2426)
);

OAI21xp5_ASAP7_75t_L g2427 ( 
.A1(n_2221),
.A2(n_1730),
.B(n_1688),
.Y(n_2427)
);

BUFx2_ASAP7_75t_L g2428 ( 
.A(n_2174),
.Y(n_2428)
);

AND2x6_ASAP7_75t_L g2429 ( 
.A(n_2094),
.B(n_1682),
.Y(n_2429)
);

OAI21xp5_ASAP7_75t_L g2430 ( 
.A1(n_2124),
.A2(n_1730),
.B(n_1688),
.Y(n_2430)
);

AOI21xp5_ASAP7_75t_L g2431 ( 
.A1(n_2176),
.A2(n_1493),
.B(n_1491),
.Y(n_2431)
);

OAI21x1_ASAP7_75t_L g2432 ( 
.A1(n_2182),
.A2(n_944),
.B(n_940),
.Y(n_2432)
);

AOI21xp5_ASAP7_75t_L g2433 ( 
.A1(n_2176),
.A2(n_1493),
.B(n_1491),
.Y(n_2433)
);

AOI21x1_ASAP7_75t_L g2434 ( 
.A1(n_2136),
.A2(n_946),
.B(n_944),
.Y(n_2434)
);

AOI21xp5_ASAP7_75t_L g2435 ( 
.A1(n_2021),
.A2(n_1493),
.B(n_1491),
.Y(n_2435)
);

OAI21xp33_ASAP7_75t_L g2436 ( 
.A1(n_2083),
.A2(n_561),
.B(n_611),
.Y(n_2436)
);

AOI21x1_ASAP7_75t_L g2437 ( 
.A1(n_2136),
.A2(n_946),
.B(n_661),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2095),
.Y(n_2438)
);

OAI21xp33_ASAP7_75t_L g2439 ( 
.A1(n_2083),
.A2(n_620),
.B(n_617),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2119),
.Y(n_2440)
);

BUFx6f_ASAP7_75t_L g2441 ( 
.A(n_2219),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2183),
.B(n_1688),
.Y(n_2442)
);

AOI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2021),
.A2(n_1515),
.B(n_1493),
.Y(n_2443)
);

OAI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_2219),
.A2(n_1724),
.B1(n_1736),
.B2(n_1695),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_SL g2445 ( 
.A(n_2088),
.B(n_1695),
.Y(n_2445)
);

OAI21x1_ASAP7_75t_SL g2446 ( 
.A1(n_2201),
.A2(n_2204),
.B(n_2202),
.Y(n_2446)
);

AOI221xp5_ASAP7_75t_L g2447 ( 
.A1(n_2077),
.A2(n_674),
.B1(n_678),
.B2(n_665),
.C(n_655),
.Y(n_2447)
);

AOI21xp5_ASAP7_75t_L g2448 ( 
.A1(n_2056),
.A2(n_1515),
.B(n_1493),
.Y(n_2448)
);

OAI22x1_ASAP7_75t_L g2449 ( 
.A1(n_2243),
.A2(n_674),
.B1(n_678),
.B2(n_665),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_2088),
.B(n_1695),
.Y(n_2450)
);

AOI21xp5_ASAP7_75t_L g2451 ( 
.A1(n_2056),
.A2(n_1515),
.B(n_1724),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_2110),
.B(n_1724),
.Y(n_2452)
);

AND2x4_ASAP7_75t_L g2453 ( 
.A(n_2096),
.B(n_1736),
.Y(n_2453)
);

OAI21x1_ASAP7_75t_SL g2454 ( 
.A1(n_2205),
.A2(n_681),
.B(n_679),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_SL g2455 ( 
.A(n_2110),
.B(n_1736),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2207),
.B(n_1688),
.Y(n_2456)
);

AOI21xp5_ASAP7_75t_L g2457 ( 
.A1(n_2210),
.A2(n_1515),
.B(n_1736),
.Y(n_2457)
);

AOI21xp5_ASAP7_75t_L g2458 ( 
.A1(n_2210),
.A2(n_1515),
.B(n_1743),
.Y(n_2458)
);

OAI21xp33_ASAP7_75t_L g2459 ( 
.A1(n_2180),
.A2(n_2216),
.B(n_2213),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2208),
.B(n_1688),
.Y(n_2460)
);

OAI21x1_ASAP7_75t_SL g2461 ( 
.A1(n_2209),
.A2(n_681),
.B(n_679),
.Y(n_2461)
);

BUFx4f_ASAP7_75t_L g2462 ( 
.A(n_2068),
.Y(n_2462)
);

INVx5_ASAP7_75t_L g2463 ( 
.A(n_2133),
.Y(n_2463)
);

AOI21xp5_ASAP7_75t_L g2464 ( 
.A1(n_2212),
.A2(n_1745),
.B(n_1743),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_2215),
.B(n_1730),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2220),
.B(n_1730),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2226),
.B(n_1730),
.Y(n_2467)
);

OAI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2124),
.A2(n_1757),
.B(n_697),
.Y(n_2468)
);

AOI21x1_ASAP7_75t_L g2469 ( 
.A1(n_2239),
.A2(n_697),
.B(n_685),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_2189),
.Y(n_2470)
);

A2O1A1Ixp33_ASAP7_75t_L g2471 ( 
.A1(n_2180),
.A2(n_2213),
.B(n_2216),
.C(n_2033),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_2105),
.B(n_704),
.Y(n_2472)
);

A2O1A1Ixp33_ASAP7_75t_L g2473 ( 
.A1(n_2143),
.A2(n_698),
.B(n_703),
.C(n_685),
.Y(n_2473)
);

BUFx2_ASAP7_75t_L g2474 ( 
.A(n_2166),
.Y(n_2474)
);

AOI21xp5_ASAP7_75t_L g2475 ( 
.A1(n_2212),
.A2(n_1751),
.B(n_1743),
.Y(n_2475)
);

NAND2xp33_ASAP7_75t_L g2476 ( 
.A(n_2035),
.B(n_1743),
.Y(n_2476)
);

A2O1A1Ixp33_ASAP7_75t_L g2477 ( 
.A1(n_2143),
.A2(n_703),
.B(n_705),
.C(n_698),
.Y(n_2477)
);

BUFx2_ASAP7_75t_L g2478 ( 
.A(n_2049),
.Y(n_2478)
);

INVxp67_ASAP7_75t_L g2479 ( 
.A(n_2075),
.Y(n_2479)
);

AO31x2_ASAP7_75t_L g2480 ( 
.A1(n_2228),
.A2(n_712),
.A3(n_718),
.B(n_705),
.Y(n_2480)
);

A2O1A1Ixp33_ASAP7_75t_L g2481 ( 
.A1(n_2194),
.A2(n_718),
.B(n_721),
.C(n_712),
.Y(n_2481)
);

O2A1O1Ixp33_ASAP7_75t_L g2482 ( 
.A1(n_2103),
.A2(n_722),
.B(n_724),
.C(n_721),
.Y(n_2482)
);

AO21x1_ASAP7_75t_L g2483 ( 
.A1(n_2229),
.A2(n_724),
.B(n_722),
.Y(n_2483)
);

AOI21xp5_ASAP7_75t_L g2484 ( 
.A1(n_2234),
.A2(n_1765),
.B(n_1751),
.Y(n_2484)
);

AOI21x1_ASAP7_75t_L g2485 ( 
.A1(n_2230),
.A2(n_729),
.B(n_726),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2232),
.Y(n_2486)
);

OAI21xp5_ASAP7_75t_L g2487 ( 
.A1(n_2227),
.A2(n_1757),
.B(n_729),
.Y(n_2487)
);

INVx3_ASAP7_75t_L g2488 ( 
.A(n_2218),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2105),
.B(n_704),
.Y(n_2489)
);

AO31x2_ASAP7_75t_L g2490 ( 
.A1(n_2238),
.A2(n_738),
.A3(n_740),
.B(n_726),
.Y(n_2490)
);

OR2x6_ASAP7_75t_L g2491 ( 
.A(n_2087),
.B(n_1751),
.Y(n_2491)
);

AOI21xp5_ASAP7_75t_L g2492 ( 
.A1(n_2234),
.A2(n_1765),
.B(n_1751),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2244),
.B(n_2245),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2130),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2145),
.B(n_1757),
.Y(n_2495)
);

A2O1A1Ixp33_ASAP7_75t_L g2496 ( 
.A1(n_2194),
.A2(n_740),
.B(n_743),
.C(n_738),
.Y(n_2496)
);

AND2x4_ASAP7_75t_L g2497 ( 
.A(n_2068),
.B(n_1765),
.Y(n_2497)
);

OAI21xp5_ASAP7_75t_L g2498 ( 
.A1(n_2227),
.A2(n_1757),
.B(n_750),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2159),
.B(n_1757),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2084),
.B(n_708),
.Y(n_2500)
);

OAI22xp33_ASAP7_75t_L g2501 ( 
.A1(n_2092),
.A2(n_623),
.B1(n_624),
.B2(n_622),
.Y(n_2501)
);

NAND2x1_ASAP7_75t_L g2502 ( 
.A(n_2087),
.B(n_1765),
.Y(n_2502)
);

OAI21x1_ASAP7_75t_L g2503 ( 
.A1(n_2164),
.A2(n_750),
.B(n_743),
.Y(n_2503)
);

OAI21x1_ASAP7_75t_L g2504 ( 
.A1(n_2190),
.A2(n_763),
.B(n_758),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2191),
.B(n_1770),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2196),
.Y(n_2506)
);

INVxp67_ASAP7_75t_SL g2507 ( 
.A(n_2135),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2199),
.B(n_1770),
.Y(n_2508)
);

OAI21xp5_ASAP7_75t_L g2509 ( 
.A1(n_2198),
.A2(n_2222),
.B(n_2217),
.Y(n_2509)
);

AOI21xp5_ASAP7_75t_L g2510 ( 
.A1(n_2098),
.A2(n_1774),
.B(n_1770),
.Y(n_2510)
);

OAI21x1_ASAP7_75t_L g2511 ( 
.A1(n_2236),
.A2(n_763),
.B(n_758),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2198),
.B(n_1770),
.Y(n_2512)
);

AND2x2_ASAP7_75t_L g2513 ( 
.A(n_2104),
.B(n_708),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2167),
.B(n_1774),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2167),
.B(n_765),
.Y(n_2515)
);

OAI21x1_ASAP7_75t_L g2516 ( 
.A1(n_2135),
.A2(n_768),
.B(n_765),
.Y(n_2516)
);

OAI21x1_ASAP7_75t_L g2517 ( 
.A1(n_2030),
.A2(n_769),
.B(n_768),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2142),
.Y(n_2518)
);

AND2x4_ASAP7_75t_L g2519 ( 
.A(n_2253),
.B(n_2141),
.Y(n_2519)
);

BUFx3_ASAP7_75t_L g2520 ( 
.A(n_2284),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_SL g2521 ( 
.A(n_2270),
.B(n_2160),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2258),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2279),
.Y(n_2523)
);

INVx4_ASAP7_75t_SL g2524 ( 
.A(n_2264),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2298),
.Y(n_2525)
);

AOI22xp33_ASAP7_75t_SL g2526 ( 
.A1(n_2334),
.A2(n_2160),
.B1(n_2036),
.B2(n_2165),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2288),
.B(n_2243),
.Y(n_2527)
);

NAND2x1p5_ASAP7_75t_L g2528 ( 
.A(n_2462),
.B(n_2296),
.Y(n_2528)
);

BUFx6f_ASAP7_75t_L g2529 ( 
.A(n_2284),
.Y(n_2529)
);

INVxp67_ASAP7_75t_SL g2530 ( 
.A(n_2493),
.Y(n_2530)
);

BUFx10_ASAP7_75t_L g2531 ( 
.A(n_2264),
.Y(n_2531)
);

BUFx6f_ASAP7_75t_L g2532 ( 
.A(n_2284),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2419),
.Y(n_2533)
);

BUFx6f_ASAP7_75t_L g2534 ( 
.A(n_2360),
.Y(n_2534)
);

O2A1O1Ixp33_ASAP7_75t_L g2535 ( 
.A1(n_2471),
.A2(n_2482),
.B(n_2347),
.C(n_2265),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2395),
.B(n_2137),
.Y(n_2536)
);

AND2x2_ASAP7_75t_L g2537 ( 
.A(n_2292),
.B(n_2179),
.Y(n_2537)
);

AOI21xp5_ASAP7_75t_L g2538 ( 
.A1(n_2260),
.A2(n_2252),
.B(n_2263),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2315),
.Y(n_2539)
);

INVxp67_ASAP7_75t_L g2540 ( 
.A(n_2303),
.Y(n_2540)
);

AND2x4_ASAP7_75t_L g2541 ( 
.A(n_2253),
.B(n_2200),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_L g2542 ( 
.A(n_2269),
.B(n_2059),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2425),
.Y(n_2543)
);

OAI21xp33_ASAP7_75t_L g2544 ( 
.A1(n_2418),
.A2(n_2447),
.B(n_2396),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2323),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2486),
.Y(n_2546)
);

INVx5_ASAP7_75t_L g2547 ( 
.A(n_2429),
.Y(n_2547)
);

AND2x4_ASAP7_75t_L g2548 ( 
.A(n_2343),
.B(n_2053),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_L g2549 ( 
.A(n_2479),
.B(n_2241),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2287),
.Y(n_2550)
);

AOI21xp33_ASAP7_75t_L g2551 ( 
.A1(n_2374),
.A2(n_2230),
.B(n_2087),
.Y(n_2551)
);

INVx1_ASAP7_75t_SL g2552 ( 
.A(n_2250),
.Y(n_2552)
);

AOI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2459),
.A2(n_2070),
.B1(n_2036),
.B2(n_2098),
.Y(n_2553)
);

BUFx2_ASAP7_75t_L g2554 ( 
.A(n_2379),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2330),
.Y(n_2555)
);

AOI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2316),
.A2(n_2098),
.B1(n_627),
.B2(n_632),
.Y(n_2556)
);

INVx2_ASAP7_75t_SL g2557 ( 
.A(n_2360),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2297),
.Y(n_2558)
);

OAI21xp33_ASAP7_75t_L g2559 ( 
.A1(n_2447),
.A2(n_638),
.B(n_626),
.Y(n_2559)
);

O2A1O1Ixp5_ASAP7_75t_L g2560 ( 
.A1(n_2252),
.A2(n_778),
.B(n_783),
.C(n_769),
.Y(n_2560)
);

INVx2_ASAP7_75t_SL g2561 ( 
.A(n_2360),
.Y(n_2561)
);

NOR2x1_ASAP7_75t_SL g2562 ( 
.A(n_2463),
.B(n_2230),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_2401),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2273),
.B(n_2142),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2346),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_R g2566 ( 
.A(n_2257),
.B(n_2025),
.Y(n_2566)
);

OAI22xp5_ASAP7_75t_L g2567 ( 
.A1(n_2288),
.A2(n_2148),
.B1(n_787),
.B2(n_793),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2361),
.B(n_2142),
.Y(n_2568)
);

BUFx5_ASAP7_75t_L g2569 ( 
.A(n_2247),
.Y(n_2569)
);

AOI22xp5_ASAP7_75t_L g2570 ( 
.A1(n_2274),
.A2(n_642),
.B1(n_643),
.B2(n_641),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_2462),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2387),
.B(n_2197),
.Y(n_2572)
);

AOI22xp5_ASAP7_75t_L g2573 ( 
.A1(n_2274),
.A2(n_646),
.B1(n_649),
.B2(n_645),
.Y(n_2573)
);

INVx2_ASAP7_75t_SL g2574 ( 
.A(n_2410),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2364),
.Y(n_2575)
);

OAI22xp5_ASAP7_75t_L g2576 ( 
.A1(n_2387),
.A2(n_2372),
.B1(n_2251),
.B2(n_2261),
.Y(n_2576)
);

AOI21xp5_ASAP7_75t_L g2577 ( 
.A1(n_2260),
.A2(n_2030),
.B(n_2197),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2251),
.B(n_2197),
.Y(n_2578)
);

OAI221xp5_ASAP7_75t_L g2579 ( 
.A1(n_2439),
.A2(n_793),
.B1(n_778),
.B2(n_653),
.C(n_656),
.Y(n_2579)
);

BUFx4f_ASAP7_75t_SL g2580 ( 
.A(n_2410),
.Y(n_2580)
);

AOI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2313),
.A2(n_2043),
.B(n_2025),
.Y(n_2581)
);

BUFx8_ASAP7_75t_SL g2582 ( 
.A(n_2406),
.Y(n_2582)
);

BUFx6f_ASAP7_75t_L g2583 ( 
.A(n_2441),
.Y(n_2583)
);

BUFx3_ASAP7_75t_L g2584 ( 
.A(n_2336),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2381),
.Y(n_2585)
);

INVx3_ASAP7_75t_L g2586 ( 
.A(n_2383),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2365),
.B(n_2025),
.Y(n_2587)
);

AND2x6_ASAP7_75t_L g2588 ( 
.A(n_2409),
.B(n_2246),
.Y(n_2588)
);

HB1xp67_ASAP7_75t_L g2589 ( 
.A(n_2386),
.Y(n_2589)
);

AOI22xp5_ASAP7_75t_L g2590 ( 
.A1(n_2449),
.A2(n_652),
.B1(n_659),
.B2(n_651),
.Y(n_2590)
);

BUFx6f_ASAP7_75t_L g2591 ( 
.A(n_2441),
.Y(n_2591)
);

NAND2x1_ASAP7_75t_L g2592 ( 
.A(n_2416),
.B(n_2133),
.Y(n_2592)
);

INVxp67_ASAP7_75t_SL g2593 ( 
.A(n_2493),
.Y(n_2593)
);

A2O1A1Ixp33_ASAP7_75t_L g2594 ( 
.A1(n_2357),
.A2(n_2148),
.B(n_667),
.C(n_672),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2353),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2402),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2411),
.Y(n_2597)
);

INVx1_ASAP7_75t_SL g2598 ( 
.A(n_2259),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2365),
.B(n_2043),
.Y(n_2599)
);

BUFx2_ASAP7_75t_L g2600 ( 
.A(n_2428),
.Y(n_2600)
);

NOR2x1_ASAP7_75t_L g2601 ( 
.A(n_2261),
.B(n_2246),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2295),
.B(n_2043),
.Y(n_2602)
);

AND2x4_ASAP7_75t_L g2603 ( 
.A(n_2491),
.B(n_2262),
.Y(n_2603)
);

AOI21xp5_ASAP7_75t_L g2604 ( 
.A1(n_2314),
.A2(n_2086),
.B(n_2081),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2370),
.Y(n_2605)
);

OR2x6_ASAP7_75t_L g2606 ( 
.A(n_2254),
.B(n_2246),
.Y(n_2606)
);

BUFx6f_ASAP7_75t_L g2607 ( 
.A(n_2441),
.Y(n_2607)
);

NAND3xp33_ASAP7_75t_L g2608 ( 
.A(n_2325),
.B(n_676),
.C(n_662),
.Y(n_2608)
);

BUFx2_ASAP7_75t_L g2609 ( 
.A(n_2390),
.Y(n_2609)
);

BUFx2_ASAP7_75t_L g2610 ( 
.A(n_2421),
.Y(n_2610)
);

BUFx2_ASAP7_75t_L g2611 ( 
.A(n_2421),
.Y(n_2611)
);

NOR2xp33_ASAP7_75t_L g2612 ( 
.A(n_2271),
.B(n_677),
.Y(n_2612)
);

AOI21xp5_ASAP7_75t_L g2613 ( 
.A1(n_2311),
.A2(n_2086),
.B(n_2081),
.Y(n_2613)
);

AND2x4_ASAP7_75t_L g2614 ( 
.A(n_2491),
.B(n_2081),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2399),
.Y(n_2615)
);

OR2x2_ASAP7_75t_L g2616 ( 
.A(n_2515),
.B(n_2086),
.Y(n_2616)
);

AND2x4_ASAP7_75t_L g2617 ( 
.A(n_2491),
.B(n_2101),
.Y(n_2617)
);

BUFx6f_ASAP7_75t_L g2618 ( 
.A(n_2478),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2325),
.A2(n_684),
.B1(n_687),
.B2(n_683),
.Y(n_2619)
);

BUFx6f_ASAP7_75t_L g2620 ( 
.A(n_2383),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2446),
.Y(n_2621)
);

O2A1O1Ixp5_ASAP7_75t_L g2622 ( 
.A1(n_2445),
.A2(n_2218),
.B(n_2133),
.C(n_2188),
.Y(n_2622)
);

AND2x4_ASAP7_75t_L g2623 ( 
.A(n_2262),
.B(n_2497),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2278),
.B(n_2101),
.Y(n_2624)
);

INVx2_ASAP7_75t_SL g2625 ( 
.A(n_2264),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2285),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2285),
.Y(n_2627)
);

INVx3_ASAP7_75t_SL g2628 ( 
.A(n_2289),
.Y(n_2628)
);

CKINVDCx11_ASAP7_75t_R g2629 ( 
.A(n_2474),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2278),
.B(n_2101),
.Y(n_2630)
);

INVx8_ASAP7_75t_L g2631 ( 
.A(n_2429),
.Y(n_2631)
);

AND2x4_ASAP7_75t_L g2632 ( 
.A(n_2497),
.B(n_2133),
.Y(n_2632)
);

INVx2_ASAP7_75t_SL g2633 ( 
.A(n_2289),
.Y(n_2633)
);

AOI21xp5_ASAP7_75t_L g2634 ( 
.A1(n_2291),
.A2(n_2133),
.B(n_2172),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2407),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2285),
.Y(n_2636)
);

INVx1_ASAP7_75t_SL g2637 ( 
.A(n_2348),
.Y(n_2637)
);

INVx6_ASAP7_75t_L g2638 ( 
.A(n_2289),
.Y(n_2638)
);

INVx2_ASAP7_75t_SL g2639 ( 
.A(n_2400),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2438),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2440),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2335),
.Y(n_2642)
);

OR2x6_ASAP7_75t_L g2643 ( 
.A(n_2317),
.B(n_2109),
.Y(n_2643)
);

BUFx6f_ASAP7_75t_L g2644 ( 
.A(n_2296),
.Y(n_2644)
);

AND2x4_ASAP7_75t_L g2645 ( 
.A(n_2426),
.B(n_2037),
.Y(n_2645)
);

AOI21xp5_ASAP7_75t_L g2646 ( 
.A1(n_2299),
.A2(n_2181),
.B(n_2184),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2283),
.B(n_688),
.Y(n_2647)
);

AOI21xp5_ASAP7_75t_L g2648 ( 
.A1(n_2305),
.A2(n_2307),
.B(n_2276),
.Y(n_2648)
);

INVxp67_ASAP7_75t_SL g2649 ( 
.A(n_2312),
.Y(n_2649)
);

INVx3_ASAP7_75t_L g2650 ( 
.A(n_2392),
.Y(n_2650)
);

AND2x4_ASAP7_75t_L g2651 ( 
.A(n_2426),
.B(n_373),
.Y(n_2651)
);

AND2x4_ASAP7_75t_L g2652 ( 
.A(n_2453),
.B(n_377),
.Y(n_2652)
);

INVx3_ASAP7_75t_R g2653 ( 
.A(n_2388),
.Y(n_2653)
);

HB1xp67_ASAP7_75t_L g2654 ( 
.A(n_2512),
.Y(n_2654)
);

NOR2xp67_ASAP7_75t_SL g2655 ( 
.A(n_2463),
.B(n_691),
.Y(n_2655)
);

INVx2_ASAP7_75t_SL g2656 ( 
.A(n_2392),
.Y(n_2656)
);

INVx3_ASAP7_75t_L g2657 ( 
.A(n_2321),
.Y(n_2657)
);

AND2x4_ASAP7_75t_L g2658 ( 
.A(n_2453),
.B(n_378),
.Y(n_2658)
);

INVx2_ASAP7_75t_SL g2659 ( 
.A(n_2518),
.Y(n_2659)
);

BUFx6f_ASAP7_75t_L g2660 ( 
.A(n_2321),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2335),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_SL g2662 ( 
.A(n_2357),
.B(n_708),
.Y(n_2662)
);

BUFx3_ASAP7_75t_L g2663 ( 
.A(n_2371),
.Y(n_2663)
);

AND2x4_ASAP7_75t_L g2664 ( 
.A(n_2470),
.B(n_381),
.Y(n_2664)
);

BUFx6f_ASAP7_75t_L g2665 ( 
.A(n_2371),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2283),
.B(n_695),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2335),
.Y(n_2667)
);

CKINVDCx5p33_ASAP7_75t_R g2668 ( 
.A(n_2373),
.Y(n_2668)
);

CKINVDCx11_ASAP7_75t_R g2669 ( 
.A(n_2494),
.Y(n_2669)
);

CKINVDCx6p67_ASAP7_75t_R g2670 ( 
.A(n_2513),
.Y(n_2670)
);

INVx3_ASAP7_75t_L g2671 ( 
.A(n_2416),
.Y(n_2671)
);

INVx3_ASAP7_75t_L g2672 ( 
.A(n_2416),
.Y(n_2672)
);

INVx2_ASAP7_75t_SL g2673 ( 
.A(n_2393),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_L g2674 ( 
.A(n_2500),
.B(n_699),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2338),
.Y(n_2675)
);

INVx3_ASAP7_75t_L g2676 ( 
.A(n_2470),
.Y(n_2676)
);

AOI22xp5_ASAP7_75t_L g2677 ( 
.A1(n_2368),
.A2(n_710),
.B1(n_713),
.B2(n_707),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_SL g2678 ( 
.A(n_2281),
.B(n_708),
.Y(n_2678)
);

BUFx2_ASAP7_75t_L g2679 ( 
.A(n_2488),
.Y(n_2679)
);

BUFx2_ASAP7_75t_L g2680 ( 
.A(n_2488),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2363),
.B(n_714),
.Y(n_2681)
);

OA21x2_ASAP7_75t_L g2682 ( 
.A1(n_2248),
.A2(n_717),
.B(n_716),
.Y(n_2682)
);

INVx1_ASAP7_75t_SL g2683 ( 
.A(n_2512),
.Y(n_2683)
);

AOI22xp5_ASAP7_75t_L g2684 ( 
.A1(n_2436),
.A2(n_719),
.B1(n_725),
.B2(n_723),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2480),
.Y(n_2685)
);

OR2x6_ASAP7_75t_L g2686 ( 
.A(n_2412),
.B(n_986),
.Y(n_2686)
);

AND2x6_ASAP7_75t_L g2687 ( 
.A(n_2376),
.B(n_1009),
.Y(n_2687)
);

AOI21xp5_ASAP7_75t_L g2688 ( 
.A1(n_2463),
.A2(n_1107),
.B(n_1084),
.Y(n_2688)
);

AOI21xp5_ASAP7_75t_L g2689 ( 
.A1(n_2463),
.A2(n_1110),
.B(n_1107),
.Y(n_2689)
);

BUFx3_ASAP7_75t_L g2690 ( 
.A(n_2472),
.Y(n_2690)
);

OR2x2_ASAP7_75t_L g2691 ( 
.A(n_2515),
.B(n_2),
.Y(n_2691)
);

NOR2xp33_ASAP7_75t_L g2692 ( 
.A(n_2501),
.B(n_728),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2480),
.Y(n_2693)
);

BUFx8_ASAP7_75t_SL g2694 ( 
.A(n_2489),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2294),
.B(n_732),
.Y(n_2695)
);

INVx1_ASAP7_75t_SL g2696 ( 
.A(n_2356),
.Y(n_2696)
);

INVx3_ASAP7_75t_L g2697 ( 
.A(n_2413),
.Y(n_2697)
);

INVx3_ASAP7_75t_L g2698 ( 
.A(n_2502),
.Y(n_2698)
);

AOI21xp5_ASAP7_75t_L g2699 ( 
.A1(n_2318),
.A2(n_1110),
.B(n_1107),
.Y(n_2699)
);

BUFx2_ASAP7_75t_L g2700 ( 
.A(n_2507),
.Y(n_2700)
);

OR2x2_ASAP7_75t_L g2701 ( 
.A(n_2480),
.B(n_3),
.Y(n_2701)
);

AOI22xp33_ASAP7_75t_L g2702 ( 
.A1(n_2362),
.A2(n_753),
.B1(n_714),
.B2(n_739),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2506),
.Y(n_2703)
);

INVx8_ASAP7_75t_L g2704 ( 
.A(n_2429),
.Y(n_2704)
);

INVx5_ASAP7_75t_L g2705 ( 
.A(n_2429),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2294),
.B(n_733),
.Y(n_2706)
);

BUFx6f_ASAP7_75t_L g2707 ( 
.A(n_2417),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2505),
.Y(n_2708)
);

INVx2_ASAP7_75t_SL g2709 ( 
.A(n_2514),
.Y(n_2709)
);

AOI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2384),
.A2(n_741),
.B1(n_746),
.B2(n_742),
.Y(n_2710)
);

OR2x6_ASAP7_75t_L g2711 ( 
.A(n_2272),
.B(n_986),
.Y(n_2711)
);

BUFx6f_ASAP7_75t_L g2712 ( 
.A(n_2306),
.Y(n_2712)
);

CKINVDCx5p33_ASAP7_75t_R g2713 ( 
.A(n_2514),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2490),
.Y(n_2714)
);

HB1xp67_ASAP7_75t_L g2715 ( 
.A(n_2509),
.Y(n_2715)
);

INVx5_ASAP7_75t_L g2716 ( 
.A(n_2247),
.Y(n_2716)
);

INVx3_ASAP7_75t_L g2717 ( 
.A(n_2306),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2312),
.B(n_747),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2490),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2358),
.Y(n_2720)
);

OR2x2_ASAP7_75t_L g2721 ( 
.A(n_2490),
.B(n_4),
.Y(n_2721)
);

OAI22xp5_ASAP7_75t_L g2722 ( 
.A1(n_2481),
.A2(n_748),
.B1(n_755),
.B2(n_754),
.Y(n_2722)
);

HB1xp67_ASAP7_75t_L g2723 ( 
.A(n_2509),
.Y(n_2723)
);

INVxp67_ASAP7_75t_L g2724 ( 
.A(n_2322),
.Y(n_2724)
);

AND2x4_ASAP7_75t_L g2725 ( 
.A(n_2430),
.B(n_382),
.Y(n_2725)
);

O2A1O1Ixp5_ASAP7_75t_SL g2726 ( 
.A1(n_2275),
.A2(n_753),
.B(n_714),
.C(n_757),
.Y(n_2726)
);

INVx4_ASAP7_75t_L g2727 ( 
.A(n_2358),
.Y(n_2727)
);

BUFx6f_ASAP7_75t_L g2728 ( 
.A(n_2247),
.Y(n_2728)
);

AO31x2_ASAP7_75t_L g2729 ( 
.A1(n_2404),
.A2(n_1058),
.A3(n_390),
.B(n_391),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2267),
.Y(n_2730)
);

NOR3xp33_ASAP7_75t_L g2731 ( 
.A(n_2350),
.B(n_761),
.C(n_760),
.Y(n_2731)
);

AND2x4_ASAP7_75t_L g2732 ( 
.A(n_2430),
.B(n_383),
.Y(n_2732)
);

AOI22xp33_ASAP7_75t_L g2733 ( 
.A1(n_2275),
.A2(n_753),
.B1(n_714),
.B2(n_762),
.Y(n_2733)
);

AOI22xp5_ASAP7_75t_L g2734 ( 
.A1(n_2483),
.A2(n_766),
.B1(n_770),
.B2(n_767),
.Y(n_2734)
);

NOR2xp33_ASAP7_75t_L g2735 ( 
.A(n_2382),
.B(n_2450),
.Y(n_2735)
);

BUFx6f_ASAP7_75t_L g2736 ( 
.A(n_2247),
.Y(n_2736)
);

AOI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2282),
.A2(n_1110),
.B(n_1107),
.Y(n_2737)
);

INVx3_ASAP7_75t_L g2738 ( 
.A(n_2266),
.Y(n_2738)
);

BUFx3_ASAP7_75t_L g2739 ( 
.A(n_2266),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2322),
.B(n_774),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2300),
.B(n_779),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2300),
.B(n_780),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2267),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2352),
.B(n_785),
.Y(n_2744)
);

OAI22xp5_ASAP7_75t_L g2745 ( 
.A1(n_2496),
.A2(n_790),
.B1(n_794),
.B2(n_792),
.Y(n_2745)
);

OAI22xp5_ASAP7_75t_SL g2746 ( 
.A1(n_2468),
.A2(n_753),
.B1(n_8),
.B2(n_5),
.Y(n_2746)
);

BUFx6f_ASAP7_75t_L g2747 ( 
.A(n_2485),
.Y(n_2747)
);

AOI21xp5_ASAP7_75t_L g2748 ( 
.A1(n_2290),
.A2(n_1110),
.B(n_1107),
.Y(n_2748)
);

INVx3_ASAP7_75t_L g2749 ( 
.A(n_2256),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2473),
.B(n_394),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2352),
.B(n_7),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2376),
.B(n_7),
.Y(n_2752)
);

AOI22xp5_ASAP7_75t_L g2753 ( 
.A1(n_2422),
.A2(n_1033),
.B1(n_1055),
.B2(n_1016),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2505),
.Y(n_2754)
);

OR2x2_ASAP7_75t_L g2755 ( 
.A(n_2380),
.B(n_2391),
.Y(n_2755)
);

INVx1_ASAP7_75t_SL g2756 ( 
.A(n_2380),
.Y(n_2756)
);

AOI22xp33_ASAP7_75t_L g2757 ( 
.A1(n_2454),
.A2(n_986),
.B1(n_1055),
.B2(n_1033),
.Y(n_2757)
);

O2A1O1Ixp5_ASAP7_75t_L g2758 ( 
.A1(n_2452),
.A2(n_1058),
.B(n_10),
.C(n_8),
.Y(n_2758)
);

AND2x4_ASAP7_75t_L g2759 ( 
.A(n_2510),
.B(n_397),
.Y(n_2759)
);

INVx3_ASAP7_75t_L g2760 ( 
.A(n_2255),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2267),
.Y(n_2761)
);

AOI21xp5_ASAP7_75t_L g2762 ( 
.A1(n_2327),
.A2(n_1117),
.B(n_1110),
.Y(n_2762)
);

O2A1O1Ixp5_ASAP7_75t_L g2763 ( 
.A1(n_2455),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2301),
.Y(n_2764)
);

INVx2_ASAP7_75t_SL g2765 ( 
.A(n_2508),
.Y(n_2765)
);

INVx3_ASAP7_75t_L g2766 ( 
.A(n_2268),
.Y(n_2766)
);

AOI21xp5_ASAP7_75t_L g2767 ( 
.A1(n_2331),
.A2(n_1119),
.B(n_1117),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2286),
.Y(n_2768)
);

AOI21x1_ASAP7_75t_L g2769 ( 
.A1(n_2434),
.A2(n_1119),
.B(n_1117),
.Y(n_2769)
);

CKINVDCx20_ASAP7_75t_R g2770 ( 
.A(n_2391),
.Y(n_2770)
);

BUFx4f_ASAP7_75t_SL g2771 ( 
.A(n_2476),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2355),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2423),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2508),
.Y(n_2774)
);

BUFx3_ASAP7_75t_L g2775 ( 
.A(n_2461),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_2444),
.Y(n_2776)
);

BUFx3_ASAP7_75t_L g2777 ( 
.A(n_2516),
.Y(n_2777)
);

OAI22xp5_ASAP7_75t_SL g2778 ( 
.A1(n_2468),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_2778)
);

OAI22xp5_ASAP7_75t_L g2779 ( 
.A1(n_2477),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_2779)
);

NOR2x1p5_ASAP7_75t_L g2780 ( 
.A(n_2469),
.B(n_986),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2432),
.Y(n_2781)
);

BUFx6f_ASAP7_75t_L g2782 ( 
.A(n_2277),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2345),
.Y(n_2783)
);

INVxp67_ASAP7_75t_L g2784 ( 
.A(n_2397),
.Y(n_2784)
);

OR2x2_ASAP7_75t_L g2785 ( 
.A(n_2397),
.B(n_14),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2522),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2523),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2533),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2543),
.Y(n_2789)
);

OAI21xp5_ASAP7_75t_L g2790 ( 
.A1(n_2608),
.A2(n_2377),
.B(n_2319),
.Y(n_2790)
);

BUFx4f_ASAP7_75t_L g2791 ( 
.A(n_2583),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2546),
.Y(n_2792)
);

AOI22xp33_ASAP7_75t_L g2793 ( 
.A1(n_2544),
.A2(n_2332),
.B1(n_2302),
.B2(n_2422),
.Y(n_2793)
);

BUFx3_ASAP7_75t_L g2794 ( 
.A(n_2529),
.Y(n_2794)
);

OAI21x1_ASAP7_75t_L g2795 ( 
.A1(n_2648),
.A2(n_2367),
.B(n_2369),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2550),
.Y(n_2796)
);

CKINVDCx20_ASAP7_75t_R g2797 ( 
.A(n_2629),
.Y(n_2797)
);

BUFx3_ASAP7_75t_L g2798 ( 
.A(n_2529),
.Y(n_2798)
);

OAI21x1_ASAP7_75t_L g2799 ( 
.A1(n_2699),
.A2(n_2737),
.B(n_2762),
.Y(n_2799)
);

INVx3_ASAP7_75t_L g2800 ( 
.A(n_2676),
.Y(n_2800)
);

NAND2x1p5_ASAP7_75t_L g2801 ( 
.A(n_2716),
.B(n_2341),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2558),
.Y(n_2802)
);

OAI21x1_ASAP7_75t_SL g2803 ( 
.A1(n_2535),
.A2(n_2359),
.B(n_2420),
.Y(n_2803)
);

OAI21x1_ASAP7_75t_L g2804 ( 
.A1(n_2767),
.A2(n_2538),
.B(n_2769),
.Y(n_2804)
);

AO21x2_ASAP7_75t_L g2805 ( 
.A1(n_2685),
.A2(n_2293),
.B(n_2342),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2575),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2585),
.Y(n_2807)
);

OAI21x1_ASAP7_75t_L g2808 ( 
.A1(n_2766),
.A2(n_2333),
.B(n_2366),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2596),
.Y(n_2809)
);

OAI21x1_ASAP7_75t_L g2810 ( 
.A1(n_2766),
.A2(n_2310),
.B(n_2280),
.Y(n_2810)
);

OAI21x1_ASAP7_75t_L g2811 ( 
.A1(n_2577),
.A2(n_2324),
.B(n_2320),
.Y(n_2811)
);

NOR2xp33_ASAP7_75t_L g2812 ( 
.A(n_2576),
.B(n_2527),
.Y(n_2812)
);

OAI21xp5_ASAP7_75t_L g2813 ( 
.A1(n_2608),
.A2(n_2308),
.B(n_2349),
.Y(n_2813)
);

AO21x2_ASAP7_75t_L g2814 ( 
.A1(n_2693),
.A2(n_2293),
.B(n_2339),
.Y(n_2814)
);

INVxp67_ASAP7_75t_SL g2815 ( 
.A(n_2715),
.Y(n_2815)
);

NAND2xp33_ASAP7_75t_L g2816 ( 
.A(n_2746),
.B(n_2329),
.Y(n_2816)
);

BUFx6f_ASAP7_75t_L g2817 ( 
.A(n_2529),
.Y(n_2817)
);

OAI21xp5_ASAP7_75t_L g2818 ( 
.A1(n_2619),
.A2(n_2517),
.B(n_2332),
.Y(n_2818)
);

INVx1_ASAP7_75t_SL g2819 ( 
.A(n_2600),
.Y(n_2819)
);

OR2x2_ASAP7_75t_L g2820 ( 
.A(n_2755),
.B(n_2249),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2597),
.Y(n_2821)
);

BUFx2_ASAP7_75t_R g2822 ( 
.A(n_2582),
.Y(n_2822)
);

OAI21x1_ASAP7_75t_L g2823 ( 
.A1(n_2768),
.A2(n_2783),
.B(n_2661),
.Y(n_2823)
);

OR2x2_ASAP7_75t_L g2824 ( 
.A(n_2756),
.B(n_2249),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2654),
.Y(n_2825)
);

AO21x2_ASAP7_75t_L g2826 ( 
.A1(n_2714),
.A2(n_2719),
.B(n_2730),
.Y(n_2826)
);

AND2x2_ASAP7_75t_L g2827 ( 
.A(n_2536),
.B(n_2249),
.Y(n_2827)
);

NOR2xp33_ASAP7_75t_L g2828 ( 
.A(n_2576),
.B(n_2437),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2530),
.Y(n_2829)
);

BUFx2_ASAP7_75t_L g2830 ( 
.A(n_2566),
.Y(n_2830)
);

OR2x6_ASAP7_75t_L g2831 ( 
.A(n_2631),
.B(n_2464),
.Y(n_2831)
);

OAI21x1_ASAP7_75t_L g2832 ( 
.A1(n_2642),
.A2(n_2414),
.B(n_2408),
.Y(n_2832)
);

BUFx3_ASAP7_75t_L g2833 ( 
.A(n_2532),
.Y(n_2833)
);

AOI221xp5_ASAP7_75t_L g2834 ( 
.A1(n_2746),
.A2(n_2487),
.B1(n_2498),
.B2(n_2302),
.C(n_2359),
.Y(n_2834)
);

OAI21x1_ASAP7_75t_L g2835 ( 
.A1(n_2748),
.A2(n_2415),
.B(n_2326),
.Y(n_2835)
);

OAI21x1_ASAP7_75t_L g2836 ( 
.A1(n_2667),
.A2(n_2634),
.B(n_2760),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2593),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2703),
.Y(n_2838)
);

OR2x6_ASAP7_75t_L g2839 ( 
.A(n_2631),
.B(n_2464),
.Y(n_2839)
);

AND2x4_ASAP7_75t_L g2840 ( 
.A(n_2606),
.B(n_2339),
.Y(n_2840)
);

AOI31xp33_ASAP7_75t_SL g2841 ( 
.A1(n_2701),
.A2(n_2424),
.A3(n_2433),
.B(n_2431),
.Y(n_2841)
);

CKINVDCx20_ASAP7_75t_R g2842 ( 
.A(n_2580),
.Y(n_2842)
);

NOR2xp33_ASAP7_75t_L g2843 ( 
.A(n_2619),
.B(n_2442),
.Y(n_2843)
);

OAI21x1_ASAP7_75t_L g2844 ( 
.A1(n_2760),
.A2(n_2781),
.B(n_2764),
.Y(n_2844)
);

OR2x6_ASAP7_75t_L g2845 ( 
.A(n_2631),
.B(n_2704),
.Y(n_2845)
);

OAI21x1_ASAP7_75t_L g2846 ( 
.A1(n_2626),
.A2(n_2309),
.B(n_2304),
.Y(n_2846)
);

OAI21x1_ASAP7_75t_L g2847 ( 
.A1(n_2627),
.A2(n_2344),
.B(n_2340),
.Y(n_2847)
);

CKINVDCx5p33_ASAP7_75t_R g2848 ( 
.A(n_2563),
.Y(n_2848)
);

OAI21x1_ASAP7_75t_L g2849 ( 
.A1(n_2636),
.A2(n_2344),
.B(n_2340),
.Y(n_2849)
);

AO21x2_ASAP7_75t_L g2850 ( 
.A1(n_2743),
.A2(n_2420),
.B(n_2337),
.Y(n_2850)
);

OAI21x1_ASAP7_75t_L g2851 ( 
.A1(n_2613),
.A2(n_2773),
.B(n_2604),
.Y(n_2851)
);

INVx3_ASAP7_75t_L g2852 ( 
.A(n_2676),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2683),
.Y(n_2853)
);

OR2x2_ASAP7_75t_L g2854 ( 
.A(n_2756),
.B(n_2341),
.Y(n_2854)
);

NOR2xp33_ASAP7_75t_L g2855 ( 
.A(n_2752),
.B(n_2442),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2683),
.Y(n_2856)
);

OAI21x1_ASAP7_75t_L g2857 ( 
.A1(n_2581),
.A2(n_2394),
.B(n_2328),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2605),
.Y(n_2858)
);

AOI22xp33_ASAP7_75t_L g2859 ( 
.A1(n_2544),
.A2(n_2487),
.B1(n_2498),
.B2(n_2337),
.Y(n_2859)
);

CKINVDCx6p67_ASAP7_75t_R g2860 ( 
.A(n_2628),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2782),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2782),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2649),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2723),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2621),
.Y(n_2865)
);

BUFx6f_ASAP7_75t_L g2866 ( 
.A(n_2532),
.Y(n_2866)
);

AND2x4_ASAP7_75t_L g2867 ( 
.A(n_2606),
.B(n_2562),
.Y(n_2867)
);

AO21x2_ASAP7_75t_L g2868 ( 
.A1(n_2761),
.A2(n_2427),
.B(n_2378),
.Y(n_2868)
);

AOI21x1_ASAP7_75t_L g2869 ( 
.A1(n_2678),
.A2(n_2375),
.B(n_2354),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2782),
.Y(n_2870)
);

NAND2x1p5_ASAP7_75t_L g2871 ( 
.A(n_2716),
.B(n_2503),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2784),
.Y(n_2872)
);

AOI22xp33_ASAP7_75t_L g2873 ( 
.A1(n_2778),
.A2(n_2511),
.B1(n_2504),
.B2(n_2460),
.Y(n_2873)
);

INVx3_ASAP7_75t_SL g2874 ( 
.A(n_2668),
.Y(n_2874)
);

BUFx2_ASAP7_75t_L g2875 ( 
.A(n_2554),
.Y(n_2875)
);

OAI22xp5_ASAP7_75t_SL g2876 ( 
.A1(n_2653),
.A2(n_2427),
.B1(n_2444),
.B2(n_2456),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2637),
.B(n_2456),
.Y(n_2877)
);

NOR2xp67_ASAP7_75t_L g2878 ( 
.A(n_2671),
.B(n_2351),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2708),
.Y(n_2879)
);

INVx1_ASAP7_75t_SL g2880 ( 
.A(n_2609),
.Y(n_2880)
);

OAI21x1_ASAP7_75t_L g2881 ( 
.A1(n_2749),
.A2(n_2389),
.B(n_2378),
.Y(n_2881)
);

O2A1O1Ixp33_ASAP7_75t_L g2882 ( 
.A1(n_2594),
.A2(n_2460),
.B(n_2466),
.C(n_2465),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_L g2883 ( 
.A(n_2735),
.B(n_2465),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2589),
.Y(n_2884)
);

BUFx2_ASAP7_75t_SL g2885 ( 
.A(n_2584),
.Y(n_2885)
);

OAI21x1_ASAP7_75t_SL g2886 ( 
.A1(n_2567),
.A2(n_2467),
.B(n_2466),
.Y(n_2886)
);

AOI221xp5_ASAP7_75t_L g2887 ( 
.A1(n_2778),
.A2(n_2467),
.B1(n_2499),
.B2(n_2495),
.C(n_2492),
.Y(n_2887)
);

OA21x2_ASAP7_75t_L g2888 ( 
.A1(n_2560),
.A2(n_2403),
.B(n_2405),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2754),
.Y(n_2889)
);

OR2x6_ASAP7_75t_L g2890 ( 
.A(n_2704),
.B(n_2475),
.Y(n_2890)
);

CKINVDCx5p33_ASAP7_75t_R g2891 ( 
.A(n_2694),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2564),
.B(n_2495),
.Y(n_2892)
);

INVx2_ASAP7_75t_SL g2893 ( 
.A(n_2532),
.Y(n_2893)
);

INVx2_ASAP7_75t_SL g2894 ( 
.A(n_2534),
.Y(n_2894)
);

NAND2xp33_ASAP7_75t_L g2895 ( 
.A(n_2716),
.B(n_2499),
.Y(n_2895)
);

INVx5_ASAP7_75t_L g2896 ( 
.A(n_2711),
.Y(n_2896)
);

AOI21xp5_ASAP7_75t_L g2897 ( 
.A1(n_2646),
.A2(n_2689),
.B(n_2688),
.Y(n_2897)
);

OAI21x1_ASAP7_75t_L g2898 ( 
.A1(n_2749),
.A2(n_2443),
.B(n_2435),
.Y(n_2898)
);

OR2x2_ASAP7_75t_L g2899 ( 
.A(n_2637),
.B(n_2385),
.Y(n_2899)
);

OAI22xp5_ASAP7_75t_L g2900 ( 
.A1(n_2556),
.A2(n_2451),
.B1(n_2484),
.B2(n_2458),
.Y(n_2900)
);

CKINVDCx20_ASAP7_75t_R g2901 ( 
.A(n_2669),
.Y(n_2901)
);

OR2x2_ASAP7_75t_L g2902 ( 
.A(n_2675),
.B(n_2398),
.Y(n_2902)
);

CKINVDCx14_ASAP7_75t_R g2903 ( 
.A(n_2670),
.Y(n_2903)
);

OAI21x1_ASAP7_75t_L g2904 ( 
.A1(n_2682),
.A2(n_2448),
.B(n_2457),
.Y(n_2904)
);

AO21x2_ASAP7_75t_L g2905 ( 
.A1(n_2772),
.A2(n_16),
.B(n_17),
.Y(n_2905)
);

OR2x6_ASAP7_75t_L g2906 ( 
.A(n_2704),
.B(n_986),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2774),
.Y(n_2907)
);

AOI21x1_ASAP7_75t_L g2908 ( 
.A1(n_2655),
.A2(n_18),
.B(n_19),
.Y(n_2908)
);

NOR2xp67_ASAP7_75t_SL g2909 ( 
.A(n_2747),
.B(n_1033),
.Y(n_2909)
);

OAI21xp5_ASAP7_75t_L g2910 ( 
.A1(n_2692),
.A2(n_407),
.B(n_401),
.Y(n_2910)
);

OAI21x1_ASAP7_75t_L g2911 ( 
.A1(n_2682),
.A2(n_409),
.B(n_408),
.Y(n_2911)
);

OAI21x1_ASAP7_75t_L g2912 ( 
.A1(n_2622),
.A2(n_411),
.B(n_410),
.Y(n_2912)
);

OAI22xp5_ASAP7_75t_L g2913 ( 
.A1(n_2556),
.A2(n_978),
.B1(n_20),
.B2(n_18),
.Y(n_2913)
);

OAI21x1_ASAP7_75t_L g2914 ( 
.A1(n_2726),
.A2(n_414),
.B(n_412),
.Y(n_2914)
);

OAI21x1_ASAP7_75t_L g2915 ( 
.A1(n_2587),
.A2(n_417),
.B(n_415),
.Y(n_2915)
);

A2O1A1Ixp33_ASAP7_75t_L g2916 ( 
.A1(n_2570),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2539),
.Y(n_2917)
);

NAND2x1p5_ASAP7_75t_L g2918 ( 
.A(n_2547),
.B(n_1033),
.Y(n_2918)
);

BUFx2_ASAP7_75t_L g2919 ( 
.A(n_2713),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2545),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2555),
.Y(n_2921)
);

OAI21xp5_ASAP7_75t_L g2922 ( 
.A1(n_2731),
.A2(n_422),
.B(n_418),
.Y(n_2922)
);

AO21x2_ASAP7_75t_L g2923 ( 
.A1(n_2551),
.A2(n_21),
.B(n_23),
.Y(n_2923)
);

OAI21xp5_ASAP7_75t_L g2924 ( 
.A1(n_2570),
.A2(n_425),
.B(n_424),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2565),
.Y(n_2925)
);

A2O1A1Ixp33_ASAP7_75t_L g2926 ( 
.A1(n_2573),
.A2(n_28),
.B(n_24),
.C(n_25),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2595),
.Y(n_2927)
);

HB1xp67_ASAP7_75t_L g2928 ( 
.A(n_2711),
.Y(n_2928)
);

OAI21xp5_ASAP7_75t_L g2929 ( 
.A1(n_2573),
.A2(n_433),
.B(n_430),
.Y(n_2929)
);

OAI21xp5_ASAP7_75t_L g2930 ( 
.A1(n_2734),
.A2(n_2733),
.B(n_2674),
.Y(n_2930)
);

AOI21x1_ASAP7_75t_L g2931 ( 
.A1(n_2521),
.A2(n_24),
.B(n_28),
.Y(n_2931)
);

HB1xp67_ASAP7_75t_L g2932 ( 
.A(n_2711),
.Y(n_2932)
);

BUFx6f_ASAP7_75t_L g2933 ( 
.A(n_2534),
.Y(n_2933)
);

NOR2xp33_ASAP7_75t_L g2934 ( 
.A(n_2785),
.B(n_33),
.Y(n_2934)
);

AO21x2_ASAP7_75t_L g2935 ( 
.A1(n_2551),
.A2(n_33),
.B(n_34),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2724),
.B(n_34),
.Y(n_2936)
);

OAI21x1_ASAP7_75t_L g2937 ( 
.A1(n_2599),
.A2(n_436),
.B(n_434),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2615),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2635),
.Y(n_2939)
);

OAI21x1_ASAP7_75t_SL g2940 ( 
.A1(n_2567),
.A2(n_35),
.B(n_36),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2572),
.B(n_36),
.Y(n_2941)
);

OAI21x1_ASAP7_75t_L g2942 ( 
.A1(n_2601),
.A2(n_439),
.B(n_437),
.Y(n_2942)
);

OAI21x1_ASAP7_75t_SL g2943 ( 
.A1(n_2553),
.A2(n_37),
.B(n_38),
.Y(n_2943)
);

OAI21x1_ASAP7_75t_L g2944 ( 
.A1(n_2601),
.A2(n_2592),
.B(n_2753),
.Y(n_2944)
);

OAI21x1_ASAP7_75t_L g2945 ( 
.A1(n_2753),
.A2(n_443),
.B(n_440),
.Y(n_2945)
);

BUFx2_ASAP7_75t_L g2946 ( 
.A(n_2679),
.Y(n_2946)
);

INVx3_ASAP7_75t_L g2947 ( 
.A(n_2671),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2640),
.Y(n_2948)
);

OAI21x1_ASAP7_75t_L g2949 ( 
.A1(n_2738),
.A2(n_447),
.B(n_444),
.Y(n_2949)
);

OAI21x1_ASAP7_75t_L g2950 ( 
.A1(n_2738),
.A2(n_2698),
.B(n_2630),
.Y(n_2950)
);

INVx5_ASAP7_75t_SL g2951 ( 
.A(n_2643),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2641),
.Y(n_2952)
);

OAI21x1_ASAP7_75t_L g2953 ( 
.A1(n_2624),
.A2(n_449),
.B(n_448),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2765),
.Y(n_2954)
);

AOI22xp33_ASAP7_75t_SL g2955 ( 
.A1(n_2662),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_2955)
);

AO31x2_ASAP7_75t_L g2956 ( 
.A1(n_2779),
.A2(n_41),
.A3(n_39),
.B(n_40),
.Y(n_2956)
);

AOI21x1_ASAP7_75t_L g2957 ( 
.A1(n_2751),
.A2(n_42),
.B(n_43),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2537),
.B(n_42),
.Y(n_2958)
);

CKINVDCx8_ASAP7_75t_R g2959 ( 
.A(n_2524),
.Y(n_2959)
);

AO32x2_ASAP7_75t_L g2960 ( 
.A1(n_2709),
.A2(n_45),
.A3(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2525),
.Y(n_2961)
);

CKINVDCx5p33_ASAP7_75t_R g2962 ( 
.A(n_2520),
.Y(n_2962)
);

NOR2xp33_ASAP7_75t_L g2963 ( 
.A(n_2707),
.B(n_44),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2700),
.Y(n_2964)
);

OAI21x1_ASAP7_75t_SL g2965 ( 
.A1(n_2553),
.A2(n_45),
.B(n_46),
.Y(n_2965)
);

OAI21x1_ASAP7_75t_L g2966 ( 
.A1(n_2698),
.A2(n_460),
.B(n_453),
.Y(n_2966)
);

OAI22xp5_ASAP7_75t_L g2967 ( 
.A1(n_2526),
.A2(n_2590),
.B1(n_2734),
.B2(n_2776),
.Y(n_2967)
);

OAI21x1_ASAP7_75t_L g2968 ( 
.A1(n_2697),
.A2(n_464),
.B(n_462),
.Y(n_2968)
);

BUFx3_ASAP7_75t_L g2969 ( 
.A(n_2534),
.Y(n_2969)
);

OAI21x1_ASAP7_75t_L g2970 ( 
.A1(n_2697),
.A2(n_2720),
.B(n_2717),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2578),
.B(n_47),
.Y(n_2971)
);

AND2x4_ASAP7_75t_L g2972 ( 
.A(n_2606),
.B(n_467),
.Y(n_2972)
);

HB1xp67_ASAP7_75t_L g2973 ( 
.A(n_2552),
.Y(n_2973)
);

AOI22xp33_ASAP7_75t_L g2974 ( 
.A1(n_2662),
.A2(n_51),
.B1(n_48),
.B2(n_50),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2721),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2680),
.Y(n_2976)
);

NOR2xp67_ASAP7_75t_L g2977 ( 
.A(n_2672),
.B(n_48),
.Y(n_2977)
);

OAI21x1_ASAP7_75t_L g2978 ( 
.A1(n_2717),
.A2(n_469),
.B(n_468),
.Y(n_2978)
);

AOI221xp5_ASAP7_75t_L g2979 ( 
.A1(n_2779),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.C(n_53),
.Y(n_2979)
);

AOI22xp33_ASAP7_75t_SL g2980 ( 
.A1(n_2725),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2980)
);

AND2x4_ASAP7_75t_L g2981 ( 
.A(n_2603),
.B(n_471),
.Y(n_2981)
);

OAI21x1_ASAP7_75t_L g2982 ( 
.A1(n_2720),
.A2(n_483),
.B(n_478),
.Y(n_2982)
);

OAI21x1_ASAP7_75t_SL g2983 ( 
.A1(n_2727),
.A2(n_54),
.B(n_56),
.Y(n_2983)
);

O2A1O1Ixp5_ASAP7_75t_L g2984 ( 
.A1(n_2758),
.A2(n_59),
.B(n_56),
.C(n_58),
.Y(n_2984)
);

NOR2xp33_ASAP7_75t_L g2985 ( 
.A(n_2707),
.B(n_59),
.Y(n_2985)
);

AOI22xp33_ASAP7_75t_L g2986 ( 
.A1(n_2559),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2986)
);

OAI21xp5_ASAP7_75t_L g2987 ( 
.A1(n_2579),
.A2(n_485),
.B(n_61),
.Y(n_2987)
);

OAI21xp5_ASAP7_75t_L g2988 ( 
.A1(n_2763),
.A2(n_62),
.B(n_63),
.Y(n_2988)
);

OAI22xp5_ASAP7_75t_L g2989 ( 
.A1(n_2590),
.A2(n_978),
.B1(n_65),
.B2(n_63),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2568),
.B(n_64),
.Y(n_2990)
);

OAI21x1_ASAP7_75t_L g2991 ( 
.A1(n_2780),
.A2(n_1055),
.B(n_1033),
.Y(n_2991)
);

OAI21xp5_ASAP7_75t_L g2992 ( 
.A1(n_2750),
.A2(n_64),
.B(n_65),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2540),
.Y(n_2993)
);

AND2x4_ASAP7_75t_L g2994 ( 
.A(n_2603),
.B(n_67),
.Y(n_2994)
);

AOI22xp5_ASAP7_75t_L g2995 ( 
.A1(n_2770),
.A2(n_2571),
.B1(n_2775),
.B2(n_2559),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2569),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2552),
.Y(n_2997)
);

OA21x2_ASAP7_75t_L g2998 ( 
.A1(n_2696),
.A2(n_2757),
.B(n_2732),
.Y(n_2998)
);

OR2x6_ASAP7_75t_L g2999 ( 
.A(n_2643),
.B(n_1055),
.Y(n_2999)
);

INVx8_ASAP7_75t_L g3000 ( 
.A(n_2643),
.Y(n_3000)
);

AOI221xp5_ASAP7_75t_L g3001 ( 
.A1(n_2722),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.C(n_71),
.Y(n_3001)
);

NAND2x1p5_ASAP7_75t_L g3002 ( 
.A(n_2547),
.B(n_1055),
.Y(n_3002)
);

OAI21x1_ASAP7_75t_L g3003 ( 
.A1(n_2672),
.A2(n_1059),
.B(n_1009),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2598),
.Y(n_3004)
);

AO21x2_ASAP7_75t_L g3005 ( 
.A1(n_2744),
.A2(n_68),
.B(n_69),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2569),
.Y(n_3006)
);

AND2x4_ASAP7_75t_L g3007 ( 
.A(n_2519),
.B(n_70),
.Y(n_3007)
);

BUFx2_ASAP7_75t_L g3008 ( 
.A(n_2618),
.Y(n_3008)
);

HB1xp67_ASAP7_75t_L g3009 ( 
.A(n_2598),
.Y(n_3009)
);

INVx3_ASAP7_75t_L g3010 ( 
.A(n_2739),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2569),
.Y(n_3011)
);

CKINVDCx9p33_ASAP7_75t_R g3012 ( 
.A(n_2610),
.Y(n_3012)
);

OAI21x1_ASAP7_75t_L g3013 ( 
.A1(n_2571),
.A2(n_1059),
.B(n_1009),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2602),
.Y(n_3014)
);

OAI21x1_ASAP7_75t_L g3015 ( 
.A1(n_2586),
.A2(n_1059),
.B(n_1009),
.Y(n_3015)
);

BUFx2_ASAP7_75t_L g3016 ( 
.A(n_2618),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_2786),
.Y(n_3017)
);

AOI22xp33_ASAP7_75t_L g3018 ( 
.A1(n_2816),
.A2(n_2690),
.B1(n_2732),
.B2(n_2725),
.Y(n_3018)
);

OR2x2_ASAP7_75t_L g3019 ( 
.A(n_2864),
.B(n_2673),
.Y(n_3019)
);

INVx1_ASAP7_75t_SL g3020 ( 
.A(n_2885),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2816),
.A2(n_2705),
.B(n_2547),
.Y(n_3021)
);

BUFx3_ASAP7_75t_L g3022 ( 
.A(n_2842),
.Y(n_3022)
);

BUFx12f_ASAP7_75t_L g3023 ( 
.A(n_2891),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_SL g3024 ( 
.A(n_2812),
.B(n_2707),
.Y(n_3024)
);

AOI221xp5_ASAP7_75t_L g3025 ( 
.A1(n_2979),
.A2(n_2745),
.B1(n_2722),
.B2(n_2702),
.C(n_2684),
.Y(n_3025)
);

AOI22xp33_ASAP7_75t_L g3026 ( 
.A1(n_2930),
.A2(n_2691),
.B1(n_2745),
.B2(n_2681),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2786),
.Y(n_3027)
);

BUFx2_ASAP7_75t_L g3028 ( 
.A(n_2946),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2787),
.Y(n_3029)
);

AO21x2_ASAP7_75t_L g3030 ( 
.A1(n_2826),
.A2(n_2666),
.B(n_2647),
.Y(n_3030)
);

OAI21xp5_ASAP7_75t_L g3031 ( 
.A1(n_2987),
.A2(n_2677),
.B(n_2684),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2787),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2789),
.Y(n_3033)
);

INVx1_ASAP7_75t_SL g3034 ( 
.A(n_2919),
.Y(n_3034)
);

INVx5_ASAP7_75t_SL g3035 ( 
.A(n_3012),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2872),
.B(n_2542),
.Y(n_3036)
);

AOI22xp33_ASAP7_75t_SL g3037 ( 
.A1(n_2967),
.A2(n_2759),
.B1(n_2638),
.B2(n_2771),
.Y(n_3037)
);

CKINVDCx20_ASAP7_75t_R g3038 ( 
.A(n_2797),
.Y(n_3038)
);

AND2x4_ASAP7_75t_L g3039 ( 
.A(n_2867),
.B(n_2524),
.Y(n_3039)
);

AOI22xp33_ASAP7_75t_L g3040 ( 
.A1(n_2924),
.A2(n_2929),
.B1(n_2812),
.B2(n_2910),
.Y(n_3040)
);

OR2x2_ASAP7_75t_L g3041 ( 
.A(n_2815),
.B(n_2696),
.Y(n_3041)
);

AOI22xp33_ASAP7_75t_L g3042 ( 
.A1(n_2859),
.A2(n_2740),
.B1(n_2741),
.B2(n_2718),
.Y(n_3042)
);

INVx4_ASAP7_75t_L g3043 ( 
.A(n_2860),
.Y(n_3043)
);

INVx3_ASAP7_75t_L g3044 ( 
.A(n_3010),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2789),
.Y(n_3045)
);

BUFx6f_ASAP7_75t_L g3046 ( 
.A(n_2959),
.Y(n_3046)
);

AND2x2_ASAP7_75t_L g3047 ( 
.A(n_2875),
.B(n_2618),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2792),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2792),
.Y(n_3049)
);

OAI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_2859),
.A2(n_2528),
.B1(n_2638),
.B2(n_2705),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2806),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2973),
.B(n_2623),
.Y(n_3052)
);

CKINVDCx6p67_ASAP7_75t_R g3053 ( 
.A(n_2797),
.Y(n_3053)
);

AOI22xp33_ASAP7_75t_L g3054 ( 
.A1(n_3001),
.A2(n_2742),
.B1(n_2695),
.B2(n_2706),
.Y(n_3054)
);

OR2x6_ASAP7_75t_L g3055 ( 
.A(n_3000),
.B(n_2728),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_3014),
.B(n_2549),
.Y(n_3056)
);

BUFx6f_ASAP7_75t_L g3057 ( 
.A(n_2817),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2973),
.B(n_3009),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_3009),
.B(n_2623),
.Y(n_3059)
);

OAI22xp5_ASAP7_75t_SL g3060 ( 
.A1(n_2901),
.A2(n_2611),
.B1(n_2574),
.B2(n_2625),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2829),
.B(n_2687),
.Y(n_3061)
);

NAND2xp33_ASAP7_75t_R g3062 ( 
.A(n_2891),
.B(n_2548),
.Y(n_3062)
);

AOI22xp33_ASAP7_75t_L g3063 ( 
.A1(n_2986),
.A2(n_2710),
.B1(n_2677),
.B2(n_2548),
.Y(n_3063)
);

AOI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_2834),
.A2(n_2759),
.B1(n_2519),
.B2(n_2633),
.Y(n_3064)
);

NAND3xp33_ASAP7_75t_L g3065 ( 
.A(n_2916),
.B(n_2926),
.C(n_2974),
.Y(n_3065)
);

BUFx4f_ASAP7_75t_SL g3066 ( 
.A(n_2842),
.Y(n_3066)
);

INVx3_ASAP7_75t_L g3067 ( 
.A(n_3010),
.Y(n_3067)
);

BUFx4f_ASAP7_75t_SL g3068 ( 
.A(n_2901),
.Y(n_3068)
);

OAI22xp33_ASAP7_75t_L g3069 ( 
.A1(n_2992),
.A2(n_2705),
.B1(n_2616),
.B2(n_2728),
.Y(n_3069)
);

AOI22xp33_ASAP7_75t_L g3070 ( 
.A1(n_2813),
.A2(n_2747),
.B1(n_2777),
.B2(n_2687),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2806),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2837),
.B(n_2687),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2821),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2821),
.Y(n_3074)
);

INVx1_ASAP7_75t_SL g3075 ( 
.A(n_2874),
.Y(n_3075)
);

AOI22xp33_ASAP7_75t_SL g3076 ( 
.A1(n_2934),
.A2(n_2569),
.B1(n_2736),
.B2(n_2728),
.Y(n_3076)
);

OAI22xp5_ASAP7_75t_L g3077 ( 
.A1(n_2986),
.A2(n_2710),
.B1(n_2736),
.B2(n_2541),
.Y(n_3077)
);

AOI22xp33_ASAP7_75t_L g3078 ( 
.A1(n_2974),
.A2(n_2747),
.B1(n_2651),
.B2(n_2658),
.Y(n_3078)
);

AOI22xp33_ASAP7_75t_L g3079 ( 
.A1(n_2955),
.A2(n_2651),
.B1(n_2658),
.B2(n_2652),
.Y(n_3079)
);

AOI22xp5_ASAP7_75t_L g3080 ( 
.A1(n_2989),
.A2(n_2541),
.B1(n_2664),
.B2(n_2632),
.Y(n_3080)
);

AND2x2_ASAP7_75t_L g3081 ( 
.A(n_2884),
.B(n_2557),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2788),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2796),
.Y(n_3083)
);

BUFx2_ASAP7_75t_L g3084 ( 
.A(n_3008),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2802),
.Y(n_3085)
);

AOI22xp33_ASAP7_75t_L g3086 ( 
.A1(n_2913),
.A2(n_2652),
.B1(n_2612),
.B2(n_2664),
.Y(n_3086)
);

INVx4_ASAP7_75t_SL g3087 ( 
.A(n_2956),
.Y(n_3087)
);

AOI22xp33_ASAP7_75t_L g3088 ( 
.A1(n_2793),
.A2(n_2663),
.B1(n_2687),
.B2(n_2645),
.Y(n_3088)
);

BUFx6f_ASAP7_75t_L g3089 ( 
.A(n_2817),
.Y(n_3089)
);

OR2x2_ASAP7_75t_L g3090 ( 
.A(n_2825),
.B(n_2729),
.Y(n_3090)
);

OAI22xp33_ASAP7_75t_L g3091 ( 
.A1(n_2995),
.A2(n_2736),
.B1(n_2727),
.B2(n_2657),
.Y(n_3091)
);

AOI22xp33_ASAP7_75t_SL g3092 ( 
.A1(n_2934),
.A2(n_2569),
.B1(n_2531),
.B2(n_2632),
.Y(n_3092)
);

OAI22xp5_ASAP7_75t_L g3093 ( 
.A1(n_2916),
.A2(n_2645),
.B1(n_2561),
.B2(n_2586),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2863),
.B(n_2657),
.Y(n_3094)
);

BUFx3_ASAP7_75t_L g3095 ( 
.A(n_2962),
.Y(n_3095)
);

BUFx6f_ASAP7_75t_L g3096 ( 
.A(n_2817),
.Y(n_3096)
);

AND2x2_ASAP7_75t_L g3097 ( 
.A(n_2819),
.B(n_3016),
.Y(n_3097)
);

AOI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_2843),
.A2(n_2617),
.B1(n_2614),
.B2(n_2531),
.Y(n_3098)
);

AOI22xp33_ASAP7_75t_L g3099 ( 
.A1(n_2793),
.A2(n_2644),
.B1(n_2665),
.B2(n_2660),
.Y(n_3099)
);

OAI22xp33_ASAP7_75t_L g3100 ( 
.A1(n_2988),
.A2(n_2686),
.B1(n_2660),
.B2(n_2665),
.Y(n_3100)
);

AND2x2_ASAP7_75t_L g3101 ( 
.A(n_2880),
.B(n_2644),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_2997),
.B(n_2644),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_3004),
.B(n_2883),
.Y(n_3103)
);

INVx3_ASAP7_75t_L g3104 ( 
.A(n_2800),
.Y(n_3104)
);

OAI21x1_ASAP7_75t_L g3105 ( 
.A1(n_2804),
.A2(n_2650),
.B(n_2729),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2883),
.B(n_2659),
.Y(n_3106)
);

OR2x2_ASAP7_75t_L g3107 ( 
.A(n_2820),
.B(n_2729),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2807),
.Y(n_3108)
);

AOI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_2922),
.A2(n_2620),
.B1(n_2665),
.B2(n_2660),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2827),
.B(n_2620),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_2976),
.B(n_2964),
.Y(n_3111)
);

OAI211xp5_ASAP7_75t_SL g3112 ( 
.A1(n_2926),
.A2(n_2639),
.B(n_2650),
.C(n_2656),
.Y(n_3112)
);

AOI22xp5_ASAP7_75t_L g3113 ( 
.A1(n_2843),
.A2(n_2614),
.B1(n_2617),
.B2(n_2620),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_2809),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2954),
.B(n_2712),
.Y(n_3115)
);

CKINVDCx5p33_ASAP7_75t_R g3116 ( 
.A(n_2848),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2838),
.Y(n_3117)
);

AO31x2_ASAP7_75t_L g3118 ( 
.A1(n_2897),
.A2(n_2588),
.A3(n_2686),
.B(n_2712),
.Y(n_3118)
);

BUFx2_ASAP7_75t_L g3119 ( 
.A(n_3012),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2917),
.Y(n_3120)
);

OAI22xp5_ASAP7_75t_L g3121 ( 
.A1(n_2980),
.A2(n_2686),
.B1(n_2591),
.B2(n_2607),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_2917),
.Y(n_3122)
);

BUFx3_ASAP7_75t_L g3123 ( 
.A(n_2962),
.Y(n_3123)
);

AOI22xp5_ASAP7_75t_L g3124 ( 
.A1(n_2828),
.A2(n_2588),
.B1(n_2591),
.B2(n_2583),
.Y(n_3124)
);

OAI21xp33_ASAP7_75t_L g3125 ( 
.A1(n_2828),
.A2(n_2712),
.B(n_2591),
.Y(n_3125)
);

INVx3_ASAP7_75t_L g3126 ( 
.A(n_2800),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2858),
.Y(n_3127)
);

AOI221xp5_ASAP7_75t_L g3128 ( 
.A1(n_2940),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.C(n_75),
.Y(n_3128)
);

CKINVDCx5p33_ASAP7_75t_R g3129 ( 
.A(n_2848),
.Y(n_3129)
);

AOI221xp5_ASAP7_75t_L g3130 ( 
.A1(n_2790),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.C(n_76),
.Y(n_3130)
);

NAND3xp33_ASAP7_75t_L g3131 ( 
.A(n_2818),
.B(n_2607),
.C(n_2583),
.Y(n_3131)
);

INVx4_ASAP7_75t_L g3132 ( 
.A(n_3000),
.Y(n_3132)
);

AOI221xp5_ASAP7_75t_L g3133 ( 
.A1(n_2984),
.A2(n_79),
.B1(n_76),
.B2(n_77),
.C(n_80),
.Y(n_3133)
);

AOI221xp5_ASAP7_75t_L g3134 ( 
.A1(n_2943),
.A2(n_84),
.B1(n_77),
.B2(n_83),
.C(n_85),
.Y(n_3134)
);

AOI221xp5_ASAP7_75t_L g3135 ( 
.A1(n_2965),
.A2(n_2975),
.B1(n_2936),
.B2(n_3005),
.C(n_2985),
.Y(n_3135)
);

OAI22xp5_ASAP7_75t_L g3136 ( 
.A1(n_2903),
.A2(n_2607),
.B1(n_2588),
.B2(n_87),
.Y(n_3136)
);

NAND3xp33_ASAP7_75t_SL g3137 ( 
.A(n_2963),
.B(n_2588),
.C(n_83),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2993),
.B(n_86),
.Y(n_3138)
);

AOI21xp5_ASAP7_75t_L g3139 ( 
.A1(n_2895),
.A2(n_2799),
.B(n_2945),
.Y(n_3139)
);

OAI22xp5_ASAP7_75t_L g3140 ( 
.A1(n_2903),
.A2(n_89),
.B1(n_86),
.B2(n_88),
.Y(n_3140)
);

OR2x2_ASAP7_75t_L g3141 ( 
.A(n_2824),
.B(n_88),
.Y(n_3141)
);

OAI21x1_ASAP7_75t_L g3142 ( 
.A1(n_2811),
.A2(n_91),
.B(n_92),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2938),
.Y(n_3143)
);

AOI21xp5_ASAP7_75t_L g3144 ( 
.A1(n_2895),
.A2(n_1119),
.B(n_1117),
.Y(n_3144)
);

INVxp67_ASAP7_75t_L g3145 ( 
.A(n_2865),
.Y(n_3145)
);

OAI21x1_ASAP7_75t_L g3146 ( 
.A1(n_2811),
.A2(n_93),
.B(n_94),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2938),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2853),
.Y(n_3148)
);

OAI221xp5_ASAP7_75t_L g3149 ( 
.A1(n_2963),
.A2(n_96),
.B1(n_93),
.B2(n_95),
.C(n_97),
.Y(n_3149)
);

OR2x6_ASAP7_75t_L g3150 ( 
.A(n_3000),
.B(n_1059),
.Y(n_3150)
);

HB1xp67_ASAP7_75t_L g3151 ( 
.A(n_2826),
.Y(n_3151)
);

AOI221xp5_ASAP7_75t_L g3152 ( 
.A1(n_3005),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.C(n_101),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2855),
.B(n_99),
.Y(n_3153)
);

NAND3xp33_ASAP7_75t_SL g3154 ( 
.A(n_2985),
.B(n_100),
.C(n_102),
.Y(n_3154)
);

AND2x4_ASAP7_75t_L g3155 ( 
.A(n_2867),
.B(n_103),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2948),
.Y(n_3156)
);

NAND2xp33_ASAP7_75t_R g3157 ( 
.A(n_2830),
.B(n_104),
.Y(n_3157)
);

AO21x2_ASAP7_75t_L g3158 ( 
.A1(n_2805),
.A2(n_105),
.B(n_108),
.Y(n_3158)
);

INVx3_ASAP7_75t_L g3159 ( 
.A(n_2852),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2948),
.Y(n_3160)
);

CKINVDCx5p33_ASAP7_75t_R g3161 ( 
.A(n_2822),
.Y(n_3161)
);

CKINVDCx5p33_ASAP7_75t_R g3162 ( 
.A(n_2874),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2855),
.B(n_105),
.Y(n_3163)
);

HB1xp67_ASAP7_75t_L g3164 ( 
.A(n_2856),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2879),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_2892),
.B(n_108),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2952),
.Y(n_3167)
);

O2A1O1Ixp33_ASAP7_75t_L g3168 ( 
.A1(n_2983),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_2952),
.Y(n_3169)
);

AOI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_2799),
.A2(n_1119),
.B(n_1117),
.Y(n_3170)
);

NOR2x1p5_ASAP7_75t_L g3171 ( 
.A(n_2931),
.B(n_1059),
.Y(n_3171)
);

OAI22xp33_ASAP7_75t_L g3172 ( 
.A1(n_2957),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_3172)
);

INVx3_ASAP7_75t_L g3173 ( 
.A(n_2852),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2879),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2889),
.Y(n_3175)
);

AND2x2_ASAP7_75t_L g3176 ( 
.A(n_2867),
.B(n_113),
.Y(n_3176)
);

OAI22xp5_ASAP7_75t_L g3177 ( 
.A1(n_2876),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2877),
.B(n_114),
.Y(n_3178)
);

AOI22xp33_ASAP7_75t_L g3179 ( 
.A1(n_2905),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2889),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_2996),
.B(n_116),
.Y(n_3181)
);

BUFx12f_ASAP7_75t_L g3182 ( 
.A(n_2990),
.Y(n_3182)
);

AOI22xp33_ASAP7_75t_L g3183 ( 
.A1(n_2905),
.A2(n_120),
.B1(n_117),
.B2(n_119),
.Y(n_3183)
);

INVx2_ASAP7_75t_SL g3184 ( 
.A(n_2794),
.Y(n_3184)
);

OAI22xp5_ASAP7_75t_L g3185 ( 
.A1(n_2999),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_3185)
);

INVx4_ASAP7_75t_L g3186 ( 
.A(n_2817),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2907),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2920),
.B(n_122),
.Y(n_3188)
);

AOI22xp33_ASAP7_75t_L g3189 ( 
.A1(n_2803),
.A2(n_1062),
.B1(n_1070),
.B2(n_1009),
.Y(n_3189)
);

AOI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_2945),
.A2(n_1122),
.B(n_1119),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_2971),
.B(n_123),
.Y(n_3191)
);

INVx2_ASAP7_75t_SL g3192 ( 
.A(n_2794),
.Y(n_3192)
);

AND2x2_ASAP7_75t_SL g3193 ( 
.A(n_2972),
.B(n_123),
.Y(n_3193)
);

OAI22xp33_ASAP7_75t_L g3194 ( 
.A1(n_2999),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_3194)
);

INVx1_ASAP7_75t_SL g3195 ( 
.A(n_2798),
.Y(n_3195)
);

CKINVDCx11_ASAP7_75t_R g3196 ( 
.A(n_2866),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2921),
.Y(n_3197)
);

NOR2x1_ASAP7_75t_SL g3198 ( 
.A(n_2831),
.B(n_124),
.Y(n_3198)
);

NAND2xp33_ASAP7_75t_SL g3199 ( 
.A(n_3007),
.B(n_125),
.Y(n_3199)
);

AOI221xp5_ASAP7_75t_L g3200 ( 
.A1(n_2941),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.C(n_129),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2925),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_2996),
.B(n_127),
.Y(n_3202)
);

CKINVDCx20_ASAP7_75t_R g3203 ( 
.A(n_2798),
.Y(n_3203)
);

BUFx4f_ASAP7_75t_L g3204 ( 
.A(n_2981),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2927),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2939),
.B(n_128),
.Y(n_3206)
);

OAI21x1_ASAP7_75t_L g3207 ( 
.A1(n_2851),
.A2(n_130),
.B(n_131),
.Y(n_3207)
);

OAI222xp33_ASAP7_75t_L g3208 ( 
.A1(n_2999),
.A2(n_2845),
.B1(n_2994),
.B2(n_2831),
.C1(n_2839),
.C2(n_2890),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_2961),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2902),
.Y(n_3210)
);

AOI22xp33_ASAP7_75t_SL g3211 ( 
.A1(n_2998),
.A2(n_2935),
.B1(n_2923),
.B2(n_2994),
.Y(n_3211)
);

AND2x4_ASAP7_75t_L g3212 ( 
.A(n_3006),
.B(n_130),
.Y(n_3212)
);

INVxp67_ASAP7_75t_L g3213 ( 
.A(n_2899),
.Y(n_3213)
);

AOI22xp33_ASAP7_75t_SL g3214 ( 
.A1(n_2998),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_3214)
);

AND2x4_ASAP7_75t_L g3215 ( 
.A(n_3006),
.B(n_132),
.Y(n_3215)
);

AND2x2_ASAP7_75t_L g3216 ( 
.A(n_3011),
.B(n_133),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_2950),
.Y(n_3217)
);

AOI22xp33_ASAP7_75t_SL g3218 ( 
.A1(n_2998),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_3218)
);

HB1xp67_ASAP7_75t_L g3219 ( 
.A(n_3213),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3127),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_3058),
.B(n_2850),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_3027),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3032),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3033),
.Y(n_3224)
);

OR2x2_ASAP7_75t_L g3225 ( 
.A(n_3213),
.B(n_2854),
.Y(n_3225)
);

OR2x2_ASAP7_75t_L g3226 ( 
.A(n_3210),
.B(n_2814),
.Y(n_3226)
);

INVx2_ASAP7_75t_SL g3227 ( 
.A(n_3039),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3045),
.Y(n_3228)
);

OA21x2_ASAP7_75t_L g3229 ( 
.A1(n_3151),
.A2(n_2836),
.B(n_2844),
.Y(n_3229)
);

INVxp67_ASAP7_75t_SL g3230 ( 
.A(n_3164),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_3103),
.B(n_2850),
.Y(n_3231)
);

OAI21x1_ASAP7_75t_L g3232 ( 
.A1(n_3170),
.A2(n_2836),
.B(n_2846),
.Y(n_3232)
);

BUFx3_ASAP7_75t_L g3233 ( 
.A(n_3023),
.Y(n_3233)
);

AO21x2_ASAP7_75t_L g3234 ( 
.A1(n_3151),
.A2(n_2844),
.B(n_2805),
.Y(n_3234)
);

BUFx3_ASAP7_75t_L g3235 ( 
.A(n_3068),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_3048),
.Y(n_3236)
);

OR2x6_ASAP7_75t_L g3237 ( 
.A(n_3144),
.B(n_2831),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_3049),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_3071),
.Y(n_3239)
);

OAI21x1_ASAP7_75t_L g3240 ( 
.A1(n_3170),
.A2(n_2846),
.B(n_2857),
.Y(n_3240)
);

INVx2_ASAP7_75t_SL g3241 ( 
.A(n_3039),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3074),
.Y(n_3242)
);

OA21x2_ASAP7_75t_L g3243 ( 
.A1(n_3139),
.A2(n_2823),
.B(n_2851),
.Y(n_3243)
);

OAI21x1_ASAP7_75t_L g3244 ( 
.A1(n_3139),
.A2(n_2857),
.B(n_2795),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3017),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3029),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_3051),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_3030),
.B(n_2840),
.Y(n_3248)
);

AND2x2_ASAP7_75t_L g3249 ( 
.A(n_3084),
.B(n_2840),
.Y(n_3249)
);

AND2x2_ASAP7_75t_L g3250 ( 
.A(n_3028),
.B(n_2840),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3073),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_3082),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3108),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_3120),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_3097),
.B(n_3047),
.Y(n_3255)
);

NAND2x1p5_ASAP7_75t_L g3256 ( 
.A(n_3144),
.B(n_2896),
.Y(n_3256)
);

INVx3_ASAP7_75t_L g3257 ( 
.A(n_3186),
.Y(n_3257)
);

AND2x4_ASAP7_75t_L g3258 ( 
.A(n_3087),
.B(n_3011),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_3122),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3083),
.Y(n_3260)
);

AO21x2_ASAP7_75t_L g3261 ( 
.A1(n_3158),
.A2(n_3190),
.B(n_3030),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3085),
.Y(n_3262)
);

BUFx3_ASAP7_75t_L g3263 ( 
.A(n_3068),
.Y(n_3263)
);

AO222x2_ASAP7_75t_L g3264 ( 
.A1(n_3157),
.A2(n_2958),
.B1(n_2994),
.B2(n_3007),
.C1(n_138),
.C2(n_139),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_3110),
.B(n_2861),
.Y(n_3265)
);

HB1xp67_ASAP7_75t_L g3266 ( 
.A(n_3164),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_3143),
.Y(n_3267)
);

OAI21x1_ASAP7_75t_L g3268 ( 
.A1(n_3105),
.A2(n_2795),
.B(n_2823),
.Y(n_3268)
);

INVx2_ASAP7_75t_SL g3269 ( 
.A(n_3044),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_3147),
.Y(n_3270)
);

AOI221xp5_ASAP7_75t_L g3271 ( 
.A1(n_3154),
.A2(n_3007),
.B1(n_2882),
.B2(n_2923),
.C(n_2935),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_3156),
.Y(n_3272)
);

OAI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_3040),
.A2(n_2977),
.B(n_2878),
.Y(n_3273)
);

NAND2x1p5_ASAP7_75t_L g3274 ( 
.A(n_3021),
.B(n_2896),
.Y(n_3274)
);

BUFx2_ASAP7_75t_L g3275 ( 
.A(n_3119),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_3052),
.B(n_2861),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_3160),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3114),
.Y(n_3278)
);

HB1xp67_ASAP7_75t_L g3279 ( 
.A(n_3145),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3165),
.Y(n_3280)
);

OR2x2_ASAP7_75t_L g3281 ( 
.A(n_3107),
.B(n_2814),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3175),
.Y(n_3282)
);

INVx2_ASAP7_75t_SL g3283 ( 
.A(n_3044),
.Y(n_3283)
);

AOI21xp5_ASAP7_75t_L g3284 ( 
.A1(n_3031),
.A2(n_2900),
.B(n_2839),
.Y(n_3284)
);

INVx2_ASAP7_75t_SL g3285 ( 
.A(n_3067),
.Y(n_3285)
);

OAI21x1_ASAP7_75t_L g3286 ( 
.A1(n_3190),
.A2(n_2808),
.B(n_2810),
.Y(n_3286)
);

BUFx6f_ASAP7_75t_L g3287 ( 
.A(n_3046),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3180),
.Y(n_3288)
);

OR2x6_ASAP7_75t_L g3289 ( 
.A(n_3021),
.B(n_2839),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3167),
.Y(n_3290)
);

AND2x2_ASAP7_75t_L g3291 ( 
.A(n_3059),
.B(n_2862),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3145),
.Y(n_3292)
);

INVx2_ASAP7_75t_L g3293 ( 
.A(n_3169),
.Y(n_3293)
);

INVx2_ASAP7_75t_SL g3294 ( 
.A(n_3067),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_3111),
.B(n_2862),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3174),
.Y(n_3296)
);

HB1xp67_ASAP7_75t_L g3297 ( 
.A(n_3041),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3117),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3197),
.Y(n_3299)
);

INVx3_ASAP7_75t_L g3300 ( 
.A(n_3186),
.Y(n_3300)
);

INVx2_ASAP7_75t_L g3301 ( 
.A(n_3217),
.Y(n_3301)
);

AO21x1_ASAP7_75t_SL g3302 ( 
.A1(n_3208),
.A2(n_2932),
.B(n_2928),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3201),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3205),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3187),
.Y(n_3305)
);

OAI21x1_ASAP7_75t_L g3306 ( 
.A1(n_3142),
.A2(n_2808),
.B(n_2810),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3148),
.Y(n_3307)
);

BUFx3_ASAP7_75t_L g3308 ( 
.A(n_3053),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3209),
.Y(n_3309)
);

INVx3_ASAP7_75t_L g3310 ( 
.A(n_3104),
.Y(n_3310)
);

OAI21x1_ASAP7_75t_L g3311 ( 
.A1(n_3146),
.A2(n_2881),
.B(n_2904),
.Y(n_3311)
);

NAND3xp33_ASAP7_75t_L g3312 ( 
.A(n_3130),
.B(n_2887),
.C(n_2928),
.Y(n_3312)
);

OA21x2_ASAP7_75t_L g3313 ( 
.A1(n_3207),
.A2(n_2904),
.B(n_2911),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3087),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3087),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3090),
.Y(n_3316)
);

CKINVDCx8_ASAP7_75t_R g3317 ( 
.A(n_3046),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_3019),
.B(n_2870),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_3094),
.Y(n_3319)
);

HB1xp67_ASAP7_75t_L g3320 ( 
.A(n_3104),
.Y(n_3320)
);

BUFx6f_ASAP7_75t_L g3321 ( 
.A(n_3046),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3126),
.Y(n_3322)
);

INVx3_ASAP7_75t_L g3323 ( 
.A(n_3126),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_3159),
.Y(n_3324)
);

AO21x2_ASAP7_75t_L g3325 ( 
.A1(n_3158),
.A2(n_2870),
.B(n_2898),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_3106),
.B(n_2932),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3159),
.Y(n_3327)
);

INVx2_ASAP7_75t_SL g3328 ( 
.A(n_3173),
.Y(n_3328)
);

AO21x1_ASAP7_75t_L g3329 ( 
.A1(n_3172),
.A2(n_2960),
.B(n_2972),
.Y(n_3329)
);

BUFx3_ASAP7_75t_L g3330 ( 
.A(n_3066),
.Y(n_3330)
);

HB1xp67_ASAP7_75t_L g3331 ( 
.A(n_3173),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_3102),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_3101),
.B(n_2896),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_3141),
.B(n_2947),
.Y(n_3334)
);

BUFx2_ASAP7_75t_L g3335 ( 
.A(n_3118),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_3081),
.Y(n_3336)
);

AND2x2_ASAP7_75t_L g3337 ( 
.A(n_3195),
.B(n_2896),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_3115),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_3181),
.Y(n_3339)
);

AO21x2_ASAP7_75t_L g3340 ( 
.A1(n_3131),
.A2(n_3172),
.B(n_3208),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3061),
.Y(n_3341)
);

OAI21xp5_ASAP7_75t_L g3342 ( 
.A1(n_3065),
.A2(n_2970),
.B(n_2937),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_3202),
.Y(n_3343)
);

OR2x2_ASAP7_75t_L g3344 ( 
.A(n_3072),
.B(n_2868),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3188),
.Y(n_3345)
);

AND2x4_ASAP7_75t_L g3346 ( 
.A(n_3118),
.B(n_2970),
.Y(n_3346)
);

HB1xp67_ASAP7_75t_L g3347 ( 
.A(n_3118),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_3035),
.B(n_2847),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_3216),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3206),
.Y(n_3350)
);

AOI22xp33_ASAP7_75t_SL g3351 ( 
.A1(n_3193),
.A2(n_2951),
.B1(n_2981),
.B2(n_2972),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3118),
.Y(n_3352)
);

INVx2_ASAP7_75t_SL g3353 ( 
.A(n_3184),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3211),
.Y(n_3354)
);

AND2x2_ASAP7_75t_L g3355 ( 
.A(n_3035),
.B(n_2847),
.Y(n_3355)
);

AO21x2_ASAP7_75t_L g3356 ( 
.A1(n_3125),
.A2(n_2898),
.B(n_2835),
.Y(n_3356)
);

AND2x2_ASAP7_75t_L g3357 ( 
.A(n_3035),
.B(n_3192),
.Y(n_3357)
);

HB1xp67_ASAP7_75t_L g3358 ( 
.A(n_3036),
.Y(n_3358)
);

CKINVDCx5p33_ASAP7_75t_R g3359 ( 
.A(n_3038),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_SL g3360 ( 
.A(n_3132),
.B(n_2947),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3056),
.B(n_3024),
.Y(n_3361)
);

INVx3_ASAP7_75t_L g3362 ( 
.A(n_3132),
.Y(n_3362)
);

HB1xp67_ASAP7_75t_L g3363 ( 
.A(n_3057),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3153),
.B(n_2849),
.Y(n_3364)
);

OAI21x1_ASAP7_75t_L g3365 ( 
.A1(n_3070),
.A2(n_2869),
.B(n_2801),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3020),
.B(n_2849),
.Y(n_3366)
);

OR2x6_ASAP7_75t_L g3367 ( 
.A(n_3055),
.B(n_2845),
.Y(n_3367)
);

BUFx2_ASAP7_75t_L g3368 ( 
.A(n_3203),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3211),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3163),
.B(n_2868),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3212),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3212),
.Y(n_3372)
);

HB1xp67_ASAP7_75t_L g3373 ( 
.A(n_3057),
.Y(n_3373)
);

OR2x2_ASAP7_75t_L g3374 ( 
.A(n_3034),
.B(n_2956),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3215),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3215),
.Y(n_3376)
);

OA21x2_ASAP7_75t_L g3377 ( 
.A1(n_3135),
.A2(n_2911),
.B(n_2944),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3057),
.Y(n_3378)
);

OAI21xp5_ASAP7_75t_L g3379 ( 
.A1(n_3037),
.A2(n_2937),
.B(n_2915),
.Y(n_3379)
);

OAI221xp5_ASAP7_75t_L g3380 ( 
.A1(n_3354),
.A2(n_3037),
.B1(n_3130),
.B2(n_3026),
.C(n_3042),
.Y(n_3380)
);

OAI22xp33_ASAP7_75t_L g3381 ( 
.A1(n_3312),
.A2(n_3137),
.B1(n_3177),
.B2(n_3064),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_3310),
.Y(n_3382)
);

OA21x2_ASAP7_75t_L g3383 ( 
.A1(n_3354),
.A2(n_3369),
.B(n_3231),
.Y(n_3383)
);

HB1xp67_ASAP7_75t_L g3384 ( 
.A(n_3266),
.Y(n_3384)
);

AOI22xp33_ASAP7_75t_L g3385 ( 
.A1(n_3329),
.A2(n_3025),
.B1(n_3154),
.B2(n_3149),
.Y(n_3385)
);

AOI22xp33_ASAP7_75t_L g3386 ( 
.A1(n_3329),
.A2(n_3025),
.B1(n_3200),
.B2(n_3042),
.Y(n_3386)
);

AND2x2_ASAP7_75t_L g3387 ( 
.A(n_3249),
.B(n_3043),
.Y(n_3387)
);

OR2x2_ASAP7_75t_L g3388 ( 
.A(n_3364),
.B(n_3178),
.Y(n_3388)
);

AND2x4_ASAP7_75t_L g3389 ( 
.A(n_3367),
.B(n_3155),
.Y(n_3389)
);

OAI211xp5_ASAP7_75t_L g3390 ( 
.A1(n_3369),
.A2(n_3152),
.B(n_3200),
.C(n_3214),
.Y(n_3390)
);

OA21x2_ASAP7_75t_L g3391 ( 
.A1(n_3314),
.A2(n_3315),
.B(n_3248),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3279),
.Y(n_3392)
);

CKINVDCx5p33_ASAP7_75t_R g3393 ( 
.A(n_3359),
.Y(n_3393)
);

AOI221xp5_ASAP7_75t_L g3394 ( 
.A1(n_3370),
.A2(n_3152),
.B1(n_3140),
.B2(n_3191),
.C(n_3135),
.Y(n_3394)
);

OAI22xp5_ASAP7_75t_L g3395 ( 
.A1(n_3351),
.A2(n_3218),
.B1(n_3214),
.B2(n_3179),
.Y(n_3395)
);

AOI22xp33_ASAP7_75t_L g3396 ( 
.A1(n_3284),
.A2(n_3026),
.B1(n_3134),
.B2(n_3137),
.Y(n_3396)
);

AOI22xp33_ASAP7_75t_L g3397 ( 
.A1(n_3271),
.A2(n_3134),
.B1(n_3133),
.B2(n_3063),
.Y(n_3397)
);

AOI22xp33_ASAP7_75t_L g3398 ( 
.A1(n_3340),
.A2(n_3133),
.B1(n_3063),
.B2(n_3054),
.Y(n_3398)
);

AOI21xp5_ASAP7_75t_L g3399 ( 
.A1(n_3379),
.A2(n_3100),
.B(n_3112),
.Y(n_3399)
);

AND2x2_ASAP7_75t_L g3400 ( 
.A(n_3249),
.B(n_3043),
.Y(n_3400)
);

OAI21x1_ASAP7_75t_L g3401 ( 
.A1(n_3274),
.A2(n_2801),
.B(n_2944),
.Y(n_3401)
);

BUFx2_ASAP7_75t_L g3402 ( 
.A(n_3275),
.Y(n_3402)
);

AND2x2_ASAP7_75t_L g3403 ( 
.A(n_3333),
.B(n_3075),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_3310),
.Y(n_3404)
);

AOI22xp33_ASAP7_75t_L g3405 ( 
.A1(n_3340),
.A2(n_3054),
.B1(n_3128),
.B2(n_3193),
.Y(n_3405)
);

OAI22xp33_ASAP7_75t_L g3406 ( 
.A1(n_3264),
.A2(n_3062),
.B1(n_3100),
.B2(n_3093),
.Y(n_3406)
);

AOI22xp33_ASAP7_75t_SL g3407 ( 
.A1(n_3340),
.A2(n_3198),
.B1(n_3077),
.B2(n_3121),
.Y(n_3407)
);

OA21x2_ASAP7_75t_L g3408 ( 
.A1(n_3314),
.A2(n_3138),
.B(n_3179),
.Y(n_3408)
);

INVx3_ASAP7_75t_L g3409 ( 
.A(n_3257),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3292),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3292),
.Y(n_3411)
);

AOI211xp5_ASAP7_75t_L g3412 ( 
.A1(n_3273),
.A2(n_3194),
.B(n_3112),
.C(n_3168),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3220),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3220),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_SL g3415 ( 
.A(n_3317),
.B(n_3162),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3252),
.Y(n_3416)
);

AOI22xp33_ASAP7_75t_SL g3417 ( 
.A1(n_3368),
.A2(n_3050),
.B1(n_3204),
.B2(n_3136),
.Y(n_3417)
);

AND2x4_ASAP7_75t_L g3418 ( 
.A(n_3367),
.B(n_3227),
.Y(n_3418)
);

AND2x2_ASAP7_75t_L g3419 ( 
.A(n_3333),
.B(n_3095),
.Y(n_3419)
);

AO21x2_ASAP7_75t_L g3420 ( 
.A1(n_3261),
.A2(n_3194),
.B(n_3176),
.Y(n_3420)
);

AOI22xp33_ASAP7_75t_L g3421 ( 
.A1(n_3345),
.A2(n_3128),
.B1(n_3218),
.B2(n_3183),
.Y(n_3421)
);

AOI22xp33_ASAP7_75t_L g3422 ( 
.A1(n_3345),
.A2(n_3183),
.B1(n_3199),
.B2(n_3086),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3252),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_3250),
.B(n_3123),
.Y(n_3424)
);

AOI22xp33_ASAP7_75t_L g3425 ( 
.A1(n_3350),
.A2(n_3086),
.B1(n_3079),
.B2(n_3018),
.Y(n_3425)
);

AND2x2_ASAP7_75t_L g3426 ( 
.A(n_3250),
.B(n_3092),
.Y(n_3426)
);

OAI21x1_ASAP7_75t_L g3427 ( 
.A1(n_3274),
.A2(n_3124),
.B(n_2832),
.Y(n_3427)
);

OAI22xp5_ASAP7_75t_L g3428 ( 
.A1(n_3317),
.A2(n_3076),
.B1(n_3092),
.B2(n_3088),
.Y(n_3428)
);

OAI22xp33_ASAP7_75t_L g3429 ( 
.A1(n_3358),
.A2(n_3204),
.B1(n_3069),
.B2(n_3080),
.Y(n_3429)
);

AOI22xp33_ASAP7_75t_L g3430 ( 
.A1(n_3350),
.A2(n_3079),
.B1(n_3185),
.B2(n_3078),
.Y(n_3430)
);

OA21x2_ASAP7_75t_L g3431 ( 
.A1(n_3315),
.A2(n_2912),
.B(n_3098),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_L g3432 ( 
.A(n_3233),
.B(n_3066),
.Y(n_3432)
);

AO22x1_ASAP7_75t_L g3433 ( 
.A1(n_3275),
.A2(n_3161),
.B1(n_3155),
.B2(n_3129),
.Y(n_3433)
);

BUFx6f_ASAP7_75t_L g3434 ( 
.A(n_3233),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_3227),
.B(n_3055),
.Y(n_3435)
);

OAI221xp5_ASAP7_75t_L g3436 ( 
.A1(n_3342),
.A2(n_3076),
.B1(n_3274),
.B2(n_3361),
.C(n_3344),
.Y(n_3436)
);

OAI221xp5_ASAP7_75t_L g3437 ( 
.A1(n_3344),
.A2(n_3168),
.B1(n_3109),
.B2(n_3078),
.C(n_3099),
.Y(n_3437)
);

NAND2x1p5_ASAP7_75t_L g3438 ( 
.A(n_3377),
.B(n_3089),
.Y(n_3438)
);

BUFx6f_ASAP7_75t_L g3439 ( 
.A(n_3287),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3253),
.Y(n_3440)
);

AOI22xp33_ASAP7_75t_L g3441 ( 
.A1(n_3377),
.A2(n_3069),
.B1(n_3088),
.B2(n_3099),
.Y(n_3441)
);

OAI21x1_ASAP7_75t_L g3442 ( 
.A1(n_3256),
.A2(n_3268),
.B(n_3244),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3341),
.B(n_3166),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_SL g3444 ( 
.A(n_3308),
.B(n_3091),
.Y(n_3444)
);

OR2x2_ASAP7_75t_L g3445 ( 
.A(n_3297),
.B(n_3113),
.Y(n_3445)
);

NAND3xp33_ASAP7_75t_L g3446 ( 
.A(n_3377),
.B(n_3091),
.C(n_2873),
.Y(n_3446)
);

AOI33xp33_ASAP7_75t_L g3447 ( 
.A1(n_3341),
.A2(n_3189),
.A3(n_2873),
.B1(n_2894),
.B2(n_2893),
.B3(n_2960),
.Y(n_3447)
);

OAI22xp5_ASAP7_75t_L g3448 ( 
.A1(n_3287),
.A2(n_2951),
.B1(n_2845),
.B2(n_2890),
.Y(n_3448)
);

AOI22xp33_ASAP7_75t_L g3449 ( 
.A1(n_3289),
.A2(n_3171),
.B1(n_3182),
.B2(n_2981),
.Y(n_3449)
);

AOI22xp5_ASAP7_75t_L g3450 ( 
.A1(n_3367),
.A2(n_3060),
.B1(n_2951),
.B2(n_2890),
.Y(n_3450)
);

AOI22xp33_ASAP7_75t_L g3451 ( 
.A1(n_3289),
.A2(n_2886),
.B1(n_3022),
.B2(n_3150),
.Y(n_3451)
);

AOI222xp33_ASAP7_75t_L g3452 ( 
.A1(n_3368),
.A2(n_3308),
.B1(n_3235),
.B2(n_3263),
.C1(n_3330),
.C2(n_3371),
.Y(n_3452)
);

OAI211xp5_ASAP7_75t_L g3453 ( 
.A1(n_3377),
.A2(n_2908),
.B(n_3196),
.C(n_2956),
.Y(n_3453)
);

AOI22xp33_ASAP7_75t_L g3454 ( 
.A1(n_3374),
.A2(n_2915),
.B1(n_2914),
.B2(n_2953),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3310),
.Y(n_3455)
);

OAI221xp5_ASAP7_75t_L g3456 ( 
.A1(n_3289),
.A2(n_3150),
.B1(n_3055),
.B2(n_3116),
.C(n_2841),
.Y(n_3456)
);

OA21x2_ASAP7_75t_L g3457 ( 
.A1(n_3301),
.A2(n_2912),
.B(n_2914),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3253),
.Y(n_3458)
);

AOI21xp33_ASAP7_75t_SL g3459 ( 
.A1(n_3359),
.A2(n_3150),
.B(n_2982),
.Y(n_3459)
);

OAI211xp5_ASAP7_75t_L g3460 ( 
.A1(n_3374),
.A2(n_2956),
.B(n_2960),
.C(n_2953),
.Y(n_3460)
);

BUFx5_ASAP7_75t_L g3461 ( 
.A(n_3352),
.Y(n_3461)
);

AOI21xp33_ASAP7_75t_L g3462 ( 
.A1(n_3289),
.A2(n_3096),
.B(n_3089),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3319),
.B(n_3089),
.Y(n_3463)
);

CKINVDCx5p33_ASAP7_75t_R g3464 ( 
.A(n_3235),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3303),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3303),
.Y(n_3466)
);

BUFx2_ASAP7_75t_L g3467 ( 
.A(n_3362),
.Y(n_3467)
);

OAI221xp5_ASAP7_75t_L g3468 ( 
.A1(n_3221),
.A2(n_2833),
.B1(n_2969),
.B2(n_2791),
.C(n_2871),
.Y(n_3468)
);

NOR3xp33_ASAP7_75t_L g3469 ( 
.A(n_3365),
.B(n_2982),
.C(n_2978),
.Y(n_3469)
);

OA21x2_ASAP7_75t_L g3470 ( 
.A1(n_3301),
.A2(n_3003),
.B(n_3015),
.Y(n_3470)
);

OR2x2_ASAP7_75t_L g3471 ( 
.A(n_3326),
.B(n_3096),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3304),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3304),
.Y(n_3473)
);

OAI211xp5_ASAP7_75t_L g3474 ( 
.A1(n_3371),
.A2(n_2960),
.B(n_2969),
.C(n_2833),
.Y(n_3474)
);

OA21x2_ASAP7_75t_L g3475 ( 
.A1(n_3335),
.A2(n_3003),
.B(n_3015),
.Y(n_3475)
);

AOI222xp33_ASAP7_75t_L g3476 ( 
.A1(n_3263),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.C1(n_139),
.C2(n_140),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3323),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3305),
.Y(n_3478)
);

AOI22xp33_ASAP7_75t_L g3479 ( 
.A1(n_3261),
.A2(n_2978),
.B1(n_2966),
.B2(n_2968),
.Y(n_3479)
);

OAI22xp5_ASAP7_75t_L g3480 ( 
.A1(n_3287),
.A2(n_2906),
.B1(n_2791),
.B2(n_2918),
.Y(n_3480)
);

HB1xp67_ASAP7_75t_L g3481 ( 
.A(n_3219),
.Y(n_3481)
);

AOI22xp33_ASAP7_75t_L g3482 ( 
.A1(n_3261),
.A2(n_2949),
.B1(n_2942),
.B2(n_2871),
.Y(n_3482)
);

AOI22xp33_ASAP7_75t_L g3483 ( 
.A1(n_3330),
.A2(n_2942),
.B1(n_2906),
.B2(n_2933),
.Y(n_3483)
);

INVx5_ASAP7_75t_SL g3484 ( 
.A(n_3287),
.Y(n_3484)
);

AOI221xp5_ASAP7_75t_L g3485 ( 
.A1(n_3372),
.A2(n_3096),
.B1(n_2933),
.B2(n_2866),
.C(n_143),
.Y(n_3485)
);

BUFx3_ASAP7_75t_L g3486 ( 
.A(n_3287),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3305),
.Y(n_3487)
);

OAI22xp5_ASAP7_75t_L g3488 ( 
.A1(n_3321),
.A2(n_2906),
.B1(n_3002),
.B2(n_2918),
.Y(n_3488)
);

AOI22xp33_ASAP7_75t_L g3489 ( 
.A1(n_3372),
.A2(n_2866),
.B1(n_2933),
.B2(n_2888),
.Y(n_3489)
);

OAI211xp5_ASAP7_75t_L g3490 ( 
.A1(n_3375),
.A2(n_3376),
.B(n_3281),
.C(n_3366),
.Y(n_3490)
);

AOI21xp5_ASAP7_75t_L g3491 ( 
.A1(n_3360),
.A2(n_3002),
.B(n_2991),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3223),
.Y(n_3492)
);

AOI22xp33_ASAP7_75t_L g3493 ( 
.A1(n_3375),
.A2(n_2866),
.B1(n_2933),
.B2(n_2888),
.Y(n_3493)
);

CKINVDCx5p33_ASAP7_75t_R g3494 ( 
.A(n_3321),
.Y(n_3494)
);

AOI221xp5_ASAP7_75t_L g3495 ( 
.A1(n_3376),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.C(n_144),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3241),
.B(n_2832),
.Y(n_3496)
);

OAI22xp5_ASAP7_75t_L g3497 ( 
.A1(n_3321),
.A2(n_3367),
.B1(n_3241),
.B2(n_3237),
.Y(n_3497)
);

BUFx6f_ASAP7_75t_L g3498 ( 
.A(n_3321),
.Y(n_3498)
);

OAI221xp5_ASAP7_75t_L g3499 ( 
.A1(n_3334),
.A2(n_2909),
.B1(n_2888),
.B2(n_146),
.C(n_147),
.Y(n_3499)
);

AOI221xp5_ASAP7_75t_L g3500 ( 
.A1(n_3316),
.A2(n_141),
.B1(n_144),
.B2(n_147),
.C(n_148),
.Y(n_3500)
);

AOI221xp5_ASAP7_75t_SL g3501 ( 
.A1(n_3366),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.C(n_151),
.Y(n_3501)
);

AND2x4_ASAP7_75t_L g3502 ( 
.A(n_3362),
.B(n_2991),
.Y(n_3502)
);

OR2x2_ASAP7_75t_L g3503 ( 
.A(n_3225),
.B(n_3013),
.Y(n_3503)
);

AOI21x1_ASAP7_75t_L g3504 ( 
.A1(n_3378),
.A2(n_149),
.B(n_152),
.Y(n_3504)
);

INVx2_ASAP7_75t_L g3505 ( 
.A(n_3323),
.Y(n_3505)
);

AOI22xp33_ASAP7_75t_L g3506 ( 
.A1(n_3321),
.A2(n_157),
.B1(n_154),
.B2(n_155),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3255),
.B(n_154),
.Y(n_3507)
);

AOI22xp33_ASAP7_75t_L g3508 ( 
.A1(n_3339),
.A2(n_3343),
.B1(n_3349),
.B2(n_3237),
.Y(n_3508)
);

INVx3_ASAP7_75t_L g3509 ( 
.A(n_3257),
.Y(n_3509)
);

INVxp33_ASAP7_75t_L g3510 ( 
.A(n_3255),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3223),
.Y(n_3511)
);

AOI22xp33_ASAP7_75t_L g3512 ( 
.A1(n_3339),
.A2(n_158),
.B1(n_155),
.B2(n_157),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3323),
.Y(n_3513)
);

INVx2_ASAP7_75t_SL g3514 ( 
.A(n_3434),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3402),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3413),
.Y(n_3516)
);

OR2x2_ASAP7_75t_L g3517 ( 
.A(n_3383),
.B(n_3316),
.Y(n_3517)
);

AOI22xp33_ASAP7_75t_SL g3518 ( 
.A1(n_3380),
.A2(n_3256),
.B1(n_3355),
.B2(n_3348),
.Y(n_3518)
);

NOR2xp33_ASAP7_75t_L g3519 ( 
.A(n_3434),
.B(n_3343),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_3418),
.B(n_3302),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3461),
.Y(n_3521)
);

OR2x2_ASAP7_75t_L g3522 ( 
.A(n_3383),
.B(n_3281),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3414),
.Y(n_3523)
);

AND2x2_ASAP7_75t_L g3524 ( 
.A(n_3418),
.B(n_3302),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3416),
.Y(n_3525)
);

AND2x2_ASAP7_75t_L g3526 ( 
.A(n_3426),
.B(n_3357),
.Y(n_3526)
);

INVxp67_ASAP7_75t_L g3527 ( 
.A(n_3481),
.Y(n_3527)
);

AND2x2_ASAP7_75t_L g3528 ( 
.A(n_3467),
.B(n_3357),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3409),
.B(n_3509),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3423),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3440),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3394),
.B(n_3319),
.Y(n_3532)
);

NAND2x1p5_ASAP7_75t_L g3533 ( 
.A(n_3401),
.B(n_3362),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3388),
.B(n_3349),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3458),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3461),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3409),
.B(n_3337),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3465),
.Y(n_3538)
);

BUFx2_ASAP7_75t_L g3539 ( 
.A(n_3434),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3461),
.Y(n_3540)
);

INVx2_ASAP7_75t_L g3541 ( 
.A(n_3461),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3461),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_3461),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3408),
.B(n_3338),
.Y(n_3544)
);

INVx3_ASAP7_75t_L g3545 ( 
.A(n_3439),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3466),
.Y(n_3546)
);

OR2x2_ASAP7_75t_L g3547 ( 
.A(n_3420),
.B(n_3226),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_3509),
.B(n_3337),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3472),
.Y(n_3549)
);

AO22x1_ASAP7_75t_L g3550 ( 
.A1(n_3395),
.A2(n_3230),
.B1(n_3300),
.B2(n_3257),
.Y(n_3550)
);

HB1xp67_ASAP7_75t_L g3551 ( 
.A(n_3481),
.Y(n_3551)
);

OAI221xp5_ASAP7_75t_L g3552 ( 
.A1(n_3386),
.A2(n_3335),
.B1(n_3256),
.B2(n_3237),
.C(n_3347),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_3438),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3473),
.Y(n_3554)
);

OR2x2_ASAP7_75t_L g3555 ( 
.A(n_3420),
.B(n_3226),
.Y(n_3555)
);

INVx2_ASAP7_75t_SL g3556 ( 
.A(n_3434),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3408),
.B(n_3338),
.Y(n_3557)
);

INVx2_ASAP7_75t_L g3558 ( 
.A(n_3438),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_3439),
.Y(n_3559)
);

NOR2xp67_ASAP7_75t_L g3560 ( 
.A(n_3490),
.B(n_3300),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3508),
.B(n_3348),
.Y(n_3561)
);

AND2x4_ASAP7_75t_L g3562 ( 
.A(n_3389),
.B(n_3346),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3478),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3439),
.Y(n_3564)
);

HB1xp67_ASAP7_75t_L g3565 ( 
.A(n_3384),
.Y(n_3565)
);

AND2x4_ASAP7_75t_SL g3566 ( 
.A(n_3389),
.B(n_3387),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3386),
.B(n_3392),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3487),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3492),
.Y(n_3569)
);

INVxp67_ASAP7_75t_L g3570 ( 
.A(n_3452),
.Y(n_3570)
);

AND2x2_ASAP7_75t_L g3571 ( 
.A(n_3508),
.B(n_3355),
.Y(n_3571)
);

OR2x2_ASAP7_75t_L g3572 ( 
.A(n_3384),
.B(n_3225),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3511),
.Y(n_3573)
);

AND2x4_ASAP7_75t_L g3574 ( 
.A(n_3439),
.B(n_3346),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3498),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3435),
.B(n_3300),
.Y(n_3576)
);

HB1xp67_ASAP7_75t_L g3577 ( 
.A(n_3410),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3411),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3498),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3405),
.B(n_3399),
.Y(n_3580)
);

INVx2_ASAP7_75t_SL g3581 ( 
.A(n_3498),
.Y(n_3581)
);

AND2x2_ASAP7_75t_L g3582 ( 
.A(n_3400),
.B(n_3363),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3498),
.Y(n_3583)
);

INVx2_ASAP7_75t_L g3584 ( 
.A(n_3503),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_3510),
.B(n_3373),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_3382),
.Y(n_3586)
);

AND2x2_ASAP7_75t_L g3587 ( 
.A(n_3404),
.B(n_3332),
.Y(n_3587)
);

CKINVDCx14_ASAP7_75t_R g3588 ( 
.A(n_3393),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3471),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3445),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3455),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3405),
.B(n_3336),
.Y(n_3592)
);

INVxp67_ASAP7_75t_L g3593 ( 
.A(n_3444),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_3477),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_SL g3595 ( 
.A(n_3406),
.B(n_3346),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3385),
.B(n_3336),
.Y(n_3596)
);

AND2x2_ASAP7_75t_L g3597 ( 
.A(n_3505),
.B(n_3513),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3486),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3463),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3403),
.B(n_3332),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3443),
.Y(n_3601)
);

BUFx2_ASAP7_75t_L g3602 ( 
.A(n_3391),
.Y(n_3602)
);

AND2x4_ASAP7_75t_L g3603 ( 
.A(n_3427),
.B(n_3346),
.Y(n_3603)
);

AND2x4_ASAP7_75t_L g3604 ( 
.A(n_3469),
.B(n_3352),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3385),
.B(n_3307),
.Y(n_3605)
);

AND2x2_ASAP7_75t_L g3606 ( 
.A(n_3391),
.B(n_3269),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3398),
.B(n_3307),
.Y(n_3607)
);

BUFx2_ASAP7_75t_L g3608 ( 
.A(n_3494),
.Y(n_3608)
);

INVx2_ASAP7_75t_L g3609 ( 
.A(n_3442),
.Y(n_3609)
);

AND2x4_ASAP7_75t_L g3610 ( 
.A(n_3469),
.B(n_3258),
.Y(n_3610)
);

AND2x4_ASAP7_75t_L g3611 ( 
.A(n_3450),
.B(n_3258),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3504),
.Y(n_3612)
);

AOI22xp33_ASAP7_75t_L g3613 ( 
.A1(n_3398),
.A2(n_3237),
.B1(n_3365),
.B2(n_3325),
.Y(n_3613)
);

OR2x2_ASAP7_75t_L g3614 ( 
.A(n_3446),
.B(n_3298),
.Y(n_3614)
);

INVx2_ASAP7_75t_L g3615 ( 
.A(n_3496),
.Y(n_3615)
);

AOI22xp33_ASAP7_75t_SL g3616 ( 
.A1(n_3390),
.A2(n_3237),
.B1(n_3325),
.B2(n_3313),
.Y(n_3616)
);

AND2x4_ASAP7_75t_L g3617 ( 
.A(n_3419),
.B(n_3258),
.Y(n_3617)
);

BUFx2_ASAP7_75t_L g3618 ( 
.A(n_3433),
.Y(n_3618)
);

OR2x2_ASAP7_75t_L g3619 ( 
.A(n_3436),
.B(n_3298),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3447),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3507),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_L g3622 ( 
.A(n_3432),
.B(n_3318),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_3497),
.B(n_3269),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3396),
.B(n_3295),
.Y(n_3624)
);

AND2x2_ASAP7_75t_L g3625 ( 
.A(n_3484),
.B(n_3283),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3474),
.Y(n_3626)
);

AND2x2_ASAP7_75t_L g3627 ( 
.A(n_3484),
.B(n_3283),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3484),
.Y(n_3628)
);

AND2x4_ASAP7_75t_L g3629 ( 
.A(n_3502),
.B(n_3258),
.Y(n_3629)
);

OR2x2_ASAP7_75t_L g3630 ( 
.A(n_3453),
.B(n_3299),
.Y(n_3630)
);

AND2x2_ASAP7_75t_L g3631 ( 
.A(n_3424),
.B(n_3407),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3396),
.B(n_3295),
.Y(n_3632)
);

AND2x2_ASAP7_75t_L g3633 ( 
.A(n_3407),
.B(n_3285),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3437),
.Y(n_3634)
);

INVxp67_ASAP7_75t_L g3635 ( 
.A(n_3415),
.Y(n_3635)
);

OAI222xp33_ASAP7_75t_L g3636 ( 
.A1(n_3397),
.A2(n_3353),
.B1(n_3294),
.B2(n_3285),
.C1(n_3328),
.C2(n_3320),
.Y(n_3636)
);

BUFx3_ASAP7_75t_L g3637 ( 
.A(n_3464),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3425),
.B(n_3260),
.Y(n_3638)
);

INVx3_ASAP7_75t_L g3639 ( 
.A(n_3502),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_SL g3640 ( 
.A(n_3406),
.B(n_3353),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_3462),
.B(n_3294),
.Y(n_3641)
);

HB1xp67_ASAP7_75t_L g3642 ( 
.A(n_3431),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3551),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3608),
.Y(n_3644)
);

NAND3xp33_ASAP7_75t_L g3645 ( 
.A(n_3640),
.B(n_3476),
.C(n_3501),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3608),
.Y(n_3646)
);

AND2x2_ASAP7_75t_L g3647 ( 
.A(n_3526),
.B(n_3265),
.Y(n_3647)
);

INVx3_ASAP7_75t_L g3648 ( 
.A(n_3566),
.Y(n_3648)
);

AOI22xp33_ASAP7_75t_L g3649 ( 
.A1(n_3595),
.A2(n_3397),
.B1(n_3381),
.B2(n_3417),
.Y(n_3649)
);

OA21x2_ASAP7_75t_L g3650 ( 
.A1(n_3640),
.A2(n_3493),
.B(n_3489),
.Y(n_3650)
);

OAI21x1_ASAP7_75t_L g3651 ( 
.A1(n_3533),
.A2(n_3493),
.B(n_3489),
.Y(n_3651)
);

AOI33xp33_ASAP7_75t_L g3652 ( 
.A1(n_3616),
.A2(n_3381),
.A3(n_3421),
.B1(n_3412),
.B2(n_3417),
.B3(n_3422),
.Y(n_3652)
);

OAI211xp5_ASAP7_75t_SL g3653 ( 
.A1(n_3580),
.A2(n_3595),
.B(n_3570),
.C(n_3634),
.Y(n_3653)
);

OAI33xp33_ASAP7_75t_L g3654 ( 
.A1(n_3620),
.A2(n_3429),
.A3(n_3428),
.B1(n_3448),
.B2(n_3228),
.B3(n_3242),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3577),
.Y(n_3655)
);

AOI211xp5_ASAP7_75t_L g3656 ( 
.A1(n_3550),
.A2(n_3429),
.B(n_3499),
.C(n_3485),
.Y(n_3656)
);

AOI221xp5_ASAP7_75t_L g3657 ( 
.A1(n_3626),
.A2(n_3421),
.B1(n_3495),
.B2(n_3500),
.C(n_3422),
.Y(n_3657)
);

INVxp67_ASAP7_75t_L g3658 ( 
.A(n_3618),
.Y(n_3658)
);

OR2x2_ASAP7_75t_L g3659 ( 
.A(n_3607),
.B(n_3425),
.Y(n_3659)
);

BUFx3_ASAP7_75t_L g3660 ( 
.A(n_3637),
.Y(n_3660)
);

OAI33xp33_ASAP7_75t_L g3661 ( 
.A1(n_3567),
.A2(n_3224),
.A3(n_3228),
.B1(n_3242),
.B2(n_3309),
.B3(n_3278),
.Y(n_3661)
);

INVx2_ASAP7_75t_L g3662 ( 
.A(n_3545),
.Y(n_3662)
);

NOR2x1p5_ASAP7_75t_L g3663 ( 
.A(n_3637),
.B(n_3456),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3565),
.Y(n_3664)
);

AOI22xp33_ASAP7_75t_L g3665 ( 
.A1(n_3618),
.A2(n_3441),
.B1(n_3430),
.B2(n_3468),
.Y(n_3665)
);

HB1xp67_ASAP7_75t_L g3666 ( 
.A(n_3515),
.Y(n_3666)
);

NAND2xp33_ASAP7_75t_SL g3667 ( 
.A(n_3631),
.B(n_3506),
.Y(n_3667)
);

OAI222xp33_ASAP7_75t_L g3668 ( 
.A1(n_3518),
.A2(n_3441),
.B1(n_3430),
.B2(n_3451),
.C1(n_3449),
.C2(n_3512),
.Y(n_3668)
);

NOR2xp33_ASAP7_75t_L g3669 ( 
.A(n_3588),
.B(n_3459),
.Y(n_3669)
);

OR2x2_ASAP7_75t_L g3670 ( 
.A(n_3605),
.B(n_3260),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3545),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3526),
.B(n_3265),
.Y(n_3672)
);

AND2x2_ASAP7_75t_L g3673 ( 
.A(n_3566),
.B(n_3276),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3516),
.Y(n_3674)
);

NOR2xp33_ASAP7_75t_L g3675 ( 
.A(n_3588),
.B(n_3378),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3523),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_SL g3677 ( 
.A(n_3635),
.B(n_3480),
.Y(n_3677)
);

AND2x2_ASAP7_75t_L g3678 ( 
.A(n_3528),
.B(n_3276),
.Y(n_3678)
);

INVx5_ASAP7_75t_L g3679 ( 
.A(n_3602),
.Y(n_3679)
);

AND2x2_ASAP7_75t_L g3680 ( 
.A(n_3528),
.B(n_3291),
.Y(n_3680)
);

NAND3xp33_ASAP7_75t_L g3681 ( 
.A(n_3593),
.B(n_3506),
.C(n_3512),
.Y(n_3681)
);

AO21x2_ASAP7_75t_L g3682 ( 
.A1(n_3560),
.A2(n_3460),
.B(n_3491),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3525),
.Y(n_3683)
);

INVxp67_ASAP7_75t_L g3684 ( 
.A(n_3539),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3530),
.Y(n_3685)
);

AOI22xp33_ASAP7_75t_L g3686 ( 
.A1(n_3631),
.A2(n_3479),
.B1(n_3483),
.B2(n_3431),
.Y(n_3686)
);

OR2x2_ASAP7_75t_L g3687 ( 
.A(n_3592),
.B(n_3262),
.Y(n_3687)
);

AO21x2_ASAP7_75t_L g3688 ( 
.A1(n_3636),
.A2(n_3234),
.B(n_3244),
.Y(n_3688)
);

AOI222xp33_ASAP7_75t_L g3689 ( 
.A1(n_3532),
.A2(n_3483),
.B1(n_3479),
.B2(n_3482),
.C1(n_3454),
.C2(n_3488),
.Y(n_3689)
);

OAI21xp5_ASAP7_75t_L g3690 ( 
.A1(n_3612),
.A2(n_3482),
.B(n_3454),
.Y(n_3690)
);

OAI21x1_ASAP7_75t_L g3691 ( 
.A1(n_3533),
.A2(n_3306),
.B(n_3268),
.Y(n_3691)
);

INVx1_ASAP7_75t_SL g3692 ( 
.A(n_3633),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3545),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_SL g3694 ( 
.A(n_3633),
.B(n_3328),
.Y(n_3694)
);

OAI21xp33_ASAP7_75t_L g3695 ( 
.A1(n_3613),
.A2(n_3278),
.B(n_3262),
.Y(n_3695)
);

AO21x2_ASAP7_75t_L g3696 ( 
.A1(n_3642),
.A2(n_3234),
.B(n_3224),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3514),
.Y(n_3697)
);

AO21x2_ASAP7_75t_L g3698 ( 
.A1(n_3544),
.A2(n_3234),
.B(n_3325),
.Y(n_3698)
);

AND2x4_ASAP7_75t_L g3699 ( 
.A(n_3514),
.B(n_3327),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3527),
.B(n_3280),
.Y(n_3700)
);

AND2x4_ASAP7_75t_L g3701 ( 
.A(n_3556),
.B(n_3327),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3531),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3535),
.Y(n_3703)
);

HB1xp67_ASAP7_75t_L g3704 ( 
.A(n_3515),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3538),
.Y(n_3705)
);

OAI221xp5_ASAP7_75t_L g3706 ( 
.A1(n_3596),
.A2(n_3313),
.B1(n_3331),
.B2(n_3457),
.C(n_3243),
.Y(n_3706)
);

HB1xp67_ASAP7_75t_L g3707 ( 
.A(n_3602),
.Y(n_3707)
);

NOR2xp33_ASAP7_75t_L g3708 ( 
.A(n_3621),
.B(n_3309),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3601),
.B(n_3280),
.Y(n_3709)
);

OAI221xp5_ASAP7_75t_L g3710 ( 
.A1(n_3552),
.A2(n_3313),
.B1(n_3457),
.B2(n_3243),
.C(n_3288),
.Y(n_3710)
);

NAND3xp33_ASAP7_75t_L g3711 ( 
.A(n_3638),
.B(n_3313),
.C(n_3243),
.Y(n_3711)
);

OR2x6_ASAP7_75t_L g3712 ( 
.A(n_3556),
.B(n_3628),
.Y(n_3712)
);

AO21x2_ASAP7_75t_L g3713 ( 
.A1(n_3557),
.A2(n_3288),
.B(n_3282),
.Y(n_3713)
);

NAND4xp25_ASAP7_75t_L g3714 ( 
.A(n_3624),
.B(n_3282),
.C(n_3296),
.D(n_3246),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3639),
.Y(n_3715)
);

OR2x2_ASAP7_75t_L g3716 ( 
.A(n_3590),
.B(n_3299),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3546),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3549),
.Y(n_3718)
);

AO21x1_ASAP7_75t_SL g3719 ( 
.A1(n_3632),
.A2(n_3246),
.B(n_3245),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3554),
.Y(n_3720)
);

OAI33xp33_ASAP7_75t_L g3721 ( 
.A1(n_3614),
.A2(n_3251),
.A3(n_3245),
.B1(n_3296),
.B2(n_3238),
.B3(n_3222),
.Y(n_3721)
);

OAI321xp33_ASAP7_75t_L g3722 ( 
.A1(n_3619),
.A2(n_3251),
.A3(n_3324),
.B1(n_3322),
.B2(n_3222),
.C(n_3236),
.Y(n_3722)
);

OAI221xp5_ASAP7_75t_L g3723 ( 
.A1(n_3619),
.A2(n_3324),
.B1(n_3322),
.B2(n_3239),
.C(n_3236),
.Y(n_3723)
);

AOI33xp33_ASAP7_75t_L g3724 ( 
.A1(n_3561),
.A2(n_3238),
.A3(n_3239),
.B1(n_3247),
.B2(n_3277),
.B3(n_3272),
.Y(n_3724)
);

AOI33xp33_ASAP7_75t_L g3725 ( 
.A1(n_3561),
.A2(n_3247),
.A3(n_3293),
.B1(n_3290),
.B2(n_3277),
.B3(n_3272),
.Y(n_3725)
);

NOR2xp67_ASAP7_75t_L g3726 ( 
.A(n_3520),
.B(n_3254),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3576),
.B(n_3291),
.Y(n_3727)
);

HB1xp67_ASAP7_75t_L g3728 ( 
.A(n_3572),
.Y(n_3728)
);

CKINVDCx5p33_ASAP7_75t_R g3729 ( 
.A(n_3628),
.Y(n_3729)
);

AND2x4_ASAP7_75t_L g3730 ( 
.A(n_3617),
.B(n_3254),
.Y(n_3730)
);

BUFx3_ASAP7_75t_L g3731 ( 
.A(n_3598),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3563),
.Y(n_3732)
);

AND2x4_ASAP7_75t_L g3733 ( 
.A(n_3617),
.B(n_3259),
.Y(n_3733)
);

NAND3xp33_ASAP7_75t_SL g3734 ( 
.A(n_3614),
.B(n_3267),
.C(n_3259),
.Y(n_3734)
);

OAI21xp5_ASAP7_75t_L g3735 ( 
.A1(n_3630),
.A2(n_3311),
.B(n_3306),
.Y(n_3735)
);

BUFx2_ASAP7_75t_L g3736 ( 
.A(n_3617),
.Y(n_3736)
);

NAND2xp33_ASAP7_75t_R g3737 ( 
.A(n_3623),
.B(n_3630),
.Y(n_3737)
);

AOI22xp33_ASAP7_75t_L g3738 ( 
.A1(n_3589),
.A2(n_3356),
.B1(n_3311),
.B2(n_3243),
.Y(n_3738)
);

INVxp67_ASAP7_75t_L g3739 ( 
.A(n_3519),
.Y(n_3739)
);

OAI221xp5_ASAP7_75t_L g3740 ( 
.A1(n_3522),
.A2(n_3475),
.B1(n_3229),
.B2(n_3293),
.C(n_3290),
.Y(n_3740)
);

AND2x2_ASAP7_75t_L g3741 ( 
.A(n_3576),
.B(n_3267),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_3582),
.B(n_3270),
.Y(n_3742)
);

OR2x2_ASAP7_75t_L g3743 ( 
.A(n_3534),
.B(n_3270),
.Y(n_3743)
);

AOI22xp5_ASAP7_75t_L g3744 ( 
.A1(n_3611),
.A2(n_3356),
.B1(n_3475),
.B2(n_3470),
.Y(n_3744)
);

OR2x6_ASAP7_75t_L g3745 ( 
.A(n_3581),
.B(n_3286),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3639),
.Y(n_3746)
);

OR2x2_ASAP7_75t_L g3747 ( 
.A(n_3599),
.B(n_3356),
.Y(n_3747)
);

NAND3xp33_ASAP7_75t_L g3748 ( 
.A(n_3522),
.B(n_3229),
.C(n_159),
.Y(n_3748)
);

BUFx3_ASAP7_75t_L g3749 ( 
.A(n_3611),
.Y(n_3749)
);

AOI221xp5_ASAP7_75t_L g3750 ( 
.A1(n_3571),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.C(n_162),
.Y(n_3750)
);

INVxp67_ASAP7_75t_L g3751 ( 
.A(n_3622),
.Y(n_3751)
);

NOR2xp33_ASAP7_75t_R g3752 ( 
.A(n_3579),
.B(n_161),
.Y(n_3752)
);

OAI33xp33_ASAP7_75t_L g3753 ( 
.A1(n_3547),
.A2(n_163),
.A3(n_164),
.B1(n_165),
.B2(n_166),
.B3(n_167),
.Y(n_3753)
);

AND2x4_ASAP7_75t_SL g3754 ( 
.A(n_3520),
.B(n_3229),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3568),
.Y(n_3755)
);

OAI21xp5_ASAP7_75t_L g3756 ( 
.A1(n_3547),
.A2(n_3286),
.B(n_3240),
.Y(n_3756)
);

INVx4_ASAP7_75t_L g3757 ( 
.A(n_3559),
.Y(n_3757)
);

OR2x2_ASAP7_75t_L g3758 ( 
.A(n_3692),
.B(n_3572),
.Y(n_3758)
);

AO21x2_ASAP7_75t_L g3759 ( 
.A1(n_3658),
.A2(n_3555),
.B(n_3559),
.Y(n_3759)
);

XNOR2xp5_ASAP7_75t_L g3760 ( 
.A(n_3649),
.B(n_3611),
.Y(n_3760)
);

OAI211xp5_ASAP7_75t_SL g3761 ( 
.A1(n_3652),
.A2(n_3555),
.B(n_3609),
.C(n_3517),
.Y(n_3761)
);

BUFx5_ASAP7_75t_L g3762 ( 
.A(n_3660),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3728),
.Y(n_3763)
);

NOR2x1_ASAP7_75t_L g3764 ( 
.A(n_3645),
.B(n_3564),
.Y(n_3764)
);

NOR3xp33_ASAP7_75t_L g3765 ( 
.A(n_3653),
.B(n_3575),
.C(n_3564),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3657),
.B(n_3585),
.Y(n_3766)
);

NAND3xp33_ASAP7_75t_L g3767 ( 
.A(n_3645),
.B(n_3583),
.C(n_3575),
.Y(n_3767)
);

AND2x2_ASAP7_75t_L g3768 ( 
.A(n_3648),
.B(n_3524),
.Y(n_3768)
);

AOI22xp33_ASAP7_75t_L g3769 ( 
.A1(n_3667),
.A2(n_3689),
.B1(n_3654),
.B2(n_3659),
.Y(n_3769)
);

AOI211x1_ASAP7_75t_L g3770 ( 
.A1(n_3668),
.A2(n_3571),
.B(n_3623),
.C(n_3641),
.Y(n_3770)
);

NOR3xp33_ASAP7_75t_L g3771 ( 
.A(n_3690),
.B(n_3583),
.C(n_3581),
.Y(n_3771)
);

INVxp67_ASAP7_75t_L g3772 ( 
.A(n_3737),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_3644),
.B(n_3585),
.Y(n_3773)
);

OR2x6_ASAP7_75t_L g3774 ( 
.A(n_3646),
.B(n_3712),
.Y(n_3774)
);

NAND4xp75_ASAP7_75t_L g3775 ( 
.A(n_3650),
.B(n_3524),
.C(n_3606),
.D(n_3641),
.Y(n_3775)
);

OR2x2_ASAP7_75t_L g3776 ( 
.A(n_3692),
.B(n_3578),
.Y(n_3776)
);

AOI22xp33_ASAP7_75t_L g3777 ( 
.A1(n_3689),
.A2(n_3562),
.B1(n_3610),
.B2(n_3582),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3648),
.B(n_3537),
.Y(n_3778)
);

OR2x2_ASAP7_75t_L g3779 ( 
.A(n_3751),
.B(n_3684),
.Y(n_3779)
);

NOR3xp33_ASAP7_75t_L g3780 ( 
.A(n_3690),
.B(n_3750),
.C(n_3681),
.Y(n_3780)
);

NOR3xp33_ASAP7_75t_L g3781 ( 
.A(n_3681),
.B(n_3609),
.C(n_3517),
.Y(n_3781)
);

NAND4xp75_ASAP7_75t_L g3782 ( 
.A(n_3650),
.B(n_3606),
.C(n_3627),
.D(n_3625),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_3739),
.B(n_3600),
.Y(n_3783)
);

NAND4xp75_ASAP7_75t_L g3784 ( 
.A(n_3735),
.B(n_3625),
.C(n_3627),
.D(n_3529),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3736),
.B(n_3537),
.Y(n_3785)
);

AND2x4_ASAP7_75t_L g3786 ( 
.A(n_3749),
.B(n_3562),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3707),
.Y(n_3787)
);

NAND4xp75_ASAP7_75t_L g3788 ( 
.A(n_3735),
.B(n_3529),
.C(n_3548),
.D(n_3553),
.Y(n_3788)
);

NAND3xp33_ASAP7_75t_L g3789 ( 
.A(n_3748),
.B(n_3679),
.C(n_3656),
.Y(n_3789)
);

OR2x2_ASAP7_75t_L g3790 ( 
.A(n_3643),
.B(n_3584),
.Y(n_3790)
);

NAND3xp33_ASAP7_75t_L g3791 ( 
.A(n_3748),
.B(n_3604),
.C(n_3610),
.Y(n_3791)
);

INVx2_ASAP7_75t_SL g3792 ( 
.A(n_3712),
.Y(n_3792)
);

AOI221xp5_ASAP7_75t_L g3793 ( 
.A1(n_3665),
.A2(n_3604),
.B1(n_3584),
.B2(n_3610),
.C(n_3573),
.Y(n_3793)
);

OR2x2_ASAP7_75t_L g3794 ( 
.A(n_3664),
.B(n_3569),
.Y(n_3794)
);

OR2x2_ASAP7_75t_L g3795 ( 
.A(n_3666),
.B(n_3548),
.Y(n_3795)
);

NAND4xp75_ASAP7_75t_L g3796 ( 
.A(n_3694),
.B(n_3558),
.C(n_3553),
.D(n_3521),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3704),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3697),
.B(n_3600),
.Y(n_3798)
);

AND2x2_ASAP7_75t_L g3799 ( 
.A(n_3647),
.B(n_3562),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3674),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3672),
.B(n_3587),
.Y(n_3801)
);

NOR3xp33_ASAP7_75t_L g3802 ( 
.A(n_3753),
.B(n_3558),
.C(n_3639),
.Y(n_3802)
);

BUFx3_ASAP7_75t_L g3803 ( 
.A(n_3731),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3729),
.B(n_3587),
.Y(n_3804)
);

AO21x2_ASAP7_75t_L g3805 ( 
.A1(n_3682),
.A2(n_3574),
.B(n_3604),
.Y(n_3805)
);

OA211x2_ASAP7_75t_L g3806 ( 
.A1(n_3669),
.A2(n_3675),
.B(n_3677),
.C(n_3695),
.Y(n_3806)
);

OR2x2_ASAP7_75t_L g3807 ( 
.A(n_3670),
.B(n_3586),
.Y(n_3807)
);

INVx2_ASAP7_75t_L g3808 ( 
.A(n_3679),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_SL g3809 ( 
.A(n_3679),
.B(n_3629),
.Y(n_3809)
);

AOI22xp33_ASAP7_75t_L g3810 ( 
.A1(n_3663),
.A2(n_3629),
.B1(n_3574),
.B2(n_3591),
.Y(n_3810)
);

AND2x2_ASAP7_75t_SL g3811 ( 
.A(n_3686),
.B(n_3574),
.Y(n_3811)
);

AND2x2_ASAP7_75t_L g3812 ( 
.A(n_3673),
.B(n_3678),
.Y(n_3812)
);

NAND4xp75_ASAP7_75t_L g3813 ( 
.A(n_3726),
.B(n_3756),
.C(n_3655),
.D(n_3671),
.Y(n_3813)
);

NAND3xp33_ASAP7_75t_L g3814 ( 
.A(n_3679),
.B(n_3591),
.C(n_3586),
.Y(n_3814)
);

NAND3xp33_ASAP7_75t_L g3815 ( 
.A(n_3757),
.B(n_3594),
.C(n_3615),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_3712),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3680),
.B(n_3594),
.Y(n_3817)
);

AND2x2_ASAP7_75t_L g3818 ( 
.A(n_3727),
.B(n_3629),
.Y(n_3818)
);

HB1xp67_ASAP7_75t_L g3819 ( 
.A(n_3757),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3724),
.B(n_3597),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3708),
.B(n_3597),
.Y(n_3821)
);

NOR3xp33_ASAP7_75t_L g3822 ( 
.A(n_3710),
.B(n_3615),
.C(n_3536),
.Y(n_3822)
);

AOI22xp5_ASAP7_75t_L g3823 ( 
.A1(n_3682),
.A2(n_3603),
.B1(n_3229),
.B2(n_3470),
.Y(n_3823)
);

AOI22xp33_ASAP7_75t_L g3824 ( 
.A1(n_3661),
.A2(n_3603),
.B1(n_3536),
.B2(n_3540),
.Y(n_3824)
);

AND2x2_ASAP7_75t_L g3825 ( 
.A(n_3742),
.B(n_3741),
.Y(n_3825)
);

OAI211xp5_ASAP7_75t_SL g3826 ( 
.A1(n_3710),
.A2(n_3540),
.B(n_3541),
.C(n_3521),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3676),
.Y(n_3827)
);

OAI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_3651),
.A2(n_3603),
.B(n_3542),
.Y(n_3828)
);

NOR3xp33_ASAP7_75t_L g3829 ( 
.A(n_3662),
.B(n_3542),
.C(n_3541),
.Y(n_3829)
);

NAND3xp33_ASAP7_75t_L g3830 ( 
.A(n_3683),
.B(n_3543),
.C(n_163),
.Y(n_3830)
);

AND2x2_ASAP7_75t_L g3831 ( 
.A(n_3730),
.B(n_3543),
.Y(n_3831)
);

AND2x2_ASAP7_75t_L g3832 ( 
.A(n_3730),
.B(n_3232),
.Y(n_3832)
);

INVx2_ASAP7_75t_L g3833 ( 
.A(n_3715),
.Y(n_3833)
);

NAND3xp33_ASAP7_75t_L g3834 ( 
.A(n_3711),
.B(n_166),
.C(n_170),
.Y(n_3834)
);

OR2x2_ASAP7_75t_L g3835 ( 
.A(n_3687),
.B(n_3232),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_SL g3836 ( 
.A(n_3722),
.B(n_3240),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3746),
.Y(n_3837)
);

NAND3xp33_ASAP7_75t_L g3838 ( 
.A(n_3711),
.B(n_170),
.C(n_171),
.Y(n_3838)
);

AND2x4_ASAP7_75t_L g3839 ( 
.A(n_3693),
.B(n_172),
.Y(n_3839)
);

OR2x2_ASAP7_75t_L g3840 ( 
.A(n_3714),
.B(n_172),
.Y(n_3840)
);

NAND4xp75_ASAP7_75t_L g3841 ( 
.A(n_3756),
.B(n_173),
.C(n_174),
.D(n_175),
.Y(n_3841)
);

AOI221xp5_ASAP7_75t_L g3842 ( 
.A1(n_3706),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.C(n_178),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3685),
.B(n_176),
.Y(n_3843)
);

NAND3xp33_ASAP7_75t_L g3844 ( 
.A(n_3702),
.B(n_178),
.C(n_181),
.Y(n_3844)
);

HB1xp67_ASAP7_75t_L g3845 ( 
.A(n_3752),
.Y(n_3845)
);

NAND4xp25_ASAP7_75t_L g3846 ( 
.A(n_3703),
.B(n_183),
.C(n_184),
.D(n_185),
.Y(n_3846)
);

OR2x2_ASAP7_75t_L g3847 ( 
.A(n_3714),
.B(n_184),
.Y(n_3847)
);

AOI22xp33_ASAP7_75t_L g3848 ( 
.A1(n_3721),
.A2(n_1072),
.B1(n_1071),
.B2(n_1070),
.Y(n_3848)
);

OR2x2_ASAP7_75t_L g3849 ( 
.A(n_3716),
.B(n_185),
.Y(n_3849)
);

OAI211xp5_ASAP7_75t_SL g3850 ( 
.A1(n_3738),
.A2(n_186),
.B(n_187),
.C(n_188),
.Y(n_3850)
);

AND2x4_ASAP7_75t_L g3851 ( 
.A(n_3774),
.B(n_3705),
.Y(n_3851)
);

AOI221xp5_ASAP7_75t_L g3852 ( 
.A1(n_3789),
.A2(n_3706),
.B1(n_3722),
.B2(n_3734),
.C(n_3740),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3845),
.B(n_3733),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_3772),
.B(n_3717),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3758),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3787),
.Y(n_3856)
);

BUFx4f_ASAP7_75t_SL g3857 ( 
.A(n_3762),
.Y(n_3857)
);

INVxp67_ASAP7_75t_L g3858 ( 
.A(n_3819),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3763),
.Y(n_3859)
);

AND2x4_ASAP7_75t_L g3860 ( 
.A(n_3774),
.B(n_3718),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3776),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3764),
.B(n_3720),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3780),
.B(n_3732),
.Y(n_3863)
);

OAI33xp33_ASAP7_75t_L g3864 ( 
.A1(n_3761),
.A2(n_3755),
.A3(n_3700),
.B1(n_3709),
.B2(n_3747),
.B3(n_3743),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3768),
.B(n_3733),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3769),
.B(n_3725),
.Y(n_3866)
);

INVx1_ASAP7_75t_SL g3867 ( 
.A(n_3803),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3797),
.Y(n_3868)
);

INVx3_ASAP7_75t_L g3869 ( 
.A(n_3805),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3778),
.B(n_3719),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3805),
.Y(n_3871)
);

OR2x2_ASAP7_75t_L g3872 ( 
.A(n_3779),
.B(n_3700),
.Y(n_3872)
);

NOR2xp33_ASAP7_75t_L g3873 ( 
.A(n_3789),
.B(n_3723),
.Y(n_3873)
);

HB1xp67_ASAP7_75t_L g3874 ( 
.A(n_3759),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3849),
.Y(n_3875)
);

AND2x2_ASAP7_75t_L g3876 ( 
.A(n_3785),
.B(n_3699),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3816),
.B(n_3699),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3812),
.B(n_3701),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3794),
.Y(n_3879)
);

INVx5_ASAP7_75t_L g3880 ( 
.A(n_3774),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3792),
.B(n_3701),
.Y(n_3881)
);

NAND2x1p5_ASAP7_75t_L g3882 ( 
.A(n_3809),
.B(n_3691),
.Y(n_3882)
);

AND2x2_ASAP7_75t_L g3883 ( 
.A(n_3786),
.B(n_3754),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3786),
.B(n_3709),
.Y(n_3884)
);

AND2x4_ASAP7_75t_L g3885 ( 
.A(n_3808),
.B(n_3759),
.Y(n_3885)
);

INVx2_ASAP7_75t_L g3886 ( 
.A(n_3762),
.Y(n_3886)
);

NOR2xp33_ASAP7_75t_L g3887 ( 
.A(n_3766),
.B(n_3713),
.Y(n_3887)
);

NAND4xp25_ASAP7_75t_L g3888 ( 
.A(n_3806),
.B(n_3740),
.C(n_3744),
.D(n_3688),
.Y(n_3888)
);

INVx2_ASAP7_75t_SL g3889 ( 
.A(n_3795),
.Y(n_3889)
);

INVx2_ASAP7_75t_L g3890 ( 
.A(n_3762),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3770),
.B(n_3713),
.Y(n_3891)
);

NAND3xp33_ASAP7_75t_L g3892 ( 
.A(n_3781),
.B(n_3745),
.C(n_3688),
.Y(n_3892)
);

NAND3xp33_ASAP7_75t_L g3893 ( 
.A(n_3771),
.B(n_3745),
.C(n_3698),
.Y(n_3893)
);

AOI22xp33_ASAP7_75t_L g3894 ( 
.A1(n_3806),
.A2(n_3698),
.B1(n_3696),
.B2(n_3745),
.Y(n_3894)
);

OR2x2_ASAP7_75t_L g3895 ( 
.A(n_3773),
.B(n_3696),
.Y(n_3895)
);

AOI22xp33_ASAP7_75t_L g3896 ( 
.A1(n_3777),
.A2(n_3811),
.B1(n_3791),
.B2(n_3760),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3762),
.Y(n_3897)
);

OR2x2_ASAP7_75t_L g3898 ( 
.A(n_3783),
.B(n_186),
.Y(n_3898)
);

AND2x2_ASAP7_75t_L g3899 ( 
.A(n_3818),
.B(n_187),
.Y(n_3899)
);

HB1xp67_ASAP7_75t_L g3900 ( 
.A(n_3834),
.Y(n_3900)
);

AND2x2_ASAP7_75t_L g3901 ( 
.A(n_3799),
.B(n_189),
.Y(n_3901)
);

OR2x2_ASAP7_75t_L g3902 ( 
.A(n_3767),
.B(n_189),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3800),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3810),
.B(n_190),
.Y(n_3904)
);

AND2x2_ASAP7_75t_L g3905 ( 
.A(n_3825),
.B(n_191),
.Y(n_3905)
);

NOR2xp33_ASAP7_75t_L g3906 ( 
.A(n_3762),
.B(n_191),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3827),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3801),
.B(n_192),
.Y(n_3908)
);

OR2x2_ASAP7_75t_L g3909 ( 
.A(n_3820),
.B(n_192),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3790),
.Y(n_3910)
);

AND2x2_ASAP7_75t_L g3911 ( 
.A(n_3765),
.B(n_193),
.Y(n_3911)
);

A2O1A1Ixp33_ASAP7_75t_SL g3912 ( 
.A1(n_3802),
.A2(n_193),
.B(n_194),
.C(n_195),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3813),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3839),
.Y(n_3914)
);

OR2x2_ASAP7_75t_L g3915 ( 
.A(n_3798),
.B(n_194),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3839),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3843),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3770),
.B(n_196),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3804),
.B(n_196),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3796),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3840),
.B(n_198),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3833),
.Y(n_3922)
);

AND2x2_ASAP7_75t_L g3923 ( 
.A(n_3837),
.B(n_198),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3807),
.Y(n_3924)
);

HB1xp67_ASAP7_75t_L g3925 ( 
.A(n_3834),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3814),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3814),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3847),
.B(n_199),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3775),
.Y(n_3929)
);

BUFx3_ASAP7_75t_L g3930 ( 
.A(n_3830),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3782),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3821),
.B(n_199),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3817),
.Y(n_3933)
);

OR2x2_ASAP7_75t_L g3934 ( 
.A(n_3791),
.B(n_203),
.Y(n_3934)
);

BUFx2_ASAP7_75t_L g3935 ( 
.A(n_3815),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3831),
.B(n_204),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_L g3937 ( 
.A(n_3793),
.B(n_3842),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3828),
.B(n_3784),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3841),
.B(n_205),
.Y(n_3939)
);

OAI22xp5_ASAP7_75t_L g3940 ( 
.A1(n_3838),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_3940)
);

NOR2xp33_ASAP7_75t_L g3941 ( 
.A(n_3838),
.B(n_207),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3844),
.Y(n_3942)
);

NOR2xp33_ASAP7_75t_L g3943 ( 
.A(n_3846),
.B(n_208),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_L g3944 ( 
.A(n_3853),
.B(n_3824),
.Y(n_3944)
);

AND2x2_ASAP7_75t_L g3945 ( 
.A(n_3865),
.B(n_3788),
.Y(n_3945)
);

NOR2xp67_ASAP7_75t_L g3946 ( 
.A(n_3869),
.B(n_3823),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3912),
.B(n_3822),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3874),
.Y(n_3948)
);

AND2x4_ASAP7_75t_L g3949 ( 
.A(n_3880),
.B(n_3829),
.Y(n_3949)
);

AOI22xp5_ASAP7_75t_L g3950 ( 
.A1(n_3900),
.A2(n_3850),
.B1(n_3836),
.B2(n_3826),
.Y(n_3950)
);

INVx1_ASAP7_75t_SL g3951 ( 
.A(n_3867),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3912),
.B(n_3832),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3874),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3885),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3885),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3885),
.Y(n_3956)
);

INVx2_ASAP7_75t_L g3957 ( 
.A(n_3880),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3869),
.Y(n_3958)
);

INVx2_ASAP7_75t_SL g3959 ( 
.A(n_3880),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3869),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_3880),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3889),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3889),
.Y(n_3963)
);

OAI22xp5_ASAP7_75t_L g3964 ( 
.A1(n_3896),
.A2(n_3823),
.B1(n_3848),
.B2(n_3835),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3871),
.Y(n_3965)
);

HB1xp67_ASAP7_75t_L g3966 ( 
.A(n_3858),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3857),
.Y(n_3967)
);

OAI21xp5_ASAP7_75t_SL g3968 ( 
.A1(n_3896),
.A2(n_208),
.B(n_209),
.Y(n_3968)
);

OR2x2_ASAP7_75t_L g3969 ( 
.A(n_3914),
.B(n_210),
.Y(n_3969)
);

OAI33xp33_ASAP7_75t_L g3970 ( 
.A1(n_3926),
.A2(n_211),
.A3(n_212),
.B1(n_213),
.B2(n_216),
.B3(n_217),
.Y(n_3970)
);

INVx3_ASAP7_75t_L g3971 ( 
.A(n_3851),
.Y(n_3971)
);

AOI211xp5_ASAP7_75t_L g3972 ( 
.A1(n_3900),
.A2(n_211),
.B(n_216),
.C(n_217),
.Y(n_3972)
);

INVx2_ASAP7_75t_L g3973 ( 
.A(n_3857),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3929),
.B(n_218),
.Y(n_3974)
);

OAI22xp33_ASAP7_75t_SL g3975 ( 
.A1(n_3891),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_3975)
);

XOR2x2_ASAP7_75t_L g3976 ( 
.A(n_3937),
.B(n_220),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3876),
.B(n_221),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3871),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3858),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3878),
.B(n_222),
.Y(n_3980)
);

INVx1_ASAP7_75t_SL g3981 ( 
.A(n_3935),
.Y(n_3981)
);

OAI31xp33_ASAP7_75t_L g3982 ( 
.A1(n_3925),
.A2(n_222),
.A3(n_223),
.B(n_224),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3929),
.B(n_226),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3855),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3905),
.Y(n_3985)
);

INVx1_ASAP7_75t_SL g3986 ( 
.A(n_3905),
.Y(n_3986)
);

OAI32xp33_ASAP7_75t_L g3987 ( 
.A1(n_3925),
.A2(n_226),
.A3(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_3987)
);

OA222x2_ASAP7_75t_L g3988 ( 
.A1(n_3927),
.A2(n_3930),
.B1(n_3862),
.B2(n_3913),
.C1(n_3918),
.C2(n_3934),
.Y(n_3988)
);

AND2x2_ASAP7_75t_L g3989 ( 
.A(n_3870),
.B(n_229),
.Y(n_3989)
);

XOR2x2_ASAP7_75t_L g3990 ( 
.A(n_3873),
.B(n_230),
.Y(n_3990)
);

OR2x2_ASAP7_75t_L g3991 ( 
.A(n_3916),
.B(n_230),
.Y(n_3991)
);

AND2x2_ASAP7_75t_L g3992 ( 
.A(n_3883),
.B(n_231),
.Y(n_3992)
);

AND2x2_ASAP7_75t_L g3993 ( 
.A(n_3899),
.B(n_232),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3931),
.B(n_233),
.Y(n_3994)
);

INVx2_ASAP7_75t_L g3995 ( 
.A(n_3851),
.Y(n_3995)
);

NAND2x1p5_ASAP7_75t_L g3996 ( 
.A(n_3901),
.B(n_234),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_3851),
.Y(n_3997)
);

AOI22xp5_ASAP7_75t_L g3998 ( 
.A1(n_3873),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_3931),
.B(n_236),
.Y(n_3999)
);

AND2x2_ASAP7_75t_L g4000 ( 
.A(n_3919),
.B(n_238),
.Y(n_4000)
);

AND2x2_ASAP7_75t_L g4001 ( 
.A(n_3884),
.B(n_238),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3910),
.Y(n_4002)
);

OAI22xp5_ASAP7_75t_L g4003 ( 
.A1(n_3913),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3860),
.Y(n_4004)
);

INVx1_ASAP7_75t_SL g4005 ( 
.A(n_3908),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3911),
.B(n_239),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3861),
.Y(n_4007)
);

NAND2x1_ASAP7_75t_L g4008 ( 
.A(n_3860),
.B(n_242),
.Y(n_4008)
);

AOI22xp5_ASAP7_75t_L g4009 ( 
.A1(n_3941),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_4009)
);

AOI22xp5_ASAP7_75t_L g4010 ( 
.A1(n_3941),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_4010)
);

AOI32xp33_ASAP7_75t_L g4011 ( 
.A1(n_3938),
.A2(n_248),
.A3(n_250),
.B1(n_251),
.B2(n_254),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3904),
.B(n_250),
.Y(n_4012)
);

OAI32xp33_ASAP7_75t_L g4013 ( 
.A1(n_3888),
.A2(n_254),
.A3(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_4013)
);

O2A1O1Ixp33_ASAP7_75t_L g4014 ( 
.A1(n_3863),
.A2(n_3887),
.B(n_3902),
.C(n_3866),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3923),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3875),
.Y(n_4016)
);

AOI22xp5_ASAP7_75t_L g4017 ( 
.A1(n_3940),
.A2(n_256),
.B1(n_258),
.B2(n_260),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3879),
.Y(n_4018)
);

NAND2xp33_ASAP7_75t_L g4019 ( 
.A(n_3920),
.B(n_261),
.Y(n_4019)
);

OR2x6_ASAP7_75t_L g4020 ( 
.A(n_3906),
.B(n_261),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3854),
.Y(n_4021)
);

INVx2_ASAP7_75t_L g4022 ( 
.A(n_3860),
.Y(n_4022)
);

NAND4xp75_ASAP7_75t_L g4023 ( 
.A(n_3852),
.B(n_262),
.C(n_263),
.D(n_264),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3856),
.Y(n_4024)
);

NAND2x2_ASAP7_75t_L g4025 ( 
.A(n_3930),
.B(n_3909),
.Y(n_4025)
);

INVx2_ASAP7_75t_L g4026 ( 
.A(n_3886),
.Y(n_4026)
);

NOR2x1_ASAP7_75t_L g4027 ( 
.A(n_3906),
.B(n_262),
.Y(n_4027)
);

AND2x2_ASAP7_75t_L g4028 ( 
.A(n_3932),
.B(n_263),
.Y(n_4028)
);

OAI31xp33_ASAP7_75t_L g4029 ( 
.A1(n_3887),
.A2(n_264),
.A3(n_265),
.B(n_266),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3859),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3936),
.B(n_265),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3924),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3986),
.B(n_3942),
.Y(n_4033)
);

OR2x2_ASAP7_75t_L g4034 ( 
.A(n_3951),
.B(n_3872),
.Y(n_4034)
);

NAND2xp33_ASAP7_75t_SL g4035 ( 
.A(n_4008),
.B(n_3920),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3954),
.Y(n_4036)
);

INVx2_ASAP7_75t_L g4037 ( 
.A(n_3971),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_L g4038 ( 
.A(n_3962),
.B(n_3868),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3945),
.B(n_3933),
.Y(n_4039)
);

OAI21xp5_ASAP7_75t_L g4040 ( 
.A1(n_3968),
.A2(n_3943),
.B(n_3939),
.Y(n_4040)
);

AOI21xp5_ASAP7_75t_L g4041 ( 
.A1(n_3968),
.A2(n_3947),
.B(n_4014),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3955),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3956),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3958),
.Y(n_4044)
);

AND2x2_ASAP7_75t_L g4045 ( 
.A(n_3992),
.B(n_3881),
.Y(n_4045)
);

INVx2_ASAP7_75t_L g4046 ( 
.A(n_3971),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3960),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3966),
.Y(n_4048)
);

NOR2xp33_ASAP7_75t_L g4049 ( 
.A(n_4005),
.B(n_3898),
.Y(n_4049)
);

INVx3_ASAP7_75t_L g4050 ( 
.A(n_3995),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3963),
.B(n_3922),
.Y(n_4051)
);

NOR2xp33_ASAP7_75t_L g4052 ( 
.A(n_3981),
.B(n_3921),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3989),
.B(n_3877),
.Y(n_4053)
);

CKINVDCx5p33_ASAP7_75t_R g4054 ( 
.A(n_4020),
.Y(n_4054)
);

NOR4xp25_ASAP7_75t_SL g4055 ( 
.A(n_3948),
.B(n_3903),
.C(n_3907),
.D(n_3917),
.Y(n_4055)
);

AOI22xp5_ASAP7_75t_L g4056 ( 
.A1(n_4023),
.A2(n_3864),
.B1(n_3892),
.B2(n_3893),
.Y(n_4056)
);

HB1xp67_ASAP7_75t_L g4057 ( 
.A(n_3959),
.Y(n_4057)
);

OR2x2_ASAP7_75t_L g4058 ( 
.A(n_3985),
.B(n_3915),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3965),
.Y(n_4059)
);

AND4x1_ASAP7_75t_L g4060 ( 
.A(n_4029),
.B(n_3943),
.C(n_3928),
.D(n_3894),
.Y(n_4060)
);

NOR2xp33_ASAP7_75t_L g4061 ( 
.A(n_3996),
.B(n_3864),
.Y(n_4061)
);

INVx2_ASAP7_75t_L g4062 ( 
.A(n_3997),
.Y(n_4062)
);

INVx2_ASAP7_75t_L g4063 ( 
.A(n_4004),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3978),
.Y(n_4064)
);

AND4x1_ASAP7_75t_L g4065 ( 
.A(n_4029),
.B(n_3894),
.C(n_3897),
.D(n_3890),
.Y(n_4065)
);

NOR2xp33_ASAP7_75t_R g4066 ( 
.A(n_4019),
.B(n_3886),
.Y(n_4066)
);

NOR2xp33_ASAP7_75t_L g4067 ( 
.A(n_3967),
.B(n_3890),
.Y(n_4067)
);

HB1xp67_ASAP7_75t_L g4068 ( 
.A(n_4022),
.Y(n_4068)
);

NOR2x1_ASAP7_75t_L g4069 ( 
.A(n_4027),
.B(n_3897),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_3977),
.B(n_3882),
.Y(n_4070)
);

INVx1_ASAP7_75t_SL g4071 ( 
.A(n_3949),
.Y(n_4071)
);

OR2x2_ASAP7_75t_L g4072 ( 
.A(n_3974),
.B(n_3895),
.Y(n_4072)
);

INVx2_ASAP7_75t_L g4073 ( 
.A(n_3949),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3953),
.Y(n_4074)
);

AND2x2_ASAP7_75t_L g4075 ( 
.A(n_3980),
.B(n_4001),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3979),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_L g4077 ( 
.A(n_3975),
.B(n_3882),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_L g4078 ( 
.A(n_3975),
.B(n_266),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_4015),
.B(n_267),
.Y(n_4079)
);

OR2x6_ASAP7_75t_L g4080 ( 
.A(n_3957),
.B(n_267),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3969),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3998),
.B(n_268),
.Y(n_4082)
);

INVx2_ASAP7_75t_SL g4083 ( 
.A(n_3961),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3998),
.B(n_268),
.Y(n_4084)
);

NAND2xp33_ASAP7_75t_SL g4085 ( 
.A(n_3952),
.B(n_269),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3991),
.Y(n_4086)
);

AND2x2_ASAP7_75t_L g4087 ( 
.A(n_3973),
.B(n_270),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3993),
.Y(n_4088)
);

AND2x2_ASAP7_75t_L g4089 ( 
.A(n_4000),
.B(n_271),
.Y(n_4089)
);

OR2x2_ASAP7_75t_L g4090 ( 
.A(n_3983),
.B(n_3994),
.Y(n_4090)
);

OAI21xp33_ASAP7_75t_L g4091 ( 
.A1(n_3950),
.A2(n_271),
.B(n_272),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_4011),
.B(n_273),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_4031),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_3990),
.B(n_273),
.Y(n_4094)
);

AND2x4_ASAP7_75t_L g4095 ( 
.A(n_3984),
.B(n_274),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_4028),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_4026),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_4007),
.B(n_274),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_4016),
.Y(n_4099)
);

AND2x2_ASAP7_75t_L g4100 ( 
.A(n_3988),
.B(n_275),
.Y(n_4100)
);

INVx2_ASAP7_75t_L g4101 ( 
.A(n_4020),
.Y(n_4101)
);

INVx3_ASAP7_75t_SL g4102 ( 
.A(n_4020),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_4032),
.Y(n_4103)
);

INVx2_ASAP7_75t_L g4104 ( 
.A(n_4002),
.Y(n_4104)
);

OR2x2_ASAP7_75t_L g4105 ( 
.A(n_3999),
.B(n_276),
.Y(n_4105)
);

INVx1_ASAP7_75t_SL g4106 ( 
.A(n_4012),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4018),
.Y(n_4107)
);

NOR3xp33_ASAP7_75t_L g4108 ( 
.A(n_4013),
.B(n_4021),
.C(n_3944),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_3988),
.B(n_276),
.Y(n_4109)
);

AOI21xp5_ASAP7_75t_L g4110 ( 
.A1(n_3946),
.A2(n_277),
.B(n_278),
.Y(n_4110)
);

AND2x4_ASAP7_75t_L g4111 ( 
.A(n_4024),
.B(n_277),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_4030),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_4006),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_3950),
.B(n_278),
.Y(n_4114)
);

NOR2xp33_ASAP7_75t_R g4115 ( 
.A(n_4025),
.B(n_279),
.Y(n_4115)
);

AOI22xp5_ASAP7_75t_L g4116 ( 
.A1(n_4100),
.A2(n_3976),
.B1(n_3964),
.B2(n_3946),
.Y(n_4116)
);

NOR2xp33_ASAP7_75t_L g4117 ( 
.A(n_4102),
.B(n_3970),
.Y(n_4117)
);

INVxp67_ASAP7_75t_SL g4118 ( 
.A(n_4109),
.Y(n_4118)
);

NAND2x1_ASAP7_75t_L g4119 ( 
.A(n_4050),
.B(n_4009),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_SL g4120 ( 
.A(n_4077),
.B(n_3982),
.Y(n_4120)
);

INVxp67_ASAP7_75t_L g4121 ( 
.A(n_4035),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_4071),
.B(n_3982),
.Y(n_4122)
);

OR2x2_ASAP7_75t_L g4123 ( 
.A(n_4050),
.B(n_4037),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_4068),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4046),
.Y(n_4125)
);

AND2x2_ASAP7_75t_L g4126 ( 
.A(n_4053),
.B(n_3972),
.Y(n_4126)
);

XNOR2x2_ASAP7_75t_L g4127 ( 
.A(n_4110),
.B(n_4009),
.Y(n_4127)
);

HB1xp67_ASAP7_75t_L g4128 ( 
.A(n_4069),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_4071),
.B(n_3972),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_4057),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_4080),
.Y(n_4131)
);

NAND4xp25_ASAP7_75t_L g4132 ( 
.A(n_4108),
.B(n_4010),
.C(n_4017),
.D(n_4003),
.Y(n_4132)
);

AND2x2_ASAP7_75t_L g4133 ( 
.A(n_4045),
.B(n_4075),
.Y(n_4133)
);

INVx2_ASAP7_75t_L g4134 ( 
.A(n_4080),
.Y(n_4134)
);

NAND2xp33_ASAP7_75t_SL g4135 ( 
.A(n_4055),
.B(n_4010),
.Y(n_4135)
);

OAI21xp5_ASAP7_75t_SL g4136 ( 
.A1(n_4056),
.A2(n_4017),
.B(n_3987),
.Y(n_4136)
);

INVx2_ASAP7_75t_L g4137 ( 
.A(n_4080),
.Y(n_4137)
);

OR2x2_ASAP7_75t_L g4138 ( 
.A(n_4101),
.B(n_280),
.Y(n_4138)
);

OR2x2_ASAP7_75t_L g4139 ( 
.A(n_4034),
.B(n_281),
.Y(n_4139)
);

AOI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_4041),
.A2(n_285),
.B(n_286),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_4054),
.B(n_287),
.Y(n_4141)
);

BUFx2_ASAP7_75t_L g4142 ( 
.A(n_4066),
.Y(n_4142)
);

AOI31xp33_ASAP7_75t_L g4143 ( 
.A1(n_4077),
.A2(n_288),
.A3(n_289),
.B(n_290),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_4073),
.B(n_288),
.Y(n_4144)
);

NOR2xp33_ASAP7_75t_L g4145 ( 
.A(n_4083),
.B(n_289),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_4062),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_SL g4147 ( 
.A(n_4065),
.B(n_290),
.Y(n_4147)
);

AND2x2_ASAP7_75t_L g4148 ( 
.A(n_4039),
.B(n_291),
.Y(n_4148)
);

AND2x2_ASAP7_75t_L g4149 ( 
.A(n_4070),
.B(n_291),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_L g4150 ( 
.A(n_4063),
.B(n_292),
.Y(n_4150)
);

OR2x2_ASAP7_75t_L g4151 ( 
.A(n_4033),
.B(n_292),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_4048),
.B(n_4041),
.Y(n_4152)
);

OAI22xp5_ASAP7_75t_L g4153 ( 
.A1(n_4061),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_4153)
);

NAND3xp33_ASAP7_75t_L g4154 ( 
.A(n_4060),
.B(n_294),
.C(n_295),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_4096),
.B(n_296),
.Y(n_4155)
);

HB1xp67_ASAP7_75t_L g4156 ( 
.A(n_4110),
.Y(n_4156)
);

NOR2xp33_ASAP7_75t_L g4157 ( 
.A(n_4078),
.B(n_297),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_4089),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_4088),
.B(n_298),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_4036),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_4042),
.Y(n_4161)
);

OAI21xp5_ASAP7_75t_L g4162 ( 
.A1(n_4114),
.A2(n_299),
.B(n_300),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4043),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_4079),
.B(n_4087),
.Y(n_4164)
);

AND2x4_ASAP7_75t_L g4165 ( 
.A(n_4081),
.B(n_299),
.Y(n_4165)
);

NOR2xp33_ASAP7_75t_L g4166 ( 
.A(n_4078),
.B(n_300),
.Y(n_4166)
);

AND2x2_ASAP7_75t_L g4167 ( 
.A(n_4049),
.B(n_301),
.Y(n_4167)
);

INVx2_ASAP7_75t_SL g4168 ( 
.A(n_4095),
.Y(n_4168)
);

NOR2xp33_ASAP7_75t_L g4169 ( 
.A(n_4033),
.B(n_301),
.Y(n_4169)
);

NAND2x1_ASAP7_75t_L g4170 ( 
.A(n_4095),
.B(n_302),
.Y(n_4170)
);

INVx2_ASAP7_75t_L g4171 ( 
.A(n_4058),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_4086),
.B(n_302),
.Y(n_4172)
);

INVx2_ASAP7_75t_L g4173 ( 
.A(n_4111),
.Y(n_4173)
);

AND2x2_ASAP7_75t_L g4174 ( 
.A(n_4106),
.B(n_303),
.Y(n_4174)
);

INVx3_ASAP7_75t_L g4175 ( 
.A(n_4111),
.Y(n_4175)
);

INVx1_ASAP7_75t_SL g4176 ( 
.A(n_4115),
.Y(n_4176)
);

NOR2x1_ASAP7_75t_L g4177 ( 
.A(n_4114),
.B(n_303),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4038),
.Y(n_4178)
);

INVx2_ASAP7_75t_L g4179 ( 
.A(n_4105),
.Y(n_4179)
);

INVx2_ASAP7_75t_L g4180 ( 
.A(n_4090),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4175),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_4128),
.Y(n_4182)
);

AOI21xp5_ASAP7_75t_L g4183 ( 
.A1(n_4135),
.A2(n_4040),
.B(n_4085),
.Y(n_4183)
);

INVxp67_ASAP7_75t_L g4184 ( 
.A(n_4118),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4128),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_4123),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_4133),
.B(n_4106),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_4118),
.B(n_4052),
.Y(n_4188)
);

AOI322xp5_ASAP7_75t_L g4189 ( 
.A1(n_4135),
.A2(n_4091),
.A3(n_4076),
.B1(n_4092),
.B2(n_4094),
.C1(n_4038),
.C2(n_4074),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4175),
.Y(n_4190)
);

AND2x2_ASAP7_75t_L g4191 ( 
.A(n_4176),
.B(n_4040),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_4134),
.Y(n_4192)
);

A2O1A1Ixp33_ASAP7_75t_L g4193 ( 
.A1(n_4140),
.A2(n_4082),
.B(n_4084),
.C(n_4092),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_4170),
.Y(n_4194)
);

AOI21xp5_ASAP7_75t_L g4195 ( 
.A1(n_4147),
.A2(n_4082),
.B(n_4084),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4137),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_4126),
.B(n_4093),
.Y(n_4197)
);

INVx1_ASAP7_75t_SL g4198 ( 
.A(n_4142),
.Y(n_4198)
);

NOR2xp33_ASAP7_75t_L g4199 ( 
.A(n_4120),
.B(n_4094),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_4148),
.B(n_4113),
.Y(n_4200)
);

OAI22xp5_ASAP7_75t_L g4201 ( 
.A1(n_4116),
.A2(n_4098),
.B1(n_4072),
.B2(n_4051),
.Y(n_4201)
);

NAND2x1_ASAP7_75t_L g4202 ( 
.A(n_4168),
.B(n_4059),
.Y(n_4202)
);

OAI22xp5_ASAP7_75t_SL g4203 ( 
.A1(n_4119),
.A2(n_4051),
.B1(n_4067),
.B2(n_4104),
.Y(n_4203)
);

AOI22xp5_ASAP7_75t_L g4204 ( 
.A1(n_4120),
.A2(n_4107),
.B1(n_4103),
.B2(n_4099),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_4156),
.B(n_4097),
.Y(n_4205)
);

AOI22xp33_ASAP7_75t_L g4206 ( 
.A1(n_4132),
.A2(n_4112),
.B1(n_4047),
.B2(n_4044),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_4131),
.Y(n_4207)
);

AND2x2_ASAP7_75t_L g4208 ( 
.A(n_4171),
.B(n_4064),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_4121),
.B(n_4098),
.Y(n_4209)
);

OAI221xp5_ASAP7_75t_L g4210 ( 
.A1(n_4136),
.A2(n_4147),
.B1(n_4152),
.B2(n_4154),
.C(n_4140),
.Y(n_4210)
);

AND2x4_ASAP7_75t_L g4211 ( 
.A(n_4121),
.B(n_304),
.Y(n_4211)
);

HB1xp67_ASAP7_75t_L g4212 ( 
.A(n_4156),
.Y(n_4212)
);

AND2x2_ASAP7_75t_L g4213 ( 
.A(n_4158),
.B(n_4130),
.Y(n_4213)
);

AND2x2_ASAP7_75t_L g4214 ( 
.A(n_4149),
.B(n_304),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_4173),
.Y(n_4215)
);

OR2x2_ASAP7_75t_L g4216 ( 
.A(n_4122),
.B(n_306),
.Y(n_4216)
);

AOI221xp5_ASAP7_75t_L g4217 ( 
.A1(n_4117),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.C(n_309),
.Y(n_4217)
);

AND2x2_ASAP7_75t_L g4218 ( 
.A(n_4167),
.B(n_308),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4124),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4139),
.Y(n_4220)
);

AOI222xp33_ASAP7_75t_SL g4221 ( 
.A1(n_4178),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.C1(n_313),
.C2(n_314),
.Y(n_4221)
);

INVx1_ASAP7_75t_SL g4222 ( 
.A(n_4129),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_4117),
.B(n_310),
.Y(n_4223)
);

OAI22xp33_ASAP7_75t_L g4224 ( 
.A1(n_4143),
.A2(n_311),
.B1(n_312),
.B2(n_314),
.Y(n_4224)
);

AOI22xp33_ASAP7_75t_L g4225 ( 
.A1(n_4127),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_4225)
);

NAND2xp33_ASAP7_75t_L g4226 ( 
.A(n_4177),
.B(n_315),
.Y(n_4226)
);

AND2x2_ASAP7_75t_L g4227 ( 
.A(n_4159),
.B(n_316),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_4145),
.B(n_318),
.Y(n_4228)
);

O2A1O1Ixp33_ASAP7_75t_SL g4229 ( 
.A1(n_4164),
.A2(n_4141),
.B(n_4151),
.C(n_4160),
.Y(n_4229)
);

A2O1A1Ixp33_ASAP7_75t_L g4230 ( 
.A1(n_4169),
.A2(n_318),
.B(n_319),
.C(n_320),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4174),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_4145),
.B(n_320),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_4138),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_L g4234 ( 
.A(n_4157),
.B(n_321),
.Y(n_4234)
);

OAI21xp33_ASAP7_75t_L g4235 ( 
.A1(n_4125),
.A2(n_321),
.B(n_324),
.Y(n_4235)
);

OAI21xp33_ASAP7_75t_L g4236 ( 
.A1(n_4146),
.A2(n_325),
.B(n_326),
.Y(n_4236)
);

NAND3xp33_ASAP7_75t_L g4237 ( 
.A(n_4169),
.B(n_325),
.C(n_327),
.Y(n_4237)
);

INVxp67_ASAP7_75t_L g4238 ( 
.A(n_4157),
.Y(n_4238)
);

AOI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_4166),
.A2(n_327),
.B(n_328),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_4166),
.B(n_328),
.Y(n_4240)
);

O2A1O1Ixp33_ASAP7_75t_L g4241 ( 
.A1(n_4153),
.A2(n_329),
.B(n_330),
.C(n_332),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_4187),
.B(n_4180),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_4184),
.B(n_4180),
.Y(n_4243)
);

AND2x2_ASAP7_75t_L g4244 ( 
.A(n_4191),
.B(n_4179),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_4181),
.B(n_4161),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4212),
.Y(n_4246)
);

OAI22xp33_ASAP7_75t_L g4247 ( 
.A1(n_4183),
.A2(n_4144),
.B1(n_4155),
.B2(n_4172),
.Y(n_4247)
);

AOI21xp5_ASAP7_75t_L g4248 ( 
.A1(n_4188),
.A2(n_4162),
.B(n_4150),
.Y(n_4248)
);

XOR2x2_ASAP7_75t_L g4249 ( 
.A(n_4199),
.B(n_4163),
.Y(n_4249)
);

AOI21xp33_ASAP7_75t_L g4250 ( 
.A1(n_4202),
.A2(n_4165),
.B(n_330),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4190),
.Y(n_4251)
);

OR2x2_ASAP7_75t_L g4252 ( 
.A(n_4188),
.B(n_4165),
.Y(n_4252)
);

OAI22xp5_ASAP7_75t_L g4253 ( 
.A1(n_4225),
.A2(n_329),
.B1(n_337),
.B2(n_338),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4226),
.Y(n_4254)
);

AOI32xp33_ASAP7_75t_L g4255 ( 
.A1(n_4198),
.A2(n_338),
.A3(n_339),
.B1(n_340),
.B2(n_342),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4211),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_SL g4257 ( 
.A(n_4194),
.B(n_339),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_4211),
.B(n_340),
.Y(n_4258)
);

OR2x2_ASAP7_75t_L g4259 ( 
.A(n_4215),
.B(n_342),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_4189),
.B(n_344),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_L g4261 ( 
.A(n_4222),
.B(n_345),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_4214),
.B(n_345),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4205),
.Y(n_4263)
);

AOI21xp33_ASAP7_75t_L g4264 ( 
.A1(n_4223),
.A2(n_346),
.B(n_347),
.Y(n_4264)
);

INVx2_ASAP7_75t_L g4265 ( 
.A(n_4218),
.Y(n_4265)
);

NAND2x1_ASAP7_75t_L g4266 ( 
.A(n_4182),
.B(n_346),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4205),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_4227),
.B(n_347),
.Y(n_4268)
);

AOI21xp33_ASAP7_75t_L g4269 ( 
.A1(n_4223),
.A2(n_348),
.B(n_349),
.Y(n_4269)
);

NOR2xp33_ASAP7_75t_L g4270 ( 
.A(n_4210),
.B(n_350),
.Y(n_4270)
);

AOI211xp5_ASAP7_75t_L g4271 ( 
.A1(n_4203),
.A2(n_351),
.B(n_353),
.C(n_354),
.Y(n_4271)
);

NAND4xp25_ASAP7_75t_SL g4272 ( 
.A(n_4206),
.B(n_351),
.C(n_353),
.D(n_354),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4213),
.Y(n_4273)
);

XNOR2xp5_ASAP7_75t_L g4274 ( 
.A(n_4197),
.B(n_355),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_SL g4275 ( 
.A(n_4224),
.B(n_4204),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4185),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_4186),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_4192),
.B(n_355),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4209),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4196),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4208),
.Y(n_4281)
);

XNOR2xp5_ASAP7_75t_L g4282 ( 
.A(n_4201),
.B(n_356),
.Y(n_4282)
);

INVx1_ASAP7_75t_SL g4283 ( 
.A(n_4216),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4200),
.Y(n_4284)
);

NAND4xp25_ASAP7_75t_L g4285 ( 
.A(n_4193),
.B(n_356),
.C(n_357),
.D(n_359),
.Y(n_4285)
);

XOR2xp5_ASAP7_75t_L g4286 ( 
.A(n_4201),
.B(n_357),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4231),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_4195),
.B(n_359),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_4207),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_4220),
.B(n_4239),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4228),
.Y(n_4291)
);

OR2x2_ASAP7_75t_L g4292 ( 
.A(n_4256),
.B(n_4219),
.Y(n_4292)
);

BUFx2_ASAP7_75t_L g4293 ( 
.A(n_4242),
.Y(n_4293)
);

XOR2x2_ASAP7_75t_L g4294 ( 
.A(n_4249),
.B(n_4274),
.Y(n_4294)
);

NOR2xp33_ASAP7_75t_L g4295 ( 
.A(n_4285),
.B(n_4235),
.Y(n_4295)
);

OR2x2_ASAP7_75t_L g4296 ( 
.A(n_4252),
.B(n_4233),
.Y(n_4296)
);

NOR2xp33_ASAP7_75t_L g4297 ( 
.A(n_4285),
.B(n_4236),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_L g4298 ( 
.A(n_4271),
.B(n_4238),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4266),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4244),
.Y(n_4300)
);

NOR3xp33_ASAP7_75t_SL g4301 ( 
.A(n_4275),
.B(n_4217),
.C(n_4237),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4258),
.Y(n_4302)
);

AOI221xp5_ASAP7_75t_L g4303 ( 
.A1(n_4286),
.A2(n_4229),
.B1(n_4241),
.B2(n_4234),
.C(n_4240),
.Y(n_4303)
);

INVx2_ASAP7_75t_SL g4304 ( 
.A(n_4246),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4243),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4259),
.Y(n_4306)
);

HB1xp67_ASAP7_75t_L g4307 ( 
.A(n_4282),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4284),
.Y(n_4308)
);

NAND2xp33_ASAP7_75t_SL g4309 ( 
.A(n_4254),
.B(n_4232),
.Y(n_4309)
);

INVx1_ASAP7_75t_SL g4310 ( 
.A(n_4283),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4271),
.B(n_4230),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_4273),
.B(n_4240),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_4255),
.B(n_4234),
.Y(n_4313)
);

AND2x2_ASAP7_75t_L g4314 ( 
.A(n_4265),
.B(n_4281),
.Y(n_4314)
);

INVxp67_ASAP7_75t_L g4315 ( 
.A(n_4270),
.Y(n_4315)
);

XOR2xp5_ASAP7_75t_L g4316 ( 
.A(n_4272),
.B(n_4221),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_SL g4317 ( 
.A(n_4250),
.B(n_4221),
.Y(n_4317)
);

AOI21xp33_ASAP7_75t_L g4318 ( 
.A1(n_4260),
.A2(n_360),
.B(n_361),
.Y(n_4318)
);

INVx2_ASAP7_75t_L g4319 ( 
.A(n_4277),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_L g4320 ( 
.A(n_4251),
.B(n_361),
.Y(n_4320)
);

CKINVDCx20_ASAP7_75t_R g4321 ( 
.A(n_4283),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_4253),
.B(n_362),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4262),
.Y(n_4323)
);

OAI21xp5_ASAP7_75t_L g4324 ( 
.A1(n_4288),
.A2(n_362),
.B(n_363),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_4253),
.B(n_364),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4261),
.Y(n_4326)
);

INVx2_ASAP7_75t_SL g4327 ( 
.A(n_4276),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_4280),
.B(n_4289),
.Y(n_4328)
);

NOR2x1_ASAP7_75t_L g4329 ( 
.A(n_4257),
.B(n_4263),
.Y(n_4329)
);

A2O1A1Ixp33_ASAP7_75t_L g4330 ( 
.A1(n_4295),
.A2(n_4267),
.B(n_4248),
.C(n_4287),
.Y(n_4330)
);

AOI21xp33_ASAP7_75t_SL g4331 ( 
.A1(n_4299),
.A2(n_4247),
.B(n_4290),
.Y(n_4331)
);

NOR2xp33_ASAP7_75t_SL g4332 ( 
.A(n_4293),
.B(n_4269),
.Y(n_4332)
);

NOR2xp67_ASAP7_75t_L g4333 ( 
.A(n_4304),
.B(n_4268),
.Y(n_4333)
);

AOI221xp5_ASAP7_75t_L g4334 ( 
.A1(n_4318),
.A2(n_4245),
.B1(n_4279),
.B2(n_4291),
.C(n_4278),
.Y(n_4334)
);

AOI22xp5_ASAP7_75t_L g4335 ( 
.A1(n_4321),
.A2(n_4264),
.B1(n_366),
.B2(n_367),
.Y(n_4335)
);

INVxp33_ASAP7_75t_SL g4336 ( 
.A(n_4316),
.Y(n_4336)
);

NAND2xp33_ASAP7_75t_SL g4337 ( 
.A(n_4301),
.B(n_364),
.Y(n_4337)
);

OAI21x1_ASAP7_75t_SL g4338 ( 
.A1(n_4324),
.A2(n_366),
.B(n_367),
.Y(n_4338)
);

NAND2xp33_ASAP7_75t_L g4339 ( 
.A(n_4310),
.B(n_368),
.Y(n_4339)
);

OAI211xp5_ASAP7_75t_SL g4340 ( 
.A1(n_4303),
.A2(n_369),
.B(n_978),
.C(n_1072),
.Y(n_4340)
);

OA22x2_ASAP7_75t_L g4341 ( 
.A1(n_4310),
.A2(n_369),
.B1(n_1072),
.B2(n_1062),
.Y(n_4341)
);

INVxp67_ASAP7_75t_L g4342 ( 
.A(n_4297),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4292),
.Y(n_4343)
);

NOR3xp33_ASAP7_75t_L g4344 ( 
.A(n_4309),
.B(n_1072),
.C(n_1062),
.Y(n_4344)
);

INVx2_ASAP7_75t_SL g4345 ( 
.A(n_4296),
.Y(n_4345)
);

AOI221xp5_ASAP7_75t_L g4346 ( 
.A1(n_4318),
.A2(n_1071),
.B1(n_1070),
.B2(n_1062),
.C(n_1072),
.Y(n_4346)
);

AOI22xp5_ASAP7_75t_L g4347 ( 
.A1(n_4300),
.A2(n_4314),
.B1(n_4317),
.B2(n_4294),
.Y(n_4347)
);

INVx1_ASAP7_75t_SL g4348 ( 
.A(n_4298),
.Y(n_4348)
);

AOI22xp5_ASAP7_75t_L g4349 ( 
.A1(n_4305),
.A2(n_1072),
.B1(n_1009),
.B2(n_1062),
.Y(n_4349)
);

NOR2x1_ASAP7_75t_L g4350 ( 
.A(n_4329),
.B(n_1071),
.Y(n_4350)
);

NOR3xp33_ASAP7_75t_L g4351 ( 
.A(n_4312),
.B(n_1062),
.C(n_1070),
.Y(n_4351)
);

AOI21xp5_ASAP7_75t_L g4352 ( 
.A1(n_4313),
.A2(n_1070),
.B(n_1071),
.Y(n_4352)
);

OAI21xp5_ASAP7_75t_L g4353 ( 
.A1(n_4308),
.A2(n_988),
.B(n_979),
.Y(n_4353)
);

AOI22xp33_ASAP7_75t_L g4354 ( 
.A1(n_4336),
.A2(n_4319),
.B1(n_4327),
.B2(n_4307),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_4345),
.Y(n_4355)
);

NOR2xp33_ASAP7_75t_L g4356 ( 
.A(n_4332),
.B(n_4311),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4339),
.Y(n_4357)
);

BUFx12f_ASAP7_75t_L g4358 ( 
.A(n_4348),
.Y(n_4358)
);

NOR2x1_ASAP7_75t_L g4359 ( 
.A(n_4343),
.B(n_4333),
.Y(n_4359)
);

NOR2xp33_ASAP7_75t_L g4360 ( 
.A(n_4331),
.B(n_4306),
.Y(n_4360)
);

A2O1A1Ixp33_ASAP7_75t_L g4361 ( 
.A1(n_4337),
.A2(n_4324),
.B(n_4322),
.C(n_4325),
.Y(n_4361)
);

AOI21xp5_ASAP7_75t_L g4362 ( 
.A1(n_4330),
.A2(n_4328),
.B(n_4320),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4338),
.Y(n_4363)
);

NAND2xp5_ASAP7_75t_L g4364 ( 
.A(n_4347),
.B(n_4320),
.Y(n_4364)
);

OAI22xp5_ASAP7_75t_L g4365 ( 
.A1(n_4335),
.A2(n_4315),
.B1(n_4326),
.B2(n_4302),
.Y(n_4365)
);

OAI221xp5_ASAP7_75t_L g4366 ( 
.A1(n_4342),
.A2(n_4323),
.B1(n_978),
.B2(n_1071),
.C(n_1070),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4341),
.Y(n_4367)
);

OAI22xp5_ASAP7_75t_SL g4368 ( 
.A1(n_4350),
.A2(n_1071),
.B1(n_1122),
.B2(n_957),
.Y(n_4368)
);

OAI21xp33_ASAP7_75t_L g4369 ( 
.A1(n_4334),
.A2(n_1122),
.B(n_955),
.Y(n_4369)
);

NOR2xp33_ASAP7_75t_L g4370 ( 
.A(n_4355),
.B(n_4358),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_SL g4371 ( 
.A(n_4359),
.B(n_4346),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4360),
.Y(n_4372)
);

OA22x2_ASAP7_75t_L g4373 ( 
.A1(n_4363),
.A2(n_4357),
.B1(n_4367),
.B2(n_4364),
.Y(n_4373)
);

AOI22xp5_ASAP7_75t_L g4374 ( 
.A1(n_4356),
.A2(n_4340),
.B1(n_4344),
.B2(n_4351),
.Y(n_4374)
);

NOR2x1_ASAP7_75t_L g4375 ( 
.A(n_4362),
.B(n_4361),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4365),
.Y(n_4376)
);

AO22x1_ASAP7_75t_L g4377 ( 
.A1(n_4354),
.A2(n_4353),
.B1(n_4352),
.B2(n_4349),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4369),
.Y(n_4378)
);

AOI22xp5_ASAP7_75t_L g4379 ( 
.A1(n_4368),
.A2(n_1122),
.B1(n_955),
.B2(n_957),
.Y(n_4379)
);

NOR2x1_ASAP7_75t_L g4380 ( 
.A(n_4366),
.B(n_1122),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4370),
.B(n_955),
.Y(n_4381)
);

AOI22xp5_ASAP7_75t_L g4382 ( 
.A1(n_4372),
.A2(n_955),
.B1(n_957),
.B2(n_1289),
.Y(n_4382)
);

AOI221xp5_ASAP7_75t_L g4383 ( 
.A1(n_4376),
.A2(n_4377),
.B1(n_4378),
.B2(n_4371),
.C(n_4374),
.Y(n_4383)
);

HB1xp67_ASAP7_75t_L g4384 ( 
.A(n_4375),
.Y(n_4384)
);

AO22x1_ASAP7_75t_SL g4385 ( 
.A1(n_4373),
.A2(n_955),
.B1(n_957),
.B2(n_1289),
.Y(n_4385)
);

NOR2xp67_ASAP7_75t_L g4386 ( 
.A(n_4379),
.B(n_988),
.Y(n_4386)
);

NOR2x1_ASAP7_75t_L g4387 ( 
.A(n_4381),
.B(n_4380),
.Y(n_4387)
);

NOR2x1_ASAP7_75t_L g4388 ( 
.A(n_4386),
.B(n_957),
.Y(n_4388)
);

AND2x4_ASAP7_75t_L g4389 ( 
.A(n_4384),
.B(n_957),
.Y(n_4389)
);

INVx1_ASAP7_75t_L g4390 ( 
.A(n_4385),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4383),
.Y(n_4391)
);

OAI221xp5_ASAP7_75t_L g4392 ( 
.A1(n_4391),
.A2(n_4382),
.B1(n_1289),
.B2(n_1218),
.C(n_1202),
.Y(n_4392)
);

OAI211xp5_ASAP7_75t_L g4393 ( 
.A1(n_4390),
.A2(n_1289),
.B(n_1218),
.C(n_1202),
.Y(n_4393)
);

NAND4xp75_ASAP7_75t_L g4394 ( 
.A(n_4393),
.B(n_4387),
.C(n_4388),
.D(n_4389),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4392),
.Y(n_4395)
);

NAND3xp33_ASAP7_75t_L g4396 ( 
.A(n_4395),
.B(n_1289),
.C(n_1218),
.Y(n_4396)
);

OR3x1_ASAP7_75t_L g4397 ( 
.A(n_4396),
.B(n_4394),
.C(n_1218),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4397),
.Y(n_4398)
);

OAI21xp5_ASAP7_75t_L g4399 ( 
.A1(n_4398),
.A2(n_988),
.B(n_979),
.Y(n_4399)
);

BUFx4f_ASAP7_75t_SL g4400 ( 
.A(n_4399),
.Y(n_4400)
);

OAI22xp5_ASAP7_75t_L g4401 ( 
.A1(n_4400),
.A2(n_1202),
.B1(n_1218),
.B2(n_988),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4401),
.Y(n_4402)
);

XNOR2x1_ASAP7_75t_L g4403 ( 
.A(n_4402),
.B(n_996),
.Y(n_4403)
);

AOI22xp33_ASAP7_75t_R g4404 ( 
.A1(n_4403),
.A2(n_988),
.B1(n_979),
.B2(n_954),
.Y(n_4404)
);

AOI322xp5_ASAP7_75t_L g4405 ( 
.A1(n_4403),
.A2(n_954),
.A3(n_979),
.B1(n_988),
.B2(n_996),
.C1(n_1024),
.C2(n_4310),
.Y(n_4405)
);

OAI22xp5_ASAP7_75t_L g4406 ( 
.A1(n_4404),
.A2(n_954),
.B1(n_979),
.B2(n_996),
.Y(n_4406)
);

AOI221xp5_ASAP7_75t_L g4407 ( 
.A1(n_4406),
.A2(n_4405),
.B1(n_979),
.B2(n_954),
.C(n_1024),
.Y(n_4407)
);

AOI211xp5_ASAP7_75t_L g4408 ( 
.A1(n_4407),
.A2(n_1024),
.B(n_996),
.C(n_954),
.Y(n_4408)
);


endmodule