module fake_jpeg_23466_n_37 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_37);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_32;

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_26),
.B1(n_6),
.B2(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx24_ASAP7_75t_SL g30 ( 
.A(n_25),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_18),
.B1(n_7),
.B2(n_9),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_29),
.Y(n_32)
);

AOI22x1_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_16),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_32),
.Y(n_35)
);

BUFx24_ASAP7_75t_SL g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_27),
.Y(n_37)
);


endmodule