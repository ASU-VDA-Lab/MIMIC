module fake_jpeg_8520_n_55 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_55);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_55;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_8),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_12),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_10),
.B1(n_20),
.B2(n_18),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_0),
.Y(n_37)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_22),
.B(n_1),
.C(n_2),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_40),
.B(n_7),
.C(n_11),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_42),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_1),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_45),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_3),
.B(n_6),
.Y(n_45)
);

OA21x2_ASAP7_75t_SL g50 ( 
.A1(n_49),
.A2(n_40),
.B(n_37),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B1(n_39),
.B2(n_46),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_38),
.C(n_41),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_49),
.B1(n_47),
.B2(n_43),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_21),
.B(n_13),
.Y(n_55)
);


endmodule