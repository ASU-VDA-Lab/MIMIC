module fake_jpeg_28982_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_SL g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_7),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_74),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_81),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_79),
.Y(n_96)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_82),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_72),
.B1(n_64),
.B2(n_66),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_67),
.B1(n_52),
.B2(n_62),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_73),
.C(n_51),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_92),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_31),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_50),
.B1(n_71),
.B2(n_68),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_50),
.B1(n_71),
.B2(n_68),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_93),
.B1(n_57),
.B2(n_53),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_69),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_66),
.B1(n_56),
.B2(n_70),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_133)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_3),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_104),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_60),
.B(n_58),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_9),
.C(n_10),
.Y(n_130)
);

NOR2x1p5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_57),
.Y(n_107)
);

AO22x1_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_57),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_110),
.B(n_3),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_135)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_0),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_8),
.B(n_9),
.Y(n_129)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_105),
.B(n_61),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_120),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_96),
.B1(n_97),
.B2(n_2),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_130),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_5),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_133),
.Y(n_151)
);

AO22x1_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_111),
.B(n_116),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_141),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_146),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_106),
.C(n_102),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_141),
.C(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_24),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_148),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_26),
.B(n_27),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_153),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_38),
.C(n_40),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_35),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_149),
.B(n_152),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_144),
.C(n_151),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_137),
.B1(n_127),
.B2(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_159),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_158),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_156),
.C(n_160),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_165),
.B1(n_160),
.B2(n_162),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_142),
.B1(n_140),
.B2(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_154),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_138),
.B(n_43),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_42),
.B(n_44),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_46),
.C(n_47),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_48),
.Y(n_172)
);


endmodule