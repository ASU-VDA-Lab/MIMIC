module fake_jpeg_2674_n_107 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_10),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_34),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

CKINVDCx11_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_32),
.Y(n_37)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_12),
.B(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_8),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_27),
.B(n_30),
.C(n_32),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_35),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_15),
.B1(n_21),
.B2(n_18),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_47),
.B1(n_24),
.B2(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_17),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_28),
.A2(n_21),
.B1(n_18),
.B2(n_15),
.Y(n_47)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_1),
.C(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_29),
.A2(n_24),
.B1(n_22),
.B2(n_14),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_25),
.B1(n_17),
.B2(n_19),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_54),
.B1(n_59),
.B2(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_63),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_61),
.Y(n_65)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_25),
.B1(n_35),
.B2(n_20),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_25),
.B1(n_35),
.B2(n_3),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_55),
.B1(n_57),
.B2(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_9),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_2),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_48),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_74),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_46),
.B1(n_52),
.B2(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_77),
.C(n_76),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_51),
.C(n_55),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_67),
.C(n_66),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_71),
.B(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_82),
.Y(n_87)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_81),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_72),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_82),
.C(n_62),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_75),
.B1(n_73),
.B2(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_90),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_93),
.B1(n_64),
.B2(n_44),
.Y(n_98)
);

OAI321xp33_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_78),
.A3(n_83),
.B1(n_81),
.B2(n_64),
.C(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_86),
.C(n_85),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_94),
.C(n_44),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_99),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_41),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_100),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_104),
.A3(n_100),
.B1(n_58),
.B2(n_42),
.C1(n_9),
.C2(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_97),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_39),
.C(n_2),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_58),
.Y(n_107)
);


endmodule