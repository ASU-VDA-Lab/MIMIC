module fake_jpeg_1083_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_5),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_8),
.B(n_1),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_20),
.B(n_22),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_7),
.A2(n_10),
.B1(n_14),
.B2(n_12),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_11),
.B1(n_0),
.B2(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_11),
.B1(n_14),
.B2(n_3),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_0),
.B(n_4),
.Y(n_29)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_21),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_19),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_29),
.Y(n_30)
);

AOI21x1_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_18),
.B(n_17),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_20),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_18),
.B1(n_17),
.B2(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_16),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_28),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_29),
.B(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_37),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_34),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_32),
.C(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_41),
.B(n_39),
.Y(n_42)
);

AOI322xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_43),
.A3(n_22),
.B1(n_24),
.B2(n_31),
.C1(n_40),
.C2(n_35),
.Y(n_44)
);

NOR3xp33_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_42),
.C(n_22),
.Y(n_45)
);


endmodule