module fake_netlist_6_3656_n_1204 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1204);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1204;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_881;
wire n_1199;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_1189;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_1033;
wire n_671;
wire n_726;
wire n_607;
wire n_1052;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_1203;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_1164;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_180;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_898;
wire n_617;
wire n_698;
wire n_233;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_284;
wire n_955;
wire n_337;
wire n_865;
wire n_1138;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1099;
wire n_1101;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_1192;
wire n_421;
wire n_781;
wire n_789;
wire n_424;
wire n_615;
wire n_1130;
wire n_181;
wire n_1127;
wire n_182;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_1187;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_1139;
wire n_198;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_718;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_1078;
wire n_923;
wire n_504;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_1196;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_720;
wire n_758;
wire n_516;
wire n_842;
wire n_525;
wire n_1163;
wire n_1173;
wire n_1180;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_772;
wire n_656;
wire n_843;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_886;
wire n_343;
wire n_953;
wire n_448;
wire n_1094;
wire n_1017;
wire n_1004;
wire n_1176;
wire n_1190;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_930;
wire n_684;
wire n_425;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_1181;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_236;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_1084;
wire n_929;
wire n_460;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_870;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_1152;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_185;
wire n_712;
wire n_1183;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1193;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_228;
wire n_1195;
wire n_356;
wire n_577;
wire n_936;
wire n_184;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_1201;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_1075;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_1198;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_689;
wire n_354;
wire n_231;
wire n_799;
wire n_505;
wire n_240;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_1194;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_249;
wire n_386;
wire n_201;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_199;
wire n_1167;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_1153;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_1185;
wire n_453;
wire n_612;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_1175;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_1188;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_288;
wire n_427;
wire n_1200;
wire n_1059;
wire n_1197;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1154;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1177;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_1191;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_1007;
wire n_649;
wire n_855;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_40),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_43),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_70),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_22),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_87),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_69),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_90),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_88),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_55),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_93),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_86),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_46),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_37),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_5),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_29),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_57),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_172),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_101),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_135),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_39),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_115),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_107),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_111),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_10),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_6),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_112),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_0),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_158),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_38),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_32),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_31),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_26),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_50),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_124),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_14),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_64),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_139),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_104),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_118),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_96),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_95),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_120),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_48),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_21),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_129),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_105),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_82),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_8),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_100),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_61),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_161),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_77),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_28),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_179),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_186),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_182),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_180),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_182),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_181),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_185),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_188),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_189),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_191),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_195),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_196),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_198),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_202),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_203),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_207),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_209),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_221),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_210),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_215),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_237),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_242),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_238),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_241),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_247),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_241),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_250),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_252),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_254),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_255),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_243),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_258),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_243),
.B(n_187),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_259),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_260),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_261),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_266),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_239),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_264),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_264),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_239),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_239),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_239),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_239),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_241),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_253),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_237),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_237),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_237),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_248),
.Y(n_310)
);

BUFx8_ASAP7_75t_SL g311 ( 
.A(n_241),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_248),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_237),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_253),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_253),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_275),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_280),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_287),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_311),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_267),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_269),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_300),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_275),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_300),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_306),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_314),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_315),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_272),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_291),
.Y(n_336)
);

INVxp33_ASAP7_75t_SL g337 ( 
.A(n_313),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_282),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_312),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_305),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_268),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_300),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_304),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_272),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_270),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_300),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_277),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_297),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_278),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_271),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_286),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_303),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_303),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_285),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_321),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_335),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_317),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_321),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_318),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_320),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_340),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_293),
.Y(n_370)
);

NOR2xp67_ASAP7_75t_L g371 ( 
.A(n_359),
.B(n_296),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_360),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_319),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_343),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_343),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_335),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_322),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_354),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_274),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_354),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_274),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_346),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_346),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_323),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_290),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_325),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_320),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_330),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_361),
.B(n_281),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_350),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_350),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_347),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_347),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_331),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_326),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_362),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_352),
.B(n_290),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_316),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_332),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_337),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_337),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_283),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_328),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_351),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_329),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_392),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_406),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_364),
.A2(n_277),
.B1(n_288),
.B2(n_336),
.Y(n_409)
);

OAI22x1_ASAP7_75t_SL g410 ( 
.A1(n_390),
.A2(n_217),
.B1(n_288),
.B2(n_294),
.Y(n_410)
);

OA21x2_ASAP7_75t_L g411 ( 
.A1(n_399),
.A2(n_345),
.B(n_349),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_399),
.Y(n_412)
);

AOI22x1_ASAP7_75t_SL g413 ( 
.A1(n_364),
.A2(n_217),
.B1(n_187),
.B2(n_219),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_393),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_394),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_406),
.Y(n_416)
);

NOR2x1_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_353),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_393),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_396),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_404),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_365),
.B(n_333),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_372),
.B(n_360),
.Y(n_422)
);

OA21x2_ASAP7_75t_L g423 ( 
.A1(n_367),
.A2(n_344),
.B(n_327),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_373),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

AOI22x1_ASAP7_75t_SL g426 ( 
.A1(n_383),
.A2(n_197),
.B1(n_219),
.B2(n_294),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_363),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_384),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_386),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_388),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_381),
.B(n_334),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_395),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_400),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_371),
.B(n_338),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_389),
.B(n_339),
.Y(n_435)
);

AOI22x1_ASAP7_75t_SL g436 ( 
.A1(n_383),
.A2(n_197),
.B1(n_308),
.B2(n_307),
.Y(n_436)
);

OAI22x1_ASAP7_75t_L g437 ( 
.A1(n_382),
.A2(n_385),
.B1(n_402),
.B2(n_401),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_403),
.Y(n_438)
);

INVx6_ASAP7_75t_L g439 ( 
.A(n_396),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_398),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_379),
.B(n_342),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_366),
.B(n_360),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_374),
.B(n_360),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_405),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_391),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_369),
.B(n_341),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_397),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_375),
.B(n_284),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_378),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_380),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_387),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_391),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_368),
.B(n_360),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_393),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_392),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_392),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_372),
.B(n_292),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_392),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_392),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_392),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_392),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_364),
.B(n_336),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_365),
.B(n_220),
.Y(n_466)
);

AOI22x1_ASAP7_75t_SL g467 ( 
.A1(n_364),
.A2(n_308),
.B1(n_307),
.B2(n_309),
.Y(n_467)
);

BUFx12f_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_370),
.B(n_295),
.Y(n_469)
);

OA21x2_ASAP7_75t_L g470 ( 
.A1(n_392),
.A2(n_348),
.B(n_324),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_370),
.B(n_200),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_365),
.B(n_222),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_370),
.B(n_200),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_392),
.A2(n_227),
.B(n_223),
.Y(n_474)
);

BUFx12f_ASAP7_75t_L g475 ( 
.A(n_394),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_L g476 ( 
.A(n_406),
.B(n_329),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_372),
.B(n_230),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_448),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_458),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_461),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_461),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_190),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_474),
.A2(n_34),
.B(n_33),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_408),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_462),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_440),
.B(n_201),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_452),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_443),
.B(n_204),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_427),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_408),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_438),
.B(n_35),
.Y(n_492)
);

OA21x2_ASAP7_75t_L g493 ( 
.A1(n_474),
.A2(n_218),
.B(n_216),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_464),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_448),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_438),
.B(n_36),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_184),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_438),
.B(n_429),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_463),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_473),
.B(n_184),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_429),
.B(n_41),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g504 ( 
.A(n_408),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_473),
.B(n_192),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_415),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_431),
.B(n_224),
.Y(n_507)
);

NAND3xp33_ASAP7_75t_L g508 ( 
.A(n_449),
.B(n_213),
.C(n_193),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_420),
.B(n_214),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_416),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_423),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_412),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_420),
.B(n_226),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_433),
.B(n_221),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_429),
.B(n_42),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_431),
.B(n_225),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_457),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_460),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_416),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_478),
.Y(n_522)
);

BUFx10_ASAP7_75t_L g523 ( 
.A(n_490),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_488),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_490),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_489),
.A2(n_449),
.B1(n_469),
.B2(n_427),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_488),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_492),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_506),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_496),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_499),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_R g532 ( 
.A(n_492),
.B(n_451),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_505),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_499),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_486),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_487),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_485),
.Y(n_537)
);

BUFx10_ASAP7_75t_L g538 ( 
.A(n_492),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_486),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_485),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_499),
.B(n_433),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_484),
.A2(n_411),
.B(n_470),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_509),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_L g544 ( 
.A(n_508),
.B(n_451),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_513),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_499),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_505),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_R g548 ( 
.A(n_500),
.B(n_451),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_513),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_509),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_492),
.Y(n_551)
);

NOR2xp67_ASAP7_75t_L g552 ( 
.A(n_507),
.B(n_453),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_514),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_494),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_514),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_519),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_497),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_497),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_515),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_518),
.B(n_444),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_L g561 ( 
.A(n_551),
.B(n_455),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_545),
.Y(n_562)
);

INVxp67_ASAP7_75t_SL g563 ( 
.A(n_532),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_549),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_523),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_553),
.Y(n_566)
);

BUFx10_ASAP7_75t_L g567 ( 
.A(n_525),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_555),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_535),
.Y(n_569)
);

OAI22xp33_ASAP7_75t_L g570 ( 
.A1(n_526),
.A2(n_483),
.B1(n_430),
.B2(n_432),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_535),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_539),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_556),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_539),
.Y(n_574)
);

OAI21xp33_ASAP7_75t_L g575 ( 
.A1(n_560),
.A2(n_469),
.B(n_417),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_554),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_550),
.A2(n_459),
.B1(n_454),
.B2(n_439),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_552),
.B(n_428),
.Y(n_578)
);

OAI22x1_ASAP7_75t_L g579 ( 
.A1(n_547),
.A2(n_465),
.B1(n_441),
.B2(n_445),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_554),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_542),
.Y(n_581)
);

CKINVDCx6p67_ASAP7_75t_R g582 ( 
.A(n_523),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_550),
.A2(n_498),
.B1(n_472),
.B2(n_502),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_541),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_541),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_543),
.B(n_498),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_559),
.A2(n_472),
.B1(n_430),
.B2(n_432),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_544),
.B(n_428),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_531),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_530),
.B(n_515),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_523),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_541),
.Y(n_592)
);

AO22x2_ASAP7_75t_L g593 ( 
.A1(n_537),
.A2(n_413),
.B1(n_426),
.B2(n_519),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_527),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_524),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_534),
.Y(n_596)
);

HAxp5_ASAP7_75t_SL g597 ( 
.A(n_559),
.B(n_410),
.CON(n_597),
.SN(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_540),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_540),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_546),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_557),
.B(n_428),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_529),
.Y(n_602)
);

INVx8_ASAP7_75t_L g603 ( 
.A(n_537),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_528),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_522),
.B(n_497),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_528),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_528),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_558),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_533),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_SL g610 ( 
.A1(n_536),
.A2(n_436),
.B1(n_409),
.B2(n_439),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_536),
.B(n_465),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_538),
.B(n_497),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_538),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_548),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_538),
.B(n_428),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_542),
.A2(n_477),
.B(n_493),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_525),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_527),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_545),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_535),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_560),
.B(n_452),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_560),
.B(n_452),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_560),
.B(n_433),
.Y(n_623)
);

BUFx8_ASAP7_75t_SL g624 ( 
.A(n_525),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_541),
.B(n_503),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_545),
.Y(n_626)
);

OA22x2_ASAP7_75t_L g627 ( 
.A1(n_526),
.A2(n_437),
.B1(n_446),
.B2(n_419),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_560),
.B(n_452),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_541),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_530),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_525),
.B(n_468),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_560),
.B(n_447),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_560),
.B(n_447),
.Y(n_633)
);

BUFx6f_ASAP7_75t_SL g634 ( 
.A(n_523),
.Y(n_634)
);

NAND3xp33_ASAP7_75t_L g635 ( 
.A(n_560),
.B(n_447),
.C(n_418),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_535),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_535),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_560),
.B(n_433),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_535),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_535),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_535),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_560),
.B(n_450),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_545),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_545),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_SL g645 ( 
.A(n_532),
.B(n_503),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_535),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_569),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_584),
.B(n_503),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_610),
.A2(n_437),
.B1(n_446),
.B2(n_439),
.Y(n_649)
);

BUFx10_ASAP7_75t_L g650 ( 
.A(n_617),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_567),
.Y(n_651)
);

INVxp33_ASAP7_75t_L g652 ( 
.A(n_590),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_600),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_566),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_603),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_566),
.B(n_479),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_584),
.B(n_503),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_621),
.B(n_622),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_562),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_603),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_623),
.B(n_479),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_624),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_571),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_600),
.Y(n_664)
);

AND2x2_ASAP7_75t_SL g665 ( 
.A(n_561),
.B(n_517),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_564),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_632),
.B(n_414),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_595),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_595),
.Y(n_669)
);

AND2x6_ASAP7_75t_L g670 ( 
.A(n_625),
.B(n_604),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_568),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_633),
.B(n_433),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_573),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_600),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_600),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_586),
.B(n_472),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_592),
.B(n_466),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_603),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_608),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_628),
.B(n_466),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_642),
.B(n_419),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_624),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_642),
.B(n_630),
.Y(n_683)
);

INVx5_ASAP7_75t_L g684 ( 
.A(n_565),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_619),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_626),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_572),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_643),
.Y(n_688)
);

AOI21x1_ASAP7_75t_L g689 ( 
.A1(n_616),
.A2(n_493),
.B(n_484),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_644),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_635),
.B(n_442),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_576),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_574),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_620),
.Y(n_694)
);

AND2x6_ASAP7_75t_L g695 ( 
.A(n_625),
.B(n_517),
.Y(n_695)
);

INVx5_ASAP7_75t_L g696 ( 
.A(n_591),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_636),
.Y(n_697)
);

AND2x6_ASAP7_75t_L g698 ( 
.A(n_604),
.B(n_517),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_623),
.B(n_480),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_608),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_580),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_638),
.B(n_480),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_639),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_639),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_611),
.B(n_414),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_640),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_618),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_585),
.B(n_517),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_608),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_618),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_640),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_637),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_585),
.B(n_466),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_575),
.B(n_520),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_638),
.B(n_481),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_629),
.B(n_520),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_563),
.B(n_481),
.Y(n_717)
);

AND2x6_ASAP7_75t_L g718 ( 
.A(n_606),
.B(n_501),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_563),
.B(n_482),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_641),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_646),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_646),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_570),
.B(n_442),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_570),
.B(n_435),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_598),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_599),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_627),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_629),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_627),
.Y(n_729)
);

AO21x2_ASAP7_75t_L g730 ( 
.A1(n_581),
.A2(n_512),
.B(n_511),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_726),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_725),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_659),
.Y(n_733)
);

NAND2x1p5_ASAP7_75t_L g734 ( 
.A(n_684),
.B(n_588),
.Y(n_734)
);

AO22x2_ASAP7_75t_L g735 ( 
.A1(n_727),
.A2(n_577),
.B1(n_581),
.B2(n_578),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_667),
.B(n_589),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_665),
.B(n_645),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_666),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_671),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_673),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_685),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_686),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_684),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_649),
.A2(n_691),
.B1(n_561),
.B2(n_724),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_688),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_668),
.B(n_608),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_690),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_669),
.B(n_674),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_721),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_664),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_654),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_709),
.B(n_596),
.Y(n_752)
);

NAND3x1_ASAP7_75t_L g753 ( 
.A(n_683),
.B(n_681),
.C(n_705),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_692),
.Y(n_754)
);

OAI221xp5_ASAP7_75t_L g755 ( 
.A1(n_649),
.A2(n_583),
.B1(n_610),
.B2(n_587),
.C(n_645),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_658),
.B(n_588),
.Y(n_756)
);

AO21x2_ASAP7_75t_L g757 ( 
.A1(n_689),
.A2(n_723),
.B(n_656),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_701),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_664),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_729),
.B(n_579),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_703),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_724),
.A2(n_583),
.B(n_587),
.C(n_578),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_647),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_656),
.B(n_601),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_684),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_704),
.B(n_601),
.Y(n_766)
);

AO22x2_ASAP7_75t_L g767 ( 
.A1(n_661),
.A2(n_613),
.B1(n_607),
.B2(n_615),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_706),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_652),
.B(n_605),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_711),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_680),
.B(n_605),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_664),
.Y(n_772)
);

OAI22xp33_ASAP7_75t_L g773 ( 
.A1(n_707),
.A2(n_605),
.B1(n_631),
.B2(n_582),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_720),
.Y(n_774)
);

INVx6_ASAP7_75t_L g775 ( 
.A(n_650),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_661),
.B(n_594),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_676),
.B(n_593),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_663),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_722),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_699),
.B(n_612),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_699),
.Y(n_781)
);

AND2x6_ASAP7_75t_L g782 ( 
.A(n_648),
.B(n_511),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_675),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_687),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_693),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_702),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_653),
.B(n_614),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_694),
.Y(n_788)
);

NAND2x1p5_ASAP7_75t_L g789 ( 
.A(n_696),
.B(n_615),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_675),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_697),
.Y(n_791)
);

OAI221xp5_ASAP7_75t_L g792 ( 
.A1(n_672),
.A2(n_611),
.B1(n_236),
.B2(n_231),
.C(n_456),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_714),
.A2(n_593),
.B1(n_439),
.B2(n_609),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_675),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_712),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_730),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_679),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_716),
.Y(n_798)
);

AO22x2_ASAP7_75t_L g799 ( 
.A1(n_715),
.A2(n_597),
.B1(n_602),
.B2(n_467),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_715),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_714),
.B(n_634),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_716),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_679),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_717),
.B(n_612),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_743),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_776),
.B(n_672),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_773),
.B(n_696),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_753),
.B(n_662),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_731),
.B(n_717),
.Y(n_809)
);

OR2x6_ASAP7_75t_L g810 ( 
.A(n_737),
.B(n_653),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_781),
.B(n_719),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_738),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_775),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_733),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_786),
.B(n_719),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_800),
.B(n_700),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_744),
.A2(n_695),
.B1(n_593),
.B2(n_651),
.Y(n_817)
);

INVxp67_ASAP7_75t_L g818 ( 
.A(n_736),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_739),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_740),
.Y(n_820)
);

NAND2xp33_ASAP7_75t_L g821 ( 
.A(n_799),
.B(n_682),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_745),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_747),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_801),
.B(n_775),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_764),
.B(n_700),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_775),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_764),
.B(n_700),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_741),
.B(n_728),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_746),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_750),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_742),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_743),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_732),
.B(n_728),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_754),
.B(n_758),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_751),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_769),
.B(n_696),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_755),
.A2(n_695),
.B1(n_634),
.B2(n_708),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_804),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_773),
.B(n_707),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_761),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_769),
.B(n_670),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_804),
.B(n_670),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_768),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_770),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_755),
.A2(n_695),
.B1(n_708),
.B2(n_612),
.Y(n_845)
);

INVxp67_ASAP7_75t_SL g846 ( 
.A(n_756),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_801),
.B(n_710),
.Y(n_847)
);

INVxp33_ASAP7_75t_L g848 ( 
.A(n_746),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_748),
.B(n_670),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_748),
.B(n_670),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_SL g851 ( 
.A(n_792),
.B(n_602),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_792),
.A2(n_713),
.B1(n_677),
.B2(n_695),
.Y(n_852)
);

NOR2xp67_ASAP7_75t_L g853 ( 
.A(n_765),
.B(n_710),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_760),
.B(n_718),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_763),
.B(n_718),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_798),
.B(n_655),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_778),
.B(n_718),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_784),
.B(n_785),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_788),
.B(n_718),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_SL g860 ( 
.A(n_787),
.B(n_650),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_772),
.Y(n_861)
);

AND3x1_ASAP7_75t_L g862 ( 
.A(n_793),
.B(n_660),
.C(n_655),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_791),
.B(n_648),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_787),
.B(n_678),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_774),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_762),
.A2(n_609),
.B(n_698),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_771),
.B(n_567),
.Y(n_867)
);

INVxp67_ASAP7_75t_SL g868 ( 
.A(n_756),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_795),
.B(n_657),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_799),
.A2(n_657),
.B1(n_698),
.B2(n_612),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_779),
.B(n_698),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_737),
.A2(n_422),
.B(n_476),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_SL g873 ( 
.A1(n_799),
.A2(n_698),
.B1(n_612),
.B2(n_456),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_766),
.B(n_730),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_752),
.B(n_660),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_772),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_749),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_766),
.B(n_678),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_793),
.A2(n_235),
.B(n_442),
.C(n_435),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_750),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_780),
.B(n_493),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_771),
.B(n_468),
.Y(n_882)
);

AND2x6_ASAP7_75t_SL g883 ( 
.A(n_777),
.B(n_434),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_846),
.B(n_780),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_812),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_805),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_851),
.A2(n_735),
.B1(n_762),
.B2(n_802),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_873),
.B(n_750),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_831),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_824),
.B(n_475),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_838),
.B(n_767),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_826),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_819),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_820),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_868),
.B(n_757),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_818),
.B(n_767),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_806),
.B(n_757),
.Y(n_897)
);

OAI21xp33_ASAP7_75t_L g898 ( 
.A1(n_870),
.A2(n_866),
.B(n_735),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_R g899 ( 
.A(n_808),
.B(n_475),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_830),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_805),
.B(n_790),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_822),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_874),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_860),
.B(n_870),
.Y(n_904)
);

INVxp33_ASAP7_75t_L g905 ( 
.A(n_847),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_813),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_861),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_825),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_848),
.B(n_767),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_827),
.B(n_735),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_828),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_832),
.B(n_790),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_832),
.B(n_797),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_842),
.B(n_829),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_875),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_840),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_814),
.B(n_796),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_821),
.A2(n_734),
.B(n_789),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_823),
.B(n_796),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_876),
.B(n_797),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_810),
.B(n_783),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_810),
.B(n_803),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_810),
.B(n_876),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_830),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_877),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_811),
.B(n_803),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_815),
.B(n_750),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_836),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_849),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_843),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_830),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_844),
.B(n_789),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_809),
.B(n_858),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_878),
.B(n_759),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_880),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_865),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_835),
.B(n_759),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_834),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_881),
.B(n_734),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_914),
.B(n_867),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_918),
.B(n_853),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_887),
.A2(n_817),
.B(n_807),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_898),
.A2(n_839),
.B(n_879),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_911),
.B(n_816),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_897),
.A2(n_882),
.B(n_864),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_900),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_888),
.A2(n_837),
.B(n_872),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_938),
.B(n_833),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_904),
.A2(n_852),
.B(n_862),
.Y(n_949)
);

OAI321xp33_ASAP7_75t_L g950 ( 
.A1(n_910),
.A2(n_852),
.A3(n_845),
.B1(n_857),
.B2(n_855),
.C(n_859),
.Y(n_950)
);

OAI21xp33_ASAP7_75t_L g951 ( 
.A1(n_895),
.A2(n_884),
.B(n_896),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_905),
.A2(n_871),
.B(n_841),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_908),
.B(n_854),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_928),
.B(n_863),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_905),
.A2(n_850),
.B(n_869),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_890),
.A2(n_856),
.B(n_883),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_933),
.A2(n_856),
.B(n_794),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_903),
.B(n_880),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_926),
.A2(n_794),
.B(n_759),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_914),
.B(n_880),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_929),
.A2(n_794),
.B(n_493),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_899),
.B(n_794),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_902),
.B(n_782),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_925),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_896),
.B(n_782),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_906),
.B(n_434),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_893),
.Y(n_967)
);

BUFx8_ASAP7_75t_SL g968 ( 
.A(n_906),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_921),
.A2(n_435),
.B(n_434),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_892),
.B(n_221),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_930),
.Y(n_971)
);

NAND2x1p5_ASAP7_75t_L g972 ( 
.A(n_923),
.B(n_782),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_892),
.B(n_0),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_921),
.A2(n_516),
.B(n_425),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_907),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_921),
.A2(n_516),
.B(n_424),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_932),
.B(n_782),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_939),
.A2(n_516),
.B(n_2),
.C(n_3),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_SL g979 ( 
.A(n_892),
.B(n_504),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_932),
.B(n_1),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_939),
.A2(n_516),
.B(n_232),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_927),
.B(n_1),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_923),
.A2(n_232),
.B(n_421),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_891),
.B(n_2),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_901),
.B(n_3),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_923),
.B(n_4),
.Y(n_986)
);

AND2x2_ASAP7_75t_SL g987 ( 
.A(n_922),
.B(n_232),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_891),
.B(n_4),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_922),
.A2(n_232),
.B(n_421),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_909),
.A2(n_229),
.B(n_228),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_885),
.B(n_5),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_901),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_934),
.A2(n_234),
.B(n_233),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_894),
.B(n_6),
.Y(n_994)
);

OA22x2_ASAP7_75t_L g995 ( 
.A1(n_942),
.A2(n_915),
.B1(n_912),
.B2(n_913),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_943),
.A2(n_894),
.B(n_912),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_970),
.A2(n_947),
.B(n_949),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_990),
.A2(n_913),
.B(n_912),
.Y(n_998)
);

NAND3xp33_ASAP7_75t_SL g999 ( 
.A(n_942),
.B(n_920),
.C(n_937),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_979),
.B(n_913),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_946),
.Y(n_1001)
);

NAND3xp33_ASAP7_75t_L g1002 ( 
.A(n_990),
.B(n_919),
.C(n_917),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_978),
.A2(n_886),
.B(n_936),
.C(n_935),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_984),
.B(n_937),
.Y(n_1004)
);

NOR3xp33_ASAP7_75t_L g1005 ( 
.A(n_950),
.B(n_886),
.C(n_924),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_987),
.A2(n_919),
.B(n_917),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_968),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_941),
.A2(n_916),
.B(n_889),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_993),
.A2(n_916),
.B(n_889),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_967),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_973),
.A2(n_886),
.B(n_924),
.C(n_935),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_979),
.A2(n_920),
.B1(n_931),
.B2(n_900),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_988),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_975),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_997),
.B(n_950),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_1003),
.A2(n_962),
.B(n_956),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_1007),
.B(n_991),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_1010),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_996),
.A2(n_994),
.B(n_983),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_995),
.A2(n_972),
.B1(n_992),
.B2(n_965),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_1007),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_1002),
.A2(n_972),
.B1(n_966),
.B2(n_952),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_1013),
.A2(n_964),
.B1(n_980),
.B2(n_955),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1004),
.B(n_986),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_999),
.A2(n_989),
.B(n_961),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1001),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_998),
.B(n_957),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_1005),
.B(n_985),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_1014),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1009),
.Y(n_1030)
);

CKINVDCx14_ASAP7_75t_R g1031 ( 
.A(n_1012),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1008),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_1011),
.A2(n_1000),
.B(n_1006),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1013),
.B(n_951),
.Y(n_1034)
);

NOR3xp33_ASAP7_75t_SL g1035 ( 
.A(n_999),
.B(n_982),
.C(n_981),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1010),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_1001),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_1001),
.B(n_946),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1010),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_1021),
.B(n_940),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1030),
.B(n_948),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_1021),
.B(n_945),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1031),
.B(n_960),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1018),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_1029),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1036),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1038),
.B(n_946),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_1042),
.A2(n_1015),
.B(n_1028),
.Y(n_1048)
);

NOR3xp33_ASAP7_75t_L g1049 ( 
.A(n_1044),
.B(n_1040),
.C(n_1043),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_1047),
.A2(n_1016),
.B(n_1033),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_1050),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_1049),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1052),
.A2(n_1048),
.B1(n_1045),
.B2(n_1040),
.Y(n_1053)
);

OR2x6_ASAP7_75t_L g1054 ( 
.A(n_1051),
.B(n_1017),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1053),
.B(n_1046),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_1054),
.A2(n_1023),
.B(n_1027),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1056),
.B(n_1032),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1055),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1058),
.B(n_1037),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1057),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1060),
.Y(n_1061)
);

AO21x2_ASAP7_75t_L g1062 ( 
.A1(n_1059),
.A2(n_1041),
.B(n_1034),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1062),
.B(n_1026),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1061),
.A2(n_1038),
.B1(n_1025),
.B2(n_1020),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1062),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1065),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1064),
.B(n_1039),
.Y(n_1067)
);

INVxp67_ASAP7_75t_SL g1068 ( 
.A(n_1063),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1067),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_1066),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_1070),
.B(n_1069),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1069),
.B(n_1068),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1072),
.B(n_1024),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_1071),
.A2(n_1023),
.B1(n_1019),
.B2(n_1022),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_1073),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1074),
.B(n_1035),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1075),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_1076),
.B(n_953),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1078),
.B(n_944),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1077),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_1080),
.B(n_7),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1079),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1079),
.B(n_954),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1081),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_1082),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_1083),
.B(n_7),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1085),
.A2(n_958),
.B1(n_900),
.B2(n_931),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1086),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1088),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1087),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1089),
.B(n_1084),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_1090),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_1091),
.B(n_8),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1092),
.B(n_971),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_1093),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1094),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1095),
.B(n_9),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1096),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_1098),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_1099)
);

INVxp67_ASAP7_75t_L g1100 ( 
.A(n_1097),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_1097),
.Y(n_1101)
);

AOI21xp33_ASAP7_75t_L g1102 ( 
.A1(n_1100),
.A2(n_12),
.B(n_13),
.Y(n_1102)
);

OA21x2_ASAP7_75t_L g1103 ( 
.A1(n_1099),
.A2(n_14),
.B(n_15),
.Y(n_1103)
);

AOI22x1_ASAP7_75t_L g1104 ( 
.A1(n_1101),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1103),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_1102),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_SL g1107 ( 
.A1(n_1105),
.A2(n_1104),
.B1(n_17),
.B2(n_18),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_1106),
.Y(n_1108)
);

NAND4xp75_ASAP7_75t_L g1109 ( 
.A(n_1108),
.B(n_16),
.C(n_18),
.D(n_19),
.Y(n_1109)
);

AND3x1_ASAP7_75t_L g1110 ( 
.A(n_1107),
.B(n_19),
.C(n_20),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1110),
.Y(n_1111)
);

NOR3xp33_ASAP7_75t_L g1112 ( 
.A(n_1109),
.B(n_20),
.C(n_21),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1111),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1112),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1113),
.B(n_22),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_L g1116 ( 
.A(n_1114),
.B(n_23),
.C(n_24),
.Y(n_1116)
);

AOI222xp33_ASAP7_75t_L g1117 ( 
.A1(n_1115),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.C1(n_26),
.C2(n_27),
.Y(n_1117)
);

OAI211xp5_ASAP7_75t_L g1118 ( 
.A1(n_1116),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_1118)
);

AOI221xp5_ASAP7_75t_L g1119 ( 
.A1(n_1116),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.C(n_44),
.Y(n_1119)
);

NAND3xp33_ASAP7_75t_L g1120 ( 
.A(n_1118),
.B(n_30),
.C(n_900),
.Y(n_1120)
);

NOR3xp33_ASAP7_75t_L g1121 ( 
.A(n_1119),
.B(n_45),
.C(n_47),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1117),
.B(n_49),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1122),
.Y(n_1123)
);

NOR2x1_ASAP7_75t_L g1124 ( 
.A(n_1120),
.B(n_51),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1123),
.A2(n_1121),
.B(n_52),
.Y(n_1125)
);

NAND4xp25_ASAP7_75t_L g1126 ( 
.A(n_1124),
.B(n_53),
.C(n_54),
.D(n_56),
.Y(n_1126)
);

INVxp67_ASAP7_75t_SL g1127 ( 
.A(n_1125),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1126),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_SL g1129 ( 
.A1(n_1127),
.A2(n_58),
.B(n_59),
.Y(n_1129)
);

NOR3xp33_ASAP7_75t_L g1130 ( 
.A(n_1128),
.B(n_60),
.C(n_62),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1129),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_1130),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.C(n_67),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1131),
.Y(n_1133)
);

XNOR2x1_ASAP7_75t_L g1134 ( 
.A(n_1132),
.B(n_68),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1133),
.Y(n_1135)
);

AOI22x1_ASAP7_75t_L g1136 ( 
.A1(n_1134),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1133),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1135),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1137),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1136),
.B(n_74),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_1139),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1138),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1142),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1141),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_1143),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_1144),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1146),
.B(n_1140),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_L g1148 ( 
.A(n_1145),
.B(n_75),
.C(n_76),
.Y(n_1148)
);

XOR2x2_ASAP7_75t_L g1149 ( 
.A(n_1147),
.B(n_78),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1148),
.A2(n_931),
.B1(n_900),
.B2(n_969),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1149),
.B(n_1150),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1149),
.A2(n_931),
.B1(n_521),
.B2(n_510),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1151),
.Y(n_1153)
);

XNOR2xp5_ASAP7_75t_L g1154 ( 
.A(n_1152),
.B(n_79),
.Y(n_1154)
);

XOR2xp5_ASAP7_75t_L g1155 ( 
.A(n_1151),
.B(n_80),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1153),
.A2(n_931),
.B1(n_521),
.B2(n_510),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1154),
.A2(n_81),
.B(n_83),
.C(n_84),
.Y(n_1157)
);

AOI21xp33_ASAP7_75t_SL g1158 ( 
.A1(n_1155),
.A2(n_85),
.B(n_89),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1153),
.B(n_91),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1158),
.A2(n_92),
.B1(n_94),
.B2(n_97),
.Y(n_1160)
);

OA21x2_ASAP7_75t_L g1161 ( 
.A1(n_1159),
.A2(n_98),
.B(n_99),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1157),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1162),
.B(n_1156),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1161),
.A2(n_102),
.B(n_103),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_SL g1165 ( 
.A1(n_1160),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_1165)
);

NOR2xp67_ASAP7_75t_L g1166 ( 
.A(n_1163),
.B(n_110),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1164),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1165),
.A2(n_113),
.B(n_114),
.Y(n_1168)
);

AOI21xp33_ASAP7_75t_SL g1169 ( 
.A1(n_1163),
.A2(n_116),
.B(n_117),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1163),
.A2(n_510),
.B1(n_521),
.B2(n_495),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1163),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_SL g1172 ( 
.A1(n_1163),
.A2(n_123),
.B(n_125),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1163),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1163),
.B(n_126),
.Y(n_1174)
);

XNOR2xp5_ASAP7_75t_L g1175 ( 
.A(n_1163),
.B(n_127),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1163),
.A2(n_128),
.B(n_130),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1163),
.A2(n_491),
.B1(n_485),
.B2(n_495),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1173),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1167),
.A2(n_1168),
.B1(n_1172),
.B2(n_1175),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_1174),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1166),
.B(n_131),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1169),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1176),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1171),
.B(n_132),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1170),
.Y(n_1185)
);

OAI221xp5_ASAP7_75t_L g1186 ( 
.A1(n_1177),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.C(n_137),
.Y(n_1186)
);

OA21x2_ASAP7_75t_L g1187 ( 
.A1(n_1178),
.A2(n_138),
.B(n_140),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1183),
.A2(n_141),
.B(n_142),
.Y(n_1188)
);

AOI222xp33_ASAP7_75t_L g1189 ( 
.A1(n_1179),
.A2(n_143),
.B1(n_144),
.B2(n_146),
.C1(n_147),
.C2(n_148),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1182),
.Y(n_1190)
);

AO221x1_ASAP7_75t_L g1191 ( 
.A1(n_1180),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.C(n_153),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1185),
.A2(n_155),
.B(n_156),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1184),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_1193)
);

OA21x2_ASAP7_75t_L g1194 ( 
.A1(n_1190),
.A2(n_1181),
.B(n_1186),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1187),
.A2(n_1193),
.B(n_1188),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1191),
.B(n_162),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1194),
.A2(n_1192),
.B1(n_1189),
.B2(n_166),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1197),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_1198),
.A2(n_1195),
.B(n_1196),
.Y(n_1199)
);

OAI221xp5_ASAP7_75t_R g1200 ( 
.A1(n_1199),
.A2(n_163),
.B1(n_164),
.B2(n_167),
.C(n_168),
.Y(n_1200)
);

AOI221xp5_ASAP7_75t_L g1201 ( 
.A1(n_1200),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.C(n_173),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1201),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_1202)
);

AOI211xp5_ASAP7_75t_L g1203 ( 
.A1(n_1202),
.A2(n_177),
.B(n_977),
.C(n_959),
.Y(n_1203)
);

AOI211xp5_ASAP7_75t_L g1204 ( 
.A1(n_1203),
.A2(n_963),
.B(n_976),
.C(n_974),
.Y(n_1204)
);


endmodule