module fake_jpeg_28956_n_415 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_415);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_415;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_30),
.Y(n_53)
);

INVx5_ASAP7_75t_SL g120 ( 
.A(n_53),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_19),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_54),
.Y(n_122)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_55),
.Y(n_141)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_13),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_57),
.B(n_60),
.Y(n_145)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_13),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_11),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_63),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_20),
.B(n_11),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_71),
.B(n_78),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_39),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_23),
.B(n_10),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_23),
.B(n_35),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_83),
.Y(n_143)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_32),
.B(n_10),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_96),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_32),
.B(n_35),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_41),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_48),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_47),
.B1(n_48),
.B2(n_46),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_98),
.A2(n_107),
.B1(n_133),
.B2(n_136),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_61),
.A2(n_47),
.B1(n_48),
.B2(n_46),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_109),
.B(n_79),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_47),
.B1(n_25),
.B2(n_26),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_46),
.B1(n_22),
.B2(n_44),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_112),
.A2(n_123),
.B1(n_124),
.B2(n_53),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_51),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_53),
.B1(n_50),
.B2(n_76),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_44),
.B1(n_45),
.B2(n_43),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_45),
.B1(n_31),
.B2(n_42),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_135),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_72),
.A2(n_94),
.B1(n_93),
.B2(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_58),
.B(n_39),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_91),
.A2(n_36),
.B1(n_26),
.B2(n_25),
.Y(n_136)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_89),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_180),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_145),
.B(n_105),
.C(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_153),
.B(n_164),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_154),
.A2(n_157),
.B1(n_183),
.B2(n_188),
.Y(n_198)
);

NAND2x1_ASAP7_75t_SL g156 ( 
.A(n_112),
.B(n_120),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_156),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_88),
.B1(n_87),
.B2(n_64),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_56),
.B1(n_52),
.B2(n_77),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_158),
.A2(n_134),
.B1(n_129),
.B2(n_103),
.Y(n_220)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

INVx4_ASAP7_75t_SL g161 ( 
.A(n_120),
.Y(n_161)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_161),
.Y(n_225)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_102),
.Y(n_164)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_169),
.B(n_170),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_102),
.Y(n_170)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_125),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_97),
.Y(n_174)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_130),
.B(n_67),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_122),
.C(n_99),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_100),
.Y(n_176)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_106),
.A2(n_80),
.B1(n_86),
.B2(n_84),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_122),
.B1(n_144),
.B2(n_132),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_111),
.B(n_42),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_54),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_123),
.A2(n_73),
.B1(n_65),
.B2(n_70),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_184),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_27),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_19),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_103),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_186),
.Y(n_223)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_138),
.A2(n_36),
.B1(n_27),
.B2(n_75),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_116),
.B(n_54),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_190),
.Y(n_204)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_108),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_108),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_192),
.A2(n_220),
.B1(n_161),
.B2(n_183),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_205),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_150),
.B(n_147),
.C(n_131),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_211),
.C(n_175),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_19),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_168),
.A2(n_131),
.B1(n_144),
.B2(n_132),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_156),
.B(n_165),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_195),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g217 ( 
.A1(n_156),
.A2(n_134),
.B1(n_129),
.B2(n_124),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_222),
.B(n_184),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_185),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_233),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_216),
.A2(n_165),
.B1(n_168),
.B2(n_167),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_245),
.B1(n_220),
.B2(n_205),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_209),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_231),
.B(n_234),
.Y(n_274)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_225),
.Y(n_232)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_175),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_236),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_238),
.A2(n_247),
.B1(n_198),
.B2(n_215),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_163),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_239),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_221),
.A2(n_161),
.B(n_190),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_249),
.B(n_204),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_153),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_244),
.C(n_206),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_178),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_248),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_178),
.C(n_187),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_221),
.A2(n_142),
.B1(n_191),
.B2(n_162),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_195),
.A2(n_155),
.B1(n_159),
.B2(n_142),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_164),
.Y(n_248)
);

NAND2xp33_ASAP7_75t_R g249 ( 
.A(n_216),
.B(n_173),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_223),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_202),
.A2(n_170),
.B(n_19),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_254),
.B(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_252),
.B(n_205),
.Y(n_258)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_208),
.Y(n_253)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_195),
.A2(n_19),
.B(n_31),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_255),
.A2(n_268),
.B1(n_247),
.B2(n_254),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_248),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_257),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_272),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_269),
.B1(n_246),
.B2(n_245),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_265),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_217),
.B1(n_198),
.B2(n_204),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_241),
.A2(n_217),
.B1(n_199),
.B2(n_204),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_233),
.B(n_217),
.Y(n_271)
);

XNOR2x1_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_276),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_226),
.B(n_243),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_229),
.B(n_213),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_275),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_228),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_253),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_236),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_252),
.B(n_212),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_230),
.Y(n_295)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_240),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_283),
.Y(n_305)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_264),
.Y(n_284)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_240),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_285),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_286),
.A2(n_291),
.B1(n_275),
.B2(n_256),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_257),
.A2(n_270),
.B1(n_263),
.B2(n_235),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_255),
.B1(n_258),
.B2(n_279),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_239),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_262),
.A2(n_227),
.B1(n_238),
.B2(n_232),
.Y(n_291)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_295),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_242),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_263),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_298),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_244),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_261),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_301),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_300),
.A2(n_267),
.B1(n_271),
.B2(n_227),
.Y(n_314)
);

OAI21xp33_ASAP7_75t_L g304 ( 
.A1(n_260),
.A2(n_251),
.B(n_227),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_304),
.A2(n_275),
.B(n_259),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_266),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_306),
.B(n_311),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_307),
.A2(n_319),
.B1(n_322),
.B2(n_302),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_266),
.C(n_276),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_325),
.C(n_326),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_298),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_314),
.A2(n_321),
.B1(n_289),
.B2(n_286),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_317),
.A2(n_289),
.B(n_285),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_273),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_196),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_300),
.A2(n_278),
.B1(n_277),
.B2(n_256),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_291),
.A2(n_278),
.B1(n_280),
.B2(n_200),
.Y(n_322)
);

NAND2x1p5_ASAP7_75t_L g323 ( 
.A(n_283),
.B(n_207),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_295),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_193),
.C(n_280),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_283),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_294),
.B(n_212),
.C(n_207),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_285),
.C(n_297),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_328),
.B(n_200),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_324),
.B(n_288),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_330),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_311),
.B(n_302),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_332),
.A2(n_315),
.B1(n_322),
.B2(n_323),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_333),
.A2(n_323),
.B(n_317),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_340),
.C(n_346),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_338),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_310),
.B(n_293),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_339),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_281),
.Y(n_337)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_337),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_290),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_325),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_308),
.B(n_284),
.C(n_282),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_309),
.Y(n_341)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_341),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_312),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_321),
.B(n_319),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_344),
.B(n_326),
.Y(n_354)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_309),
.Y(n_345)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_345),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_320),
.C(n_314),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_335),
.A2(n_316),
.B(n_305),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_347),
.A2(n_166),
.B(n_155),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_331),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_355),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_357),
.A2(n_362),
.B1(n_361),
.B2(n_359),
.Y(n_367)
);

AOI322xp5_ASAP7_75t_L g358 ( 
.A1(n_335),
.A2(n_315),
.A3(n_312),
.B1(n_313),
.B2(n_224),
.C1(n_151),
.C2(n_172),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_358),
.B(n_342),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_359),
.B(n_361),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_224),
.C(n_214),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_360),
.B(n_334),
.C(n_338),
.Y(n_365)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_335),
.Y(n_362)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_362),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_353),
.A2(n_331),
.B(n_339),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_363),
.A2(n_347),
.B(n_352),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_373),
.C(n_73),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_366),
.A2(n_369),
.B1(n_374),
.B2(n_360),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_367),
.B(n_351),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_368),
.B(n_356),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_357),
.A2(n_346),
.B1(n_343),
.B2(n_186),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_343),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_355),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_349),
.B(n_214),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_371),
.B(n_372),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_117),
.C(n_127),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_348),
.A2(n_171),
.B1(n_127),
.B2(n_152),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_378),
.A2(n_364),
.B1(n_370),
.B2(n_2),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_379),
.B(n_382),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_351),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_381),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_376),
.B(n_356),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_383),
.B(n_384),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_352),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_385),
.A2(n_1),
.B(n_2),
.Y(n_396)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_375),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_386),
.B(n_364),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_31),
.C(n_3),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_373),
.B(n_31),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_388),
.A2(n_372),
.B1(n_369),
.B2(n_367),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_394),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_393),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_377),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_395),
.A2(n_382),
.B1(n_3),
.B2(n_4),
.Y(n_402)
);

O2A1O1Ixp33_ASAP7_75t_SL g404 ( 
.A1(n_396),
.A2(n_392),
.B(n_394),
.C(n_393),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_397),
.B(n_1),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_391),
.B(n_380),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_402),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_389),
.A2(n_387),
.B(n_379),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_400),
.A2(n_398),
.B(n_401),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_403),
.B(n_3),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_397),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_405),
.A2(n_7),
.B(n_8),
.Y(n_411)
);

MAJx2_ASAP7_75t_L g409 ( 
.A(n_406),
.B(n_401),
.C(n_5),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_408),
.A2(n_4),
.B(n_5),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_409),
.A2(n_410),
.B(n_411),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_412),
.Y(n_413)
);

OAI221xp5_ASAP7_75t_L g414 ( 
.A1(n_413),
.A2(n_407),
.B1(n_8),
.B2(n_9),
.C(n_7),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_8),
.Y(n_415)
);


endmodule