module real_jpeg_17087_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_355),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_0),
.B(n_356),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_1),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_2),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_2),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_3),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_3),
.Y(n_208)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_4),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_4),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_5),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_5),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_5),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_5),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_5),
.B(n_280),
.Y(n_279)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_6),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_6),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g185 ( 
.A(n_6),
.B(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_6),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_6),
.B(n_204),
.Y(n_203)
);

AND2x4_ASAP7_75t_SL g207 ( 
.A(n_6),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_6),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_6),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_7),
.Y(n_187)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_8),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_9),
.Y(n_356)
);

AND2x4_ASAP7_75t_SL g24 ( 
.A(n_10),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_29),
.Y(n_28)
);

NAND2x1p5_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_33),
.Y(n_32)
);

NAND2x1_ASAP7_75t_L g65 ( 
.A(n_10),
.B(n_66),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_10),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_10),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_10),
.B(n_59),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_10),
.B(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_11),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_11),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_12),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_12),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_12),
.B(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_12),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_12),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_12),
.B(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_175),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_173),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_150),
.Y(n_18)
);

AND2x4_ASAP7_75t_SL g174 ( 
.A(n_19),
.B(n_150),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_86),
.C(n_111),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_20),
.B(n_86),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_60),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_21),
.B(n_61),
.C(n_72),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.C(n_46),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_22),
.B(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_22)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_23),
.A2(n_36),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_31),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_28),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_24),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_24),
.A2(n_63),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_24),
.B(n_89),
.C(n_95),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_24),
.A2(n_63),
.B1(n_139),
.B2(n_195),
.Y(n_261)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_40),
.B(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_28),
.B(n_32),
.C(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_28),
.A2(n_40),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_28),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_28),
.A2(n_116),
.B1(n_192),
.B2(n_198),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_29),
.Y(n_280)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_31),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_31),
.B(n_32),
.C(n_246),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_32),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_32),
.A2(n_37),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_32),
.A2(n_37),
.B1(n_246),
.B2(n_250),
.Y(n_245)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_36),
.A2(n_202),
.B(n_207),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_37),
.B(n_79),
.C(n_102),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_38),
.B(n_46),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_39),
.Y(n_271)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_40),
.A2(n_117),
.B1(n_203),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_40),
.A2(n_75),
.B1(n_117),
.B2(n_132),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_40),
.B(n_75),
.C(n_259),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_43),
.B(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_56),
.Y(n_46)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_48),
.A2(n_49),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_48),
.A2(n_49),
.B1(n_95),
.B2(n_96),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_52),
.C(n_110),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_49),
.A2(n_96),
.B(n_185),
.C(n_225),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_56),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_56),
.A2(n_81),
.B1(n_110),
.B2(n_131),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_56),
.B(n_131),
.C(n_189),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_56),
.A2(n_110),
.B1(n_246),
.B2(n_250),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_90),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_57),
.B(n_140),
.Y(n_139)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_72),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_62),
.B(n_65),
.C(n_68),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_63),
.B(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_65),
.A2(n_71),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_65),
.A2(n_71),
.B1(n_171),
.B2(n_172),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_65),
.B(n_96),
.C(n_126),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_73),
.C(n_83),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_67),
.A2(n_68),
.B1(n_142),
.B2(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_68),
.B(n_134),
.C(n_142),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_68),
.B(n_83),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_68),
.B(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_68),
.B(n_79),
.C(n_259),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_70),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_73),
.A2(n_74),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.C(n_81),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_75),
.A2(n_81),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_79),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_79),
.A2(n_101),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AO21x1_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_119),
.B(n_128),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_81),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_81),
.B(n_120),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_83),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_135),
.C(n_139),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_97),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_87),
.B(n_98),
.C(n_109),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_93),
.B2(n_94),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_89),
.A2(n_279),
.B(n_281),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_89),
.B(n_279),
.Y(n_281)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_95),
.B(n_126),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_95),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_95),
.B(n_232),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_109),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_110),
.B(n_250),
.C(n_291),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_111),
.B(n_328),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_133),
.C(n_146),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_112),
.B(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.C(n_129),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_118),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_120),
.A2(n_121),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_126),
.Y(n_128)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_125),
.A2(n_126),
.B1(n_207),
.B2(n_209),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_125),
.A2(n_126),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_126),
.A2(n_207),
.B(n_223),
.C(n_225),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_126),
.B(n_207),
.Y(n_225)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_129),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_133),
.A2(n_146),
.B1(n_147),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_133),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_134),
.B(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_135),
.A2(n_139),
.B1(n_195),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_135),
.Y(n_303)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_139),
.Y(n_195)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_142),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_164),
.Y(n_152)
);

XNOR2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_163),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_162),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI321xp33_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_309),
.A3(n_342),
.B1(n_348),
.B2(n_353),
.C(n_354),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_284),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_263),
.B(n_283),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_240),
.B(n_262),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_220),
.B(n_239),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_199),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_199),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_191),
.C(n_196),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_185),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_185),
.A2(n_189),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_191),
.A2(n_196),
.B1(n_197),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_191),
.A2(n_192),
.B(n_195),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_210),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_211),
.C(n_219),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_206),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_231),
.B(n_233),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_218),
.B2(n_219),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_215),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_215),
.A2(n_259),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_229),
.B(n_238),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_226),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_235),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_234),
.B(n_237),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_242),
.Y(n_262)
);

XOR2x2_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_252),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_251),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_251),
.C(n_252),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_246),
.Y(n_250)
);

OR2x6_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_257),
.C(n_261),
.Y(n_267)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_265),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_275),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_268),
.C(n_275),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_272),
.C(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_282),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_278),
.C(n_282),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_281),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_285),
.B(n_286),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_299),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_287),
.B(n_300),
.C(n_308),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_297),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_293),
.B2(n_294),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_290),
.B(n_293),
.C(n_297),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_308),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_304),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_306),
.C(n_307),
.Y(n_316)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_329),
.Y(n_309)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_327),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_311),
.B(n_327),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.C(n_323),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_312),
.B(n_324),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_317),
.C(n_318),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_319),
.B1(n_320),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AOI31xp67_ASAP7_75t_L g348 ( 
.A1(n_329),
.A2(n_343),
.A3(n_349),
.B(n_352),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_332),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_332),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_337),
.C(n_338),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_333),
.A2(n_334),
.B1(n_338),
.B2(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_337),
.B(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_338),
.Y(n_346)
);

XNOR2x1_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_347),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_344),
.B(n_347),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);


endmodule