module real_aes_15890_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVx1_ASAP7_75t_L g465 ( .A(n_0), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_1), .A2(n_3), .B1(n_242), .B2(n_243), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_2), .A2(n_21), .B1(n_169), .B2(n_178), .Y(n_186) );
INVx1_ASAP7_75t_L g671 ( .A(n_3), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_4), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g542 ( .A(n_4), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_5), .A2(n_47), .B1(n_85), .B2(n_130), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g108 ( .A1(n_6), .A2(n_10), .B1(n_109), .B2(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g473 ( .A(n_7), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_8), .Y(n_177) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_9), .Y(n_87) );
OAI22xp33_ASAP7_75t_L g550 ( .A1(n_11), .A2(n_17), .B1(n_551), .B2(n_554), .Y(n_550) );
OAI22xp33_ASAP7_75t_L g591 ( .A1(n_11), .A2(n_17), .B1(n_592), .B2(n_595), .Y(n_591) );
INVx1_ASAP7_75t_L g472 ( .A(n_12), .Y(n_472) );
INVx1_ASAP7_75t_L g479 ( .A(n_12), .Y(n_479) );
INVx1_ASAP7_75t_L g578 ( .A(n_13), .Y(n_578) );
OAI211xp5_ASAP7_75t_L g607 ( .A1(n_13), .A2(n_608), .B(n_611), .C(n_615), .Y(n_607) );
INVx1_ASAP7_75t_L g482 ( .A(n_14), .Y(n_482) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_15), .Y(n_658) );
INVx2_ASAP7_75t_L g463 ( .A(n_16), .Y(n_463) );
OAI21x1_ASAP7_75t_L g117 ( .A1(n_18), .A2(n_43), .B(n_118), .Y(n_117) );
XNOR2xp5_ASAP7_75t_L g451 ( .A(n_19), .B(n_452), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_20), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_22), .B(n_90), .Y(n_198) );
INVx4_ASAP7_75t_R g152 ( .A(n_23), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_24), .B(n_169), .Y(n_204) );
INVx1_ASAP7_75t_L g247 ( .A(n_25), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_SL g175 ( .A1(n_26), .A2(n_89), .B(n_109), .C(n_176), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_27), .A2(n_40), .B1(n_109), .B2(n_112), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_28), .A2(n_31), .B1(n_580), .B2(n_582), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_28), .A2(n_31), .B1(n_600), .B2(n_603), .Y(n_599) );
INVx1_ASAP7_75t_L g506 ( .A(n_29), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_30), .Y(n_172) );
BUFx2_ASAP7_75t_L g656 ( .A(n_32), .Y(n_656) );
INVx1_ASAP7_75t_L g572 ( .A(n_33), .Y(n_572) );
INVx2_ASAP7_75t_L g462 ( .A(n_34), .Y(n_462) );
INVx1_ASAP7_75t_L g503 ( .A(n_34), .Y(n_503) );
INVx1_ASAP7_75t_L g201 ( .A(n_35), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_36), .B(n_109), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_37), .Y(n_220) );
INVx2_ASAP7_75t_L g643 ( .A(n_38), .Y(n_643) );
INVx1_ASAP7_75t_L g508 ( .A(n_39), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_41), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_42), .A2(n_71), .B1(n_109), .B2(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g488 ( .A(n_44), .Y(n_488) );
BUFx3_ASAP7_75t_L g666 ( .A(n_45), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_46), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_46), .Y(n_655) );
BUFx3_ASAP7_75t_L g470 ( .A(n_48), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_49), .Y(n_120) );
AND2x4_ASAP7_75t_L g93 ( .A(n_50), .B(n_94), .Y(n_93) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_50), .Y(n_629) );
INVx1_ASAP7_75t_L g118 ( .A(n_51), .Y(n_118) );
INVx1_ASAP7_75t_L g497 ( .A(n_52), .Y(n_497) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_53), .Y(n_515) );
INVx1_ASAP7_75t_L g494 ( .A(n_54), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_55), .A2(n_73), .B1(n_112), .B2(n_240), .Y(n_239) );
AO22x1_ASAP7_75t_L g133 ( .A1(n_56), .A2(n_63), .B1(n_134), .B2(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g94 ( .A(n_57), .Y(n_94) );
AND2x2_ASAP7_75t_L g179 ( .A(n_58), .B(n_180), .Y(n_179) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_59), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_60), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_61), .B(n_130), .Y(n_226) );
BUFx2_ASAP7_75t_L g679 ( .A(n_61), .Y(n_679) );
OAI211xp5_ASAP7_75t_L g560 ( .A1(n_62), .A2(n_561), .B(n_562), .C(n_568), .Y(n_560) );
INVx1_ASAP7_75t_L g622 ( .A(n_62), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_64), .B(n_169), .Y(n_221) );
INVx2_ASAP7_75t_L g90 ( .A(n_65), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_66), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_67), .B(n_180), .Y(n_195) );
INVx1_ASAP7_75t_L g673 ( .A(n_68), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_69), .B(n_116), .Y(n_131) );
BUFx3_ASAP7_75t_L g524 ( .A(n_70), .Y(n_524) );
INVx1_ASAP7_75t_L g557 ( .A(n_70), .Y(n_557) );
INVx1_ASAP7_75t_L g460 ( .A(n_72), .Y(n_460) );
INVx2_ASAP7_75t_L g501 ( .A(n_72), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_74), .B(n_180), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g147 ( .A1(n_75), .A2(n_114), .B(n_130), .C(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g664 ( .A(n_75), .Y(n_664) );
AND2x2_ASAP7_75t_L g156 ( .A(n_76), .B(n_157), .Y(n_156) );
NAND2xp33_ASAP7_75t_L g225 ( .A(n_77), .B(n_153), .Y(n_225) );
INVx1_ASAP7_75t_SL g685 ( .A(n_77), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_95), .B(n_450), .Y(n_78) );
BUFx2_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
NOR2xp33_ASAP7_75t_L g80 ( .A(n_81), .B(n_91), .Y(n_80) );
AO21x2_ASAP7_75t_L g688 ( .A1(n_81), .A2(n_630), .B(n_689), .Y(n_688) );
NAND2xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_88), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_86), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx3_ASAP7_75t_L g109 ( .A(n_87), .Y(n_109) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_87), .Y(n_112) );
INVx1_ASAP7_75t_L g130 ( .A(n_87), .Y(n_130) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_87), .Y(n_135) );
INVx1_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_87), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_87), .Y(n_154) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_87), .Y(n_169) );
INVx1_ASAP7_75t_L g171 ( .A(n_87), .Y(n_171) );
INVx2_ASAP7_75t_L g178 ( .A(n_87), .Y(n_178) );
OAI22x1_ASAP7_75t_L g107 ( .A1(n_88), .A2(n_108), .B1(n_111), .B2(n_113), .Y(n_107) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_88), .A2(n_126), .B1(n_186), .B2(n_187), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_88), .A2(n_113), .B1(n_239), .B2(n_241), .Y(n_238) );
INVx6_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_89), .B(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_89), .A2(n_225), .B(n_226), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_89), .A2(n_125), .B(n_133), .C(n_139), .Y(n_268) );
BUFx8_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g114 ( .A(n_90), .Y(n_114) );
INVx2_ASAP7_75t_L g128 ( .A(n_90), .Y(n_128) );
INVx1_ASAP7_75t_L g174 ( .A(n_90), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_91), .A2(n_147), .B(n_150), .Y(n_146) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AO31x2_ASAP7_75t_L g106 ( .A1(n_92), .A2(n_107), .A3(n_115), .B(n_119), .Y(n_106) );
BUFx10_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
BUFx10_ASAP7_75t_L g189 ( .A(n_93), .Y(n_189) );
INVx1_ASAP7_75t_L g245 ( .A(n_93), .Y(n_245) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_94), .Y(n_631) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
NOR2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_364), .Y(n_97) );
NAND4xp75_ASAP7_75t_L g98 ( .A(n_99), .B(n_269), .C(n_311), .D(n_335), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI211xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_158), .B(n_206), .C(n_248), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g355 ( .A(n_103), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g449 ( .A(n_103), .B(n_386), .Y(n_449) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_122), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g264 ( .A(n_105), .B(n_216), .Y(n_264) );
AND2x2_ASAP7_75t_L g305 ( .A(n_105), .B(n_266), .Y(n_305) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g212 ( .A(n_106), .B(n_142), .Y(n_212) );
OR2x2_ASAP7_75t_L g230 ( .A(n_106), .B(n_142), .Y(n_230) );
INVx2_ASAP7_75t_L g256 ( .A(n_106), .Y(n_256) );
AND2x2_ASAP7_75t_L g286 ( .A(n_106), .B(n_216), .Y(n_286) );
AND2x2_ASAP7_75t_L g315 ( .A(n_106), .B(n_141), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_106), .B(n_267), .Y(n_351) );
INVx4_ASAP7_75t_L g110 ( .A(n_109), .Y(n_110) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_110), .A2(n_220), .B(n_221), .C(n_222), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_112), .B(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g242 ( .A(n_112), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_113), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g121 ( .A(n_116), .Y(n_121) );
OAI21xp33_ASAP7_75t_L g139 ( .A1(n_116), .A2(n_131), .B(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_117), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
INVx2_ASAP7_75t_L g157 ( .A(n_121), .Y(n_157) );
BUFx2_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_121), .B(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_121), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g328 ( .A(n_122), .B(n_257), .Y(n_328) );
INVx2_ASAP7_75t_L g423 ( .A(n_122), .Y(n_423) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_141), .Y(n_122) );
INVx2_ASAP7_75t_L g211 ( .A(n_123), .Y(n_211) );
AND2x4_ASAP7_75t_L g254 ( .A(n_123), .B(n_142), .Y(n_254) );
AOI21x1_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_132), .B(n_138), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B(n_131), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_126), .A2(n_203), .B(n_204), .Y(n_202) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g223 ( .A(n_128), .Y(n_223) );
INVxp67_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
OAI21xp33_ASAP7_75t_SL g197 ( .A1(n_136), .A2(n_198), .B(n_199), .Y(n_197) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_140), .A2(n_166), .B(n_175), .Y(n_165) );
AND2x2_ASAP7_75t_L g413 ( .A(n_141), .B(n_211), .Y(n_413) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g277 ( .A(n_142), .Y(n_277) );
AND2x2_ASAP7_75t_L g334 ( .A(n_142), .B(n_216), .Y(n_334) );
AND2x2_ASAP7_75t_L g349 ( .A(n_142), .B(n_257), .Y(n_349) );
AND2x2_ASAP7_75t_L g371 ( .A(n_142), .B(n_211), .Y(n_371) );
AO21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_146), .B(n_156), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI22xp33_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B1(n_154), .B2(n_155), .Y(n_151) );
INVx2_ASAP7_75t_L g240 ( .A(n_153), .Y(n_240) );
OAI211xp5_ASAP7_75t_SL g418 ( .A1(n_158), .A2(n_419), .B(n_421), .C(n_428), .Y(n_418) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_192), .Y(n_159) );
INVxp67_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OR2x2_ASAP7_75t_L g405 ( .A(n_161), .B(n_341), .Y(n_405) );
OR2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_182), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_162), .B(n_194), .Y(n_304) );
INVxp67_ASAP7_75t_L g318 ( .A(n_162), .Y(n_318) );
AND2x2_ASAP7_75t_L g338 ( .A(n_162), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_162), .B(n_251), .Y(n_345) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g234 ( .A(n_163), .Y(n_234) );
AOI21x1_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_179), .Y(n_163) );
AO31x2_ASAP7_75t_L g237 ( .A1(n_164), .A2(n_238), .A3(n_244), .B(n_246), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_173), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
INVx2_ASAP7_75t_L g243 ( .A(n_171), .Y(n_243) );
BUFx4f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_174), .B(n_201), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
INVx2_ASAP7_75t_L g188 ( .A(n_180), .Y(n_188) );
NOR2x1_ASAP7_75t_L g227 ( .A(n_180), .B(n_228), .Y(n_227) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g205 ( .A(n_181), .B(n_189), .Y(n_205) );
OR2x2_ASAP7_75t_L g279 ( .A(n_182), .B(n_261), .Y(n_279) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OR2x2_ASAP7_75t_L g327 ( .A(n_183), .B(n_234), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_183), .B(n_237), .Y(n_333) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g233 ( .A(n_184), .B(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g302 ( .A(n_184), .B(n_237), .Y(n_302) );
BUFx2_ASAP7_75t_L g309 ( .A(n_184), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_184), .B(n_237), .Y(n_389) );
AO31x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_188), .A3(n_189), .B(n_190), .Y(n_184) );
INVx1_ASAP7_75t_L g228 ( .A(n_189), .Y(n_228) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AND2x4_ASAP7_75t_L g319 ( .A(n_193), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g448 ( .A(n_193), .B(n_233), .Y(n_448) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g251 ( .A(n_194), .Y(n_251) );
AND2x2_ASAP7_75t_L g262 ( .A(n_194), .B(n_237), .Y(n_262) );
AND2x2_ASAP7_75t_L g308 ( .A(n_194), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g341 ( .A(n_194), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_194), .B(n_252), .Y(n_358) );
AND2x2_ASAP7_75t_L g397 ( .A(n_194), .B(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_202), .B(n_205), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_213), .B(n_231), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_208), .A2(n_376), .B1(n_377), .B2(n_379), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_212), .Y(n_208) );
AND2x2_ASAP7_75t_L g373 ( .A(n_209), .B(n_264), .Y(n_373) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g288 ( .A(n_210), .Y(n_288) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g437 ( .A(n_211), .B(n_257), .Y(n_437) );
AND2x2_ASAP7_75t_L g401 ( .A(n_212), .B(n_296), .Y(n_401) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_229), .Y(n_213) );
OR2x2_ASAP7_75t_L g298 ( .A(n_214), .B(n_275), .Y(n_298) );
OR2x2_ASAP7_75t_L g410 ( .A(n_214), .B(n_230), .Y(n_410) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g273 ( .A(n_215), .Y(n_273) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g257 ( .A(n_216), .Y(n_257) );
BUFx3_ASAP7_75t_L g339 ( .A(n_216), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
OAI21x1_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_224), .B(n_227), .Y(n_218) );
INVx2_ASAP7_75t_SL g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g407 ( .A(n_230), .B(n_266), .Y(n_407) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
AND2x2_ASAP7_75t_L g249 ( .A(n_233), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g290 ( .A(n_233), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g427 ( .A(n_233), .Y(n_427) );
INVx1_ASAP7_75t_L g446 ( .A(n_233), .Y(n_446) );
INVx2_ASAP7_75t_L g261 ( .A(n_234), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_234), .B(n_237), .Y(n_310) );
INVx1_ASAP7_75t_L g374 ( .A(n_235), .Y(n_374) );
BUFx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g435 ( .A(n_236), .Y(n_435) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g252 ( .A(n_237), .Y(n_252) );
INVx1_ASAP7_75t_L g342 ( .A(n_237), .Y(n_342) );
INVx2_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_253), .B1(n_258), .B2(n_263), .Y(n_248) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g291 ( .A(n_251), .Y(n_291) );
AND2x2_ASAP7_75t_L g293 ( .A(n_251), .B(n_278), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_251), .B(n_261), .Y(n_353) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx3_ASAP7_75t_L g284 ( .A(n_254), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_254), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g378 ( .A(n_254), .B(n_362), .Y(n_378) );
INVx1_ASAP7_75t_L g282 ( .A(n_255), .Y(n_282) );
AOI222xp33_ASAP7_75t_L g292 ( .A1(n_255), .A2(n_293), .B1(n_294), .B2(n_299), .C1(n_305), .C2(n_306), .Y(n_292) );
OAI21xp33_ASAP7_75t_SL g322 ( .A1(n_255), .A2(n_323), .B(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g346 ( .A(n_255), .B(n_265), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_255), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
OR2x2_ASAP7_75t_L g275 ( .A(n_256), .B(n_267), .Y(n_275) );
INVx1_ASAP7_75t_L g363 ( .A(n_256), .Y(n_363) );
BUFx2_ASAP7_75t_L g297 ( .A(n_257), .Y(n_297) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_262), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_260), .B(n_301), .Y(n_330) );
OR2x2_ASAP7_75t_L g442 ( .A(n_260), .B(n_302), .Y(n_442) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g325 ( .A(n_262), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g440 ( .A(n_262), .Y(n_440) );
OAI31xp33_ASAP7_75t_L g421 ( .A1(n_263), .A2(n_422), .A3(n_424), .B(n_425), .Y(n_421) );
AND2x4_ASAP7_75t_SL g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_264), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_292), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_278), .B(n_280), .Y(n_270) );
NOR2x1_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x6_ASAP7_75t_L g391 ( .A(n_273), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g323 ( .A(n_276), .Y(n_323) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g414 ( .A(n_277), .B(n_351), .Y(n_414) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_279), .A2(n_368), .B1(n_370), .B2(n_372), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g428 ( .A1(n_279), .A2(n_340), .B(n_402), .C(n_429), .Y(n_428) );
AOI21xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_285), .B(n_289), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND4xp25_ASAP7_75t_L g381 ( .A(n_284), .B(n_382), .C(n_383), .D(n_385), .Y(n_381) );
NAND2x1_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_286), .B(n_288), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_286), .B(n_371), .Y(n_394) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g360 ( .A(n_291), .B(n_320), .Y(n_360) );
NAND2xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_298), .A2(n_442), .B1(n_443), .B2(n_445), .Y(n_441) );
AOI221x1_ASAP7_75t_L g380 ( .A1(n_299), .A2(n_381), .B1(n_387), .B2(n_390), .C(n_393), .Y(n_380) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g320 ( .A(n_302), .Y(n_320) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g332 ( .A(n_304), .B(n_333), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g395 ( .A(n_305), .B(n_386), .Y(n_395) );
O2A1O1Ixp5_ASAP7_75t_L g408 ( .A1(n_306), .A2(n_390), .B(n_409), .C(n_411), .Y(n_408) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx2_ASAP7_75t_L g357 ( .A(n_309), .Y(n_357) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_321), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_313), .A2(n_331), .B1(n_401), .B2(n_402), .C(n_404), .Y(n_400) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g337 ( .A(n_315), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_315), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g436 ( .A(n_315), .B(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
NAND2x1_ASAP7_75t_L g415 ( .A(n_318), .B(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g439 ( .A(n_318), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g379 ( .A(n_319), .Y(n_379) );
AOI222xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_325), .B1(n_328), .B2(n_329), .C1(n_331), .C2(n_334), .Y(n_321) );
INVx1_ASAP7_75t_L g406 ( .A(n_325), .Y(n_406) );
INVx1_ASAP7_75t_L g369 ( .A(n_326), .Y(n_369) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g403 ( .A(n_327), .Y(n_403) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g344 ( .A(n_333), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g398 ( .A(n_333), .Y(n_398) );
AND2x2_ASAP7_75t_L g361 ( .A(n_334), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_354), .Y(n_335) );
AOI222xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_340), .B1(n_343), .B2(n_346), .C1(n_347), .C2(n_352), .Y(n_336) );
INVx3_ASAP7_75t_L g386 ( .A(n_339), .Y(n_386) );
BUFx2_ASAP7_75t_L g444 ( .A(n_339), .Y(n_444) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g416 ( .A(n_341), .Y(n_416) );
OR2x2_ASAP7_75t_L g426 ( .A(n_341), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx2_ASAP7_75t_SL g384 ( .A(n_349), .Y(n_384) );
AND2x2_ASAP7_75t_L g429 ( .A(n_350), .B(n_386), .Y(n_429) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_351), .Y(n_382) );
INVxp67_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g388 ( .A(n_353), .B(n_389), .Y(n_388) );
NOR2x1_ASAP7_75t_L g354 ( .A(n_355), .B(n_359), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
OR2x2_ASAP7_75t_L g445 ( .A(n_358), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g376 ( .A(n_360), .Y(n_376) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g383 ( .A(n_363), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g433 ( .A(n_363), .Y(n_433) );
NAND4xp75_ASAP7_75t_L g364 ( .A(n_365), .B(n_399), .C(n_417), .D(n_430), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_380), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_374), .B(n_375), .Y(n_366) );
INVxp33_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_369), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g392 ( .A(n_371), .Y(n_392) );
AND2x2_ASAP7_75t_L g432 ( .A(n_371), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g402 ( .A(n_374), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g420 ( .A(n_385), .Y(n_420) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI22xp33_ASAP7_75t_SL g411 ( .A1(n_388), .A2(n_412), .B1(n_414), .B2(n_415), .Y(n_411) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI21xp33_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_395), .B(n_396), .Y(n_393) );
INVx1_ASAP7_75t_L g424 ( .A(n_395), .Y(n_424) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_408), .Y(n_399) );
AOI21xp5_ASAP7_75t_SL g404 ( .A1(n_405), .A2(n_406), .B(n_407), .Y(n_404) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_447), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B1(n_436), .B2(n_438), .C(n_441), .Y(n_431) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B1(n_628), .B2(n_632), .C(n_680), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_452), .A2(n_681), .B1(n_684), .B2(n_686), .Y(n_680) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND3x1_ASAP7_75t_L g453 ( .A(n_454), .B(n_549), .C(n_590), .Y(n_453) );
NOR2xp33_ASAP7_75t_SL g454 ( .A(n_455), .B(n_511), .Y(n_454) );
OAI33xp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_464), .A3(n_481), .B1(n_493), .B2(n_499), .B3(n_505), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_461), .Y(n_457) );
AND2x2_ASAP7_75t_SL g540 ( .A(n_458), .B(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_458), .Y(n_627) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx2_ASAP7_75t_L g589 ( .A(n_459), .Y(n_589) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx2_ASAP7_75t_L g648 ( .A(n_461), .Y(n_648) );
NAND2xp33_ASAP7_75t_SL g461 ( .A(n_462), .B(n_463), .Y(n_461) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_462), .Y(n_625) );
INVx1_ASAP7_75t_L g642 ( .A(n_462), .Y(n_642) );
INVx3_ASAP7_75t_L g504 ( .A(n_463), .Y(n_504) );
BUFx3_ASAP7_75t_L g618 ( .A(n_463), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B1(n_473), .B2(n_474), .Y(n_464) );
OAI22xp33_ASAP7_75t_L g525 ( .A1(n_465), .A2(n_506), .B1(n_526), .B2(n_530), .Y(n_525) );
BUFx4f_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx3_ASAP7_75t_L g507 ( .A(n_469), .Y(n_507) );
OR2x4_ASAP7_75t_L g594 ( .A(n_469), .B(n_504), .Y(n_594) );
OR2x4_ASAP7_75t_L g602 ( .A(n_469), .B(n_597), .Y(n_602) );
OR2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_470), .Y(n_480) );
INVx2_ASAP7_75t_L g487 ( .A(n_470), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_470), .B(n_479), .Y(n_492) );
AND2x4_ASAP7_75t_L g613 ( .A(n_470), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVxp67_ASAP7_75t_L g486 ( .A(n_472), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_473), .A2(n_508), .B1(n_544), .B2(n_547), .Y(n_543) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g510 ( .A(n_476), .Y(n_510) );
BUFx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx3_ASAP7_75t_L g610 ( .A(n_477), .Y(n_610) );
NAND2x1p5_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
BUFx2_ASAP7_75t_L g621 ( .A(n_478), .Y(n_621) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g614 ( .A(n_479), .Y(n_614) );
BUFx2_ASAP7_75t_L g619 ( .A(n_480), .Y(n_619) );
INVx2_ASAP7_75t_L g640 ( .A(n_480), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B1(n_488), .B2(n_489), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_482), .A2(n_494), .B1(n_513), .B2(n_518), .Y(n_512) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx8_ASAP7_75t_L g496 ( .A(n_485), .Y(n_496) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_485), .Y(n_598) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_488), .A2(n_497), .B1(n_536), .B2(n_538), .Y(n_535) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx3_ASAP7_75t_L g498 ( .A(n_490), .Y(n_498) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx2_ASAP7_75t_L g606 ( .A(n_492), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_497), .B2(n_498), .Y(n_493) );
INVx2_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
AND2x4_ASAP7_75t_L g522 ( .A(n_500), .B(n_523), .Y(n_522) );
BUFx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2x1p5_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g597 ( .A(n_504), .Y(n_597) );
OR2x6_ASAP7_75t_L g605 ( .A(n_504), .B(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g612 ( .A(n_504), .B(n_613), .Y(n_612) );
AND2x4_ASAP7_75t_L g641 ( .A(n_504), .B(n_642), .Y(n_641) );
OAI22xp33_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B1(n_508), .B2(n_509), .Y(n_505) );
INVxp67_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
OAI33xp33_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_521), .A3(n_525), .B1(n_535), .B2(n_539), .B3(n_543), .Y(n_511) );
BUFx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g546 ( .A(n_514), .Y(n_546) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
NAND2x1_ASAP7_75t_L g520 ( .A(n_515), .B(n_517), .Y(n_520) );
OR2x2_ASAP7_75t_L g529 ( .A(n_515), .B(n_517), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_515), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g559 ( .A(n_515), .Y(n_559) );
AND2x2_ASAP7_75t_L g567 ( .A(n_515), .B(n_517), .Y(n_567) );
BUFx2_ASAP7_75t_L g571 ( .A(n_515), .Y(n_571) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g534 ( .A(n_517), .Y(n_534) );
AND2x2_ASAP7_75t_L g558 ( .A(n_517), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g577 ( .A(n_517), .Y(n_577) );
BUFx4f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx4_ASAP7_75t_L g548 ( .A(n_519), .Y(n_548) );
BUFx4f_ASAP7_75t_L g561 ( .A(n_519), .Y(n_561) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x4_ASAP7_75t_L g541 ( .A(n_524), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g553 ( .A(n_524), .Y(n_553) );
BUFx2_ASAP7_75t_L g570 ( .A(n_524), .Y(n_570) );
AND2x4_ASAP7_75t_L g575 ( .A(n_524), .B(n_576), .Y(n_575) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x6_ASAP7_75t_L g551 ( .A(n_527), .B(n_552), .Y(n_551) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g537 ( .A(n_528), .Y(n_537) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx8_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g538 ( .A(n_532), .Y(n_538) );
OR2x2_ASAP7_75t_L g584 ( .A(n_532), .B(n_570), .Y(n_584) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx4f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x6_ASAP7_75t_L g581 ( .A(n_537), .B(n_556), .Y(n_581) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g587 ( .A(n_542), .Y(n_587) );
INVx4_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx4_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OAI31xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_560), .A3(n_579), .B(n_585), .Y(n_549) );
INVxp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g564 ( .A(n_553), .Y(n_564) );
CKINVDCx16_ASAP7_75t_R g554 ( .A(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_572), .B1(n_573), .B2(n_578), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_572), .A2(n_616), .B1(n_620), .B2(n_622), .Y(n_615) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OAI31xp33_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_599), .A3(n_607), .B(n_623), .Y(n_590) );
INVx2_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
CKINVDCx8_ASAP7_75t_R g611 ( .A(n_612), .Y(n_611) );
AND2x4_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
AND2x4_ASAP7_75t_L g620 ( .A(n_617), .B(n_621), .Y(n_620) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g650 ( .A(n_629), .Y(n_650) );
BUFx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_631), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g689 ( .A(n_631), .B(n_650), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_651), .B1(n_675), .B2(n_679), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx12f_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx3_ASAP7_75t_L g682 ( .A(n_635), .Y(n_682) );
BUFx8_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI211xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_643), .B(n_644), .C(n_649), .Y(n_636) );
AND2x2_ASAP7_75t_L g678 ( .A(n_637), .B(n_644), .Y(n_678) );
INVx4_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x6_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_639), .B(n_645), .C(n_648), .Y(n_644) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx3_ASAP7_75t_L g647 ( .A(n_643), .Y(n_647) );
INVx2_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
BUFx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g677 ( .A(n_649), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_651), .A2(n_679), .B1(n_682), .B2(n_683), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_661), .B2(n_662), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_653) );
INVx1_ASAP7_75t_L g659 ( .A(n_654), .Y(n_659) );
INVx1_ASAP7_75t_L g657 ( .A(n_656), .Y(n_657) );
INVx2_ASAP7_75t_L g660 ( .A(n_658), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_668), .B1(n_669), .B2(n_674), .Y(n_662) );
INVx1_ASAP7_75t_L g674 ( .A(n_663), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_666), .B2(n_667), .Y(n_663) );
INVx1_ASAP7_75t_L g667 ( .A(n_664), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_672), .B2(n_673), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
BUFx2_ASAP7_75t_L g683 ( .A(n_676), .Y(n_683) );
OR2x6_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_687), .Y(n_686) );
CKINVDCx16_ASAP7_75t_R g687 ( .A(n_688), .Y(n_687) );
endmodule