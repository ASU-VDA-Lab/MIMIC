module fake_jpeg_22148_n_38 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_20),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_1),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_21),
.B(n_23),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_2),
.B1(n_3),
.B2(n_11),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_8),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_12),
.A2(n_10),
.B1(n_14),
.B2(n_16),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_10),
.A2(n_11),
.B1(n_9),
.B2(n_12),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_20),
.B(n_21),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_18),
.B1(n_25),
.B2(n_28),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_22),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_30),
.C(n_31),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_36),
.Y(n_37)
);

BUFx24_ASAP7_75t_SL g38 ( 
.A(n_37),
.Y(n_38)
);


endmodule