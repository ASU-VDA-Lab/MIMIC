module fake_jpeg_22673_n_75 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_75);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_75;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_22;
wire n_47;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_59;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_74;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_10),
.Y(n_23)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_0),
.B(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_7),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_11),
.B(n_12),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_42),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_2),
.Y(n_43)
);

O2A1O1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_21),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_44)
);

A2O1A1O1Ixp25_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_46),
.B(n_50),
.C(n_51),
.D(n_26),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_6),
.B1(n_29),
.B2(n_36),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_20),
.B(n_22),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_48),
.B(n_49),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_20),
.B(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_36),
.Y(n_51)
);

OAI21x1_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_54),
.B(n_46),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_40),
.B1(n_37),
.B2(n_44),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_38),
.B(n_43),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_61),
.C(n_64),
.Y(n_67)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_63),
.Y(n_66)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_57),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_67),
.A2(n_57),
.B(n_55),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_60),
.C(n_52),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_72),
.C(n_46),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_68),
.C(n_39),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_54),
.B1(n_59),
.B2(n_71),
.Y(n_75)
);


endmodule