module fake_jpeg_2440_n_26 (n_3, n_2, n_1, n_0, n_4, n_26);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_26;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_0),
.Y(n_5)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_1),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_12),
.C(n_13),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_2),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_10),
.A2(n_7),
.B1(n_9),
.B2(n_8),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_17),
.B1(n_5),
.B2(n_2),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_7),
.B1(n_5),
.B2(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_19),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_4),
.C(n_16),
.Y(n_20)
);

AOI21x1_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_20),
.B(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_16),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_24),
.C(n_22),
.Y(n_26)
);


endmodule