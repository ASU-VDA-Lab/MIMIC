module real_jpeg_850_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_3),
.A2(n_28),
.B1(n_38),
.B2(n_39),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_4),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_4),
.A2(n_34),
.B1(n_62),
.B2(n_63),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_4),
.A2(n_34),
.B1(n_57),
.B2(n_58),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_4),
.B(n_55),
.C(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_4),
.B(n_54),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_4),
.B(n_39),
.C(n_74),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_4),
.B(n_30),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_4),
.B(n_42),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_25),
.C(n_43),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_4),
.B(n_99),
.Y(n_196)
);

BUFx4f_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_6),
.A2(n_48),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_48),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_6),
.A2(n_48),
.B1(n_57),
.B2(n_58),
.Y(n_97)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_125),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_124),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_101),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_17),
.B(n_101),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_78),
.C(n_86),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_18),
.A2(n_19),
.B1(n_78),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_49),
.B2(n_50),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_20),
.B(n_51),
.C(n_71),
.Y(n_102)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_35),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_22),
.A2(n_35),
.B1(n_36),
.B2(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_22),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_29),
.B(n_31),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_23),
.A2(n_29),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_30),
.Y(n_32)
);

AO22x1_ASAP7_75t_SL g42 ( 
.A1(n_24),
.A2(n_25),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_25),
.B(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_29),
.B(n_81),
.Y(n_116)
);

OA21x2_ASAP7_75t_L g148 ( 
.A1(n_29),
.A2(n_31),
.B(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_33),
.B(n_116),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_35),
.A2(n_36),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_35),
.B(n_190),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_35),
.A2(n_36),
.B1(n_109),
.B2(n_111),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_35),
.B(n_109),
.C(n_204),
.Y(n_210)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_46),
.B2(n_47),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_37),
.A2(n_41),
.B1(n_46),
.B2(n_47),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_37),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_37),
.A2(n_41),
.B(n_46),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_45)
);

AOI22x1_ASAP7_75t_L g76 ( 
.A1(n_38),
.A2(n_39),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_39),
.B(n_189),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_46),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_70),
.B2(n_71),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_51),
.B(n_109),
.C(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_51),
.A2(n_52),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OA21x2_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_61),
.B(n_66),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_55),
.B(n_62),
.C(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_67),
.B1(n_68),
.B2(n_88),
.Y(n_87)
);

AO22x1_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_62),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_58),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_58),
.B(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B(n_77),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_84),
.A2(n_85),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_84),
.A2(n_85),
.B1(n_169),
.B2(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_85),
.B(n_164),
.C(n_169),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_85),
.B(n_94),
.C(n_196),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.C(n_96),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_87),
.A2(n_96),
.B1(n_112),
.B2(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_89),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_93),
.A2(n_94),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_94),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_94),
.B(n_184),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_95),
.Y(n_149)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_147),
.C(n_148),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_96),
.A2(n_131),
.B1(n_165),
.B2(n_168),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

AO21x1_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_99),
.B(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_113),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_111),
.B1(n_139),
.B2(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_117),
.B1(n_118),
.B2(n_123),
.Y(n_113)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

OAI211xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_150),
.B(n_156),
.C(n_157),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_140),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_140),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_135),
.C(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.C(n_146),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_148),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_158),
.C(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_153),
.Y(n_156)
);

OAI21x1_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_175),
.B(n_212),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_163),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

NOR2xp67_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_187),
.Y(n_191)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_206),
.B(n_211),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_200),
.B(n_205),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_192),
.B(n_199),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_186),
.B(n_191),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_183),
.B(n_185),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_188),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_198),
.Y(n_199)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_202),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_210),
.Y(n_211)
);


endmodule