module fake_jpeg_10809_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_66),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_0),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_62),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_57),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_86),
.Y(n_93)
);

CKINVDCx6p67_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_49),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_56),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_63),
.B1(n_44),
.B2(n_55),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_88),
.B1(n_101),
.B2(n_100),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_44),
.B1(n_55),
.B2(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_98),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_67),
.B1(n_60),
.B2(n_61),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_53),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_59),
.B1(n_48),
.B2(n_45),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_2),
.B(n_3),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_80),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_4),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_23),
.B1(n_42),
.B2(n_41),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_1),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_21),
.Y(n_104)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_28),
.A3(n_39),
.B1(n_38),
.B2(n_36),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_76),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_108),
.C(n_109),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_19),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_25),
.C(n_40),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_4),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_5),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_121),
.B1(n_11),
.B2(n_12),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_6),
.Y(n_116)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_120),
.B1(n_122),
.B2(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_8),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_119),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_10),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_104),
.C(n_33),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_108),
.C(n_112),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_131),
.A2(n_132),
.B(n_107),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_18),
.B1(n_26),
.B2(n_27),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_118),
.Y(n_133)
);

NOR4xp25_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.C(n_135),
.D(n_43),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_12),
.B1(n_34),
.B2(n_35),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_110),
.B(n_123),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_139),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_142),
.A3(n_141),
.B1(n_138),
.B2(n_129),
.C1(n_140),
.C2(n_127),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_128),
.B(n_124),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_143),
.C(n_130),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_132),
.Y(n_150)
);


endmodule