module fake_jpeg_17808_n_356 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_356);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_7),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_41),
.B(n_11),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_49),
.Y(n_69)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_47),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_21),
.A2(n_7),
.B1(n_12),
.B2(n_2),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_20),
.B1(n_16),
.B2(n_24),
.Y(n_91)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_57),
.Y(n_74)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_65),
.Y(n_79)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_30),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_37),
.B1(n_18),
.B2(n_30),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_71),
.A2(n_76),
.B1(n_95),
.B2(n_99),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_85),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_75),
.A2(n_93),
.B(n_89),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_21),
.B1(n_20),
.B2(n_24),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_19),
.B(n_26),
.C(n_28),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_77),
.A2(n_0),
.B(n_1),
.C(n_72),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_22),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_81),
.B(n_88),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_22),
.Y(n_88)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_91),
.A2(n_0),
.B(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_33),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_92),
.B(n_115),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_33),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_98),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_28),
.B1(n_26),
.B2(n_19),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_31),
.B1(n_9),
.B2(n_2),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_96),
.A2(n_101),
.B1(n_111),
.B2(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_31),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_31),
.B1(n_35),
.B2(n_15),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_35),
.B1(n_15),
.B2(n_14),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_105),
.B1(n_118),
.B2(n_12),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_38),
.A2(n_8),
.B1(n_13),
.B2(n_2),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_43),
.A2(n_35),
.B1(n_15),
.B2(n_14),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_8),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_8),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_SL g108 ( 
.A(n_50),
.Y(n_108)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_46),
.A2(n_9),
.B1(n_13),
.B2(n_3),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_59),
.A2(n_9),
.B1(n_12),
.B2(n_4),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_57),
.B(n_10),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_0),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_55),
.A2(n_10),
.B1(n_12),
.B2(n_5),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_114),
.A2(n_110),
.B1(n_116),
.B2(n_68),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_115),
.B(n_113),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_63),
.B(n_11),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_117),
.A2(n_15),
.B(n_6),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_56),
.A2(n_60),
.B1(n_62),
.B2(n_47),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_77),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_119),
.B(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_61),
.B1(n_48),
.B2(n_42),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_122),
.A2(n_125),
.B1(n_132),
.B2(n_145),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_15),
.B(n_35),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_123),
.A2(n_138),
.B(n_162),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_127),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_61),
.B1(n_48),
.B2(n_42),
.Y(n_125)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_70),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_79),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_134),
.Y(n_183)
);

AOI22x1_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_48),
.B1(n_61),
.B2(n_6),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_7),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_141),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_142),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_72),
.A2(n_0),
.B(n_1),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_93),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_74),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_152),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_144),
.A2(n_165),
.B(n_127),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_102),
.A2(n_116),
.B1(n_82),
.B2(n_103),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_100),
.A2(n_102),
.B1(n_87),
.B2(n_70),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_124),
.B1(n_132),
.B2(n_121),
.Y(n_182)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_73),
.A2(n_110),
.B1(n_89),
.B2(n_68),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_126),
.B(n_133),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_73),
.A2(n_110),
.B1(n_90),
.B2(n_78),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_90),
.A2(n_78),
.B1(n_82),
.B2(n_103),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_83),
.A2(n_84),
.B1(n_109),
.B2(n_87),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_159),
.A2(n_83),
.B1(n_84),
.B2(n_104),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_109),
.A2(n_76),
.B1(n_93),
.B2(n_107),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_160),
.A2(n_166),
.B1(n_164),
.B2(n_129),
.Y(n_191)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_162),
.B(n_163),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_163),
.B(n_131),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_106),
.B(n_74),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_69),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_85),
.B(n_69),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_169),
.B(n_206),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_188),
.B1(n_135),
.B2(n_152),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_80),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_179),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_104),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_182),
.A2(n_186),
.B1(n_187),
.B2(n_191),
.Y(n_212)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_202),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_119),
.A2(n_144),
.B1(n_146),
.B2(n_120),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_148),
.B1(n_132),
.B2(n_143),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_140),
.A2(n_130),
.B1(n_161),
.B2(n_141),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

HAxp5_ASAP7_75t_SL g208 ( 
.A(n_190),
.B(n_122),
.CON(n_208),
.SN(n_208)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_137),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_204),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_196),
.A2(n_197),
.B(n_200),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_126),
.A2(n_138),
.B(n_133),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_122),
.A2(n_165),
.B(n_125),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_160),
.B(n_142),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_165),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_192),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_207),
.B(n_204),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_208),
.A2(n_242),
.B(n_243),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_201),
.A2(n_151),
.B1(n_122),
.B2(n_160),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_209),
.A2(n_210),
.B1(n_214),
.B2(n_240),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_219),
.B(n_223),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_171),
.A2(n_151),
.B1(n_160),
.B2(n_145),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_135),
.B(n_197),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_203),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_221),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_193),
.A2(n_135),
.B(n_200),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_171),
.A2(n_181),
.B1(n_198),
.B2(n_172),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_226),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_174),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_227),
.B(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_174),
.B(n_169),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_229),
.B(n_237),
.Y(n_257)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_183),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_235),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_239),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_206),
.B(n_178),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_167),
.B(n_170),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_238),
.Y(n_252)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_181),
.A2(n_182),
.B1(n_187),
.B2(n_171),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_241),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_176),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_177),
.B(n_207),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_250),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g254 ( 
.A(n_224),
.B(n_179),
.CI(n_186),
.CON(n_254),
.SN(n_254)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_254),
.B(n_268),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_227),
.A2(n_190),
.B(n_184),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_255),
.A2(n_261),
.B(n_262),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_216),
.B(n_195),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_260),
.C(n_270),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_184),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_225),
.A2(n_167),
.B1(n_170),
.B2(n_180),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_219),
.A2(n_177),
.B(n_176),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_180),
.B1(n_185),
.B2(n_194),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_272),
.B1(n_210),
.B2(n_240),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_224),
.A2(n_219),
.B(n_212),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_266),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_212),
.A2(n_223),
.B(n_213),
.Y(n_266)
);

NAND3xp33_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_235),
.C(n_226),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_232),
.Y(n_269)
);

OA22x2_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_271),
.B1(n_242),
.B2(n_221),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_223),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_236),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_240),
.A2(n_225),
.B1(n_209),
.B2(n_214),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_278),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_277),
.A2(n_291),
.B1(n_297),
.B2(n_261),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_228),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_218),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_280),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_218),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_234),
.C(n_229),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_282),
.C(n_287),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_270),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_237),
.C(n_213),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_243),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_289),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_273),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_249),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_256),
.A2(n_240),
.B1(n_238),
.B2(n_231),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_220),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_288),
.Y(n_301)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

OAI321xp33_ASAP7_75t_L g295 ( 
.A1(n_257),
.A2(n_211),
.A3(n_222),
.B1(n_215),
.B2(n_239),
.C(n_241),
.Y(n_295)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_258),
.A3(n_249),
.B1(n_255),
.B2(n_253),
.C1(n_254),
.C2(n_244),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_215),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_298),
.C(n_269),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_246),
.A2(n_217),
.B1(n_230),
.B2(n_272),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_244),
.B(n_217),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_246),
.B1(n_263),
.B2(n_266),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_300),
.B(n_301),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_303),
.Y(n_322)
);

NAND3xp33_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_279),
.C(n_278),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_277),
.A2(n_254),
.B1(n_262),
.B2(n_258),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_313),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_253),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_316),
.C(n_287),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_282),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_297),
.A2(n_271),
.B1(n_245),
.B2(n_251),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_276),
.A2(n_245),
.B1(n_251),
.B2(n_267),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_289),
.Y(n_327)
);

NAND2x1_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_264),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_274),
.B(n_285),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_275),
.B(n_264),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_321),
.Y(n_334)
);

OAI31xp33_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_283),
.A3(n_292),
.B(n_280),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_319),
.A2(n_325),
.B(n_311),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_330),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_296),
.C(n_298),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_326),
.C(n_329),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_281),
.C(n_276),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_327),
.B(n_313),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_328),
.B(n_305),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_283),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_309),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_301),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_332),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_333),
.A2(n_336),
.B1(n_308),
.B2(n_300),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_309),
.Y(n_337)
);

OAI221xp5_ASAP7_75t_L g344 ( 
.A1(n_337),
.A2(n_338),
.B1(n_339),
.B2(n_284),
.C(n_286),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_322),
.B(n_318),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_324),
.B(n_299),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_341),
.B(n_345),
.Y(n_349)
);

NAND3xp33_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_304),
.C(n_319),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_342),
.B(n_344),
.Y(n_347)
);

OAI221xp5_ASAP7_75t_L g345 ( 
.A1(n_333),
.A2(n_291),
.B1(n_294),
.B2(n_321),
.C(n_326),
.Y(n_345)
);

NAND4xp25_ASAP7_75t_SL g346 ( 
.A(n_335),
.B(n_289),
.C(n_302),
.D(n_307),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_346),
.B(n_329),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_334),
.C(n_337),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_SL g351 ( 
.A(n_348),
.B(n_334),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_350),
.A2(n_307),
.B(n_335),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_351),
.B(n_352),
.Y(n_353)
);

OAI321xp33_ASAP7_75t_L g354 ( 
.A1(n_353),
.A2(n_347),
.A3(n_349),
.B1(n_323),
.B2(n_348),
.C(n_340),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_340),
.C(n_317),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_230),
.Y(n_356)
);


endmodule