module fake_jpeg_14328_n_132 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_16),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_37),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_18),
.A2(n_1),
.B(n_2),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_19),
.C(n_15),
.Y(n_60)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_6),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_22),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_23),
.B1(n_26),
.B2(n_25),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_64),
.B1(n_45),
.B2(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_60),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_30),
.A2(n_24),
.B1(n_25),
.B2(n_20),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_40),
.B1(n_5),
.B2(n_3),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_26),
.B1(n_23),
.B2(n_18),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_61),
.B1(n_62),
.B2(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_12),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_56),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_27),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_19),
.B1(n_15),
.B2(n_14),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_28),
.A2(n_14),
.B1(n_27),
.B2(n_4),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_72),
.B(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_75),
.Y(n_91)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_9),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_48),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_51),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_54),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_63),
.B1(n_68),
.B2(n_46),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_63),
.B1(n_68),
.B2(n_46),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_67),
.C(n_85),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_65),
.B(n_54),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_100),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_65),
.B(n_67),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_87),
.B(n_91),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_98),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_100),
.B1(n_88),
.B2(n_96),
.Y(n_105)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_89),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_75),
.C(n_71),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_76),
.B(n_73),
.C(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_84),
.B1(n_83),
.B2(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_109),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_107),
.B(n_110),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_97),
.B1(n_99),
.B2(n_94),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_92),
.B(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_111),
.B(n_113),
.Y(n_119)
);

OA21x2_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_88),
.B(n_105),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_114),
.Y(n_121)
);

AO221x1_ASAP7_75t_L g118 ( 
.A1(n_115),
.A2(n_102),
.B1(n_110),
.B2(n_104),
.C(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_119),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_112),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_120),
.B(n_121),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_115),
.B(n_116),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_116),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_120),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_121),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_124),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_128),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_122),
.Y(n_132)
);


endmodule