module fake_jpeg_22296_n_111 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_27),
.Y(n_39)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_30),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_0),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_41),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_16),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2x1_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_14),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_19),
.B1(n_13),
.B2(n_17),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_19),
.B1(n_13),
.B2(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_24),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_56),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_35),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_31),
.B1(n_27),
.B2(n_26),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_13),
.B1(n_32),
.B2(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_16),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_55),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_16),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

AND2x6_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_0),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_48),
.Y(n_66)
);

AOI22x1_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_43),
.B1(n_32),
.B2(n_37),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_50),
.B1(n_37),
.B2(n_55),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_71),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_52),
.B1(n_58),
.B2(n_23),
.Y(n_78)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_38),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_78),
.B1(n_64),
.B2(n_67),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_53),
.B(n_59),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_52),
.C(n_51),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_80),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_24),
.C(n_23),
.Y(n_80)
);

XNOR2x1_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_16),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_60),
.B(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_75),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_88),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_85),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_21),
.B(n_18),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_75),
.C(n_62),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_88),
.C(n_85),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_94),
.B(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_97),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_72),
.Y(n_97)
);

AOI322xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_93),
.A3(n_72),
.B1(n_15),
.B2(n_36),
.C1(n_8),
.C2(n_9),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

AO21x1_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_15),
.B(n_10),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_102),
.B(n_98),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_105),
.B(n_106),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_18),
.C(n_15),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_5),
.C(n_2),
.Y(n_106)
);

AOI322xp5_ASAP7_75t_L g108 ( 
.A1(n_104),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.C1(n_36),
.C2(n_102),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_108),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_107),
.C(n_36),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_1),
.Y(n_111)
);


endmodule