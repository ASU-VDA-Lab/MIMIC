module fake_netlist_1_7336_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
CKINVDCx16_ASAP7_75t_R g11 ( .A(n_6), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_7), .Y(n_13) );
INVx1_ASAP7_75t_SL g14 ( .A(n_10), .Y(n_14) );
INVx2_ASAP7_75t_SL g15 ( .A(n_9), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_3), .Y(n_16) );
CKINVDCx16_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
O2A1O1Ixp5_ASAP7_75t_L g19 ( .A1(n_15), .A2(n_0), .B(n_1), .C(n_2), .Y(n_19) );
NOR2x1_ASAP7_75t_R g20 ( .A(n_16), .B(n_0), .Y(n_20) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
OAI21xp33_ASAP7_75t_SL g22 ( .A1(n_15), .A2(n_1), .B(n_2), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_21), .B(n_13), .Y(n_23) );
NOR2xp33_ASAP7_75t_R g24 ( .A(n_18), .B(n_17), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_18), .B(n_11), .Y(n_25) );
CKINVDCx16_ASAP7_75t_R g26 ( .A(n_20), .Y(n_26) );
NOR4xp25_ASAP7_75t_SL g27 ( .A(n_26), .B(n_13), .C(n_20), .D(n_22), .Y(n_27) );
NAND2xp67_ASAP7_75t_L g28 ( .A(n_25), .B(n_19), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_23), .B(n_14), .Y(n_29) );
OAI22xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_27), .B1(n_28), .B2(n_24), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
INVx1_ASAP7_75t_SL g32 ( .A(n_31), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_3), .Y(n_33) );
CKINVDCx20_ASAP7_75t_R g34 ( .A(n_33), .Y(n_34) );
BUFx2_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
AOI22xp5_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_5), .B1(n_12), .B2(n_34), .Y(n_36) );
endmodule