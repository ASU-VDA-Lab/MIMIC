module fake_ariane_1464_n_2065 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_439, n_222, n_478, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_503, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_384, n_468, n_61, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_496, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_2065);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_439;
input n_222;
input n_478;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_503;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_384;
input n_468;
input n_61;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;

output n_2065;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_1383;
wire n_603;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_813;
wire n_1985;
wire n_995;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_1751;
wire n_533;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_650;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_1913;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_552;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_1467;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_1156;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1854;
wire n_666;
wire n_1747;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_519;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_937;
wire n_1474;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_523;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_849;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_242),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_188),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_52),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_53),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_387),
.Y(n_514)
);

CKINVDCx14_ASAP7_75t_R g515 ( 
.A(n_183),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_310),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_495),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_497),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_129),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_265),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_65),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_298),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_352),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_21),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_404),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_459),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_315),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_109),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_108),
.Y(n_529)
);

BUFx10_ASAP7_75t_L g530 ( 
.A(n_259),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_149),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_122),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_8),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_500),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_181),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_77),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_337),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_471),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_446),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_508),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_144),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_283),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_305),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_481),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_250),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_475),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_324),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_152),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_297),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_79),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_487),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_244),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_58),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_428),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_170),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_186),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_379),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_174),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_21),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_12),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_105),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_119),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_16),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_496),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_135),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_368),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_331),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_483),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_413),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_462),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_59),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_489),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_157),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_455),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_360),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_8),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_338),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_73),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_437),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_198),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_123),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_166),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_207),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_144),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_23),
.Y(n_585)
);

CKINVDCx16_ASAP7_75t_R g586 ( 
.A(n_451),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_169),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_72),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_124),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_341),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_256),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_279),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_35),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_36),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_76),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_449),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_93),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_191),
.Y(n_598)
);

BUFx5_ASAP7_75t_L g599 ( 
.A(n_384),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_494),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_445),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_359),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_427),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_443),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_486),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_439),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_132),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_478),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_35),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_401),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_235),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_442),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_46),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_433),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_392),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_336),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_499),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_261),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_363),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_498),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_412),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_447),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_304),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_414),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_419),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_426),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_181),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_4),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_69),
.Y(n_629)
);

BUFx2_ASAP7_75t_SL g630 ( 
.A(n_67),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_237),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_94),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_343),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_295),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_507),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_51),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_388),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_292),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_163),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_10),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_104),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_66),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_307),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_434),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_477),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_266),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_243),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_228),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_177),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_480),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_385),
.Y(n_651)
);

CKINVDCx16_ASAP7_75t_R g652 ( 
.A(n_458),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_67),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_420),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_362),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_43),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_249),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_502),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_202),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_11),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_46),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_484),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_161),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_441),
.Y(n_664)
);

CKINVDCx16_ASAP7_75t_R g665 ( 
.A(n_196),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_171),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_476),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_470),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_482),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_24),
.Y(n_670)
);

BUFx2_ASAP7_75t_SL g671 ( 
.A(n_464),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_306),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_66),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_260),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_485),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_403),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_469),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_345),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_215),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_128),
.Y(n_680)
);

CKINVDCx16_ASAP7_75t_R g681 ( 
.A(n_289),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_245),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_225),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_264),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_380),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_168),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_118),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_223),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_488),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_490),
.Y(n_690)
);

CKINVDCx16_ASAP7_75t_R g691 ( 
.A(n_479),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_106),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_205),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_328),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_472),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_31),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_161),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_364),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_316),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_98),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_18),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_222),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_491),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_167),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_229),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_88),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_238),
.Y(n_707)
);

BUFx5_ASAP7_75t_L g708 ( 
.A(n_501),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_474),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_457),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_79),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_399),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_216),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_503),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_202),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_98),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_89),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_339),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_196),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_492),
.Y(n_720)
);

INVx4_ASAP7_75t_R g721 ( 
.A(n_322),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_296),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_77),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_192),
.Y(n_724)
);

BUFx10_ASAP7_75t_L g725 ( 
.A(n_44),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_20),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_506),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_406),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_141),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_102),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_189),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_493),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_247),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_367),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_182),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_227),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_436),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_43),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_153),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_44),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_101),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_176),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_407),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_54),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_473),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_174),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_38),
.Y(n_747)
);

CKINVDCx14_ASAP7_75t_R g748 ( 
.A(n_27),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_31),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_80),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_117),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_375),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_299),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_335),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_185),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_28),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_208),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_282),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_146),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_241),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_330),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_12),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_134),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_533),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_665),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_533),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_608),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_535),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_535),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_707),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_565),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_526),
.B(n_0),
.Y(n_772)
);

INVxp67_ASAP7_75t_SL g773 ( 
.A(n_565),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_585),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_585),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_515),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_706),
.Y(n_777)
);

INVxp33_ASAP7_75t_SL g778 ( 
.A(n_571),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_603),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_515),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_722),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_706),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_723),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_744),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_748),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_511),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_723),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_512),
.Y(n_788)
);

INVxp67_ASAP7_75t_SL g789 ( 
.A(n_741),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_741),
.Y(n_790)
);

INVxp33_ASAP7_75t_SL g791 ( 
.A(n_696),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_513),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_731),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_748),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_716),
.Y(n_795)
);

CKINVDCx16_ASAP7_75t_R g796 ( 
.A(n_527),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_524),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_521),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_528),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_731),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_529),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_541),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_553),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_513),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_560),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_561),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_562),
.Y(n_807)
);

CKINVDCx16_ASAP7_75t_R g808 ( 
.A(n_586),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_581),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_582),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_687),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_731),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_588),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_607),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_609),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_613),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_632),
.Y(n_817)
);

INVxp33_ASAP7_75t_L g818 ( 
.A(n_700),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_531),
.Y(n_819)
);

INVxp33_ASAP7_75t_SL g820 ( 
.A(n_709),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_636),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_642),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_656),
.Y(n_823)
);

CKINVDCx16_ASAP7_75t_R g824 ( 
.A(n_652),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_663),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_731),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_670),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_532),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_679),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_713),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_681),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_691),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_629),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_630),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_719),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_536),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_603),
.Y(n_837)
);

INVxp67_ASAP7_75t_SL g838 ( 
.A(n_700),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_726),
.Y(n_839)
);

INVxp33_ASAP7_75t_SL g840 ( 
.A(n_760),
.Y(n_840)
);

INVxp33_ASAP7_75t_L g841 ( 
.A(n_740),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_548),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_740),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_534),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_550),
.Y(n_845)
);

INVxp67_ASAP7_75t_SL g846 ( 
.A(n_750),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_687),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_750),
.Y(n_848)
);

INVxp33_ASAP7_75t_SL g849 ( 
.A(n_555),
.Y(n_849)
);

CKINVDCx16_ASAP7_75t_R g850 ( 
.A(n_629),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_558),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_779),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_767),
.Y(n_853)
);

CKINVDCx16_ASAP7_75t_R g854 ( 
.A(n_796),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_779),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_779),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_779),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_793),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_800),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_797),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_837),
.Y(n_861)
);

OAI21x1_ASAP7_75t_L g862 ( 
.A1(n_812),
.A2(n_545),
.B(n_538),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_837),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_785),
.B(n_554),
.Y(n_864)
);

OAI22x1_ASAP7_75t_SL g865 ( 
.A1(n_792),
.A2(n_746),
.B1(n_578),
.B2(n_701),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_837),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_801),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_773),
.B(n_596),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_784),
.Y(n_869)
);

INVx4_ASAP7_75t_L g870 ( 
.A(n_837),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_812),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_802),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_826),
.A2(n_552),
.B(n_549),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_777),
.B(n_564),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_826),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_844),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_795),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_803),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_782),
.B(n_572),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_789),
.B(n_715),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_844),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_805),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_806),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_818),
.B(n_629),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_807),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_809),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_764),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_838),
.B(n_755),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_765),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_820),
.A2(n_746),
.B1(n_597),
.B2(n_556),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_810),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_813),
.Y(n_892)
);

AND2x6_ASAP7_75t_L g893 ( 
.A(n_772),
.B(n_534),
.Y(n_893)
);

OAI22x1_ASAP7_75t_R g894 ( 
.A1(n_792),
.A2(n_756),
.B1(n_757),
.B2(n_751),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_786),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_814),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_815),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_816),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_776),
.B(n_600),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_776),
.B(n_544),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_817),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_821),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_822),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_823),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_825),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_827),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_843),
.B(n_647),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_766),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_829),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_820),
.A2(n_517),
.B1(n_621),
.B2(n_620),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_818),
.B(n_841),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_780),
.B(n_794),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_830),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_835),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_911),
.B(n_850),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_886),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_853),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_854),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_853),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_895),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_895),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_889),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_889),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_910),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_865),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_890),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_886),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_908),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_884),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_898),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_898),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_901),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_901),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_876),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_876),
.Y(n_935)
);

CKINVDCx6p67_ASAP7_75t_R g936 ( 
.A(n_869),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_876),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_R g938 ( 
.A(n_912),
.B(n_770),
.Y(n_938)
);

NOR2xp67_ASAP7_75t_L g939 ( 
.A(n_877),
.B(n_831),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_869),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_905),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_905),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_876),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_908),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_894),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_899),
.B(n_808),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_877),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_882),
.B(n_824),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_881),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_880),
.B(n_781),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_882),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_914),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_881),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_900),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_882),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_892),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_892),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_892),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_907),
.B(n_833),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_900),
.B(n_780),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_892),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_881),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_902),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_902),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_R g965 ( 
.A(n_887),
.B(n_831),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_902),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_907),
.B(n_833),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_902),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_904),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_R g970 ( 
.A(n_887),
.B(n_832),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_881),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_852),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_914),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_852),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_864),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_904),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_904),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_904),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_914),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_914),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_864),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_858),
.B(n_794),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_906),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_906),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_R g985 ( 
.A(n_859),
.B(n_832),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_906),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_906),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_909),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_863),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_909),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_909),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_909),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_874),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_864),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_879),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_860),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_880),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_994),
.B(n_868),
.Y(n_998)
);

OAI22xp33_ASAP7_75t_L g999 ( 
.A1(n_947),
.A2(n_840),
.B1(n_517),
.B2(n_621),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_916),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_972),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_927),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_993),
.B(n_849),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_930),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_931),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_995),
.B(n_849),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_943),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_922),
.Y(n_1008)
);

AND2x6_ASAP7_75t_L g1009 ( 
.A(n_959),
.B(n_868),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_959),
.B(n_868),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_959),
.B(n_893),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_972),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_929),
.A2(n_893),
.B1(n_967),
.B2(n_960),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_974),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_936),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_997),
.B(n_840),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_974),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_967),
.B(n_893),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_967),
.B(n_893),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_915),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_918),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_943),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_989),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_943),
.Y(n_1024)
);

INVx4_ASAP7_75t_SL g1025 ( 
.A(n_996),
.Y(n_1025)
);

OR2x6_ASAP7_75t_L g1026 ( 
.A(n_975),
.B(n_880),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_950),
.B(n_788),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_952),
.B(n_893),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_981),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_928),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_989),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_956),
.B(n_907),
.Y(n_1032)
);

AND2x6_ASAP7_75t_L g1033 ( 
.A(n_932),
.B(n_888),
.Y(n_1033)
);

AND2x6_ASAP7_75t_L g1034 ( 
.A(n_933),
.B(n_888),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_946),
.B(n_948),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_939),
.B(n_867),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_941),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_942),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_934),
.Y(n_1039)
);

OAI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_926),
.A2(n_643),
.B1(n_646),
.B2(n_620),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_944),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_940),
.B(n_828),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_946),
.B(n_798),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_938),
.B(n_799),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_918),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_948),
.B(n_819),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_934),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_L g1048 ( 
.A(n_917),
.B(n_842),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_943),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_935),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_951),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_965),
.B(n_970),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_920),
.B(n_845),
.Y(n_1053)
);

INVxp67_ASAP7_75t_SL g1054 ( 
.A(n_935),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_919),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_937),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_955),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_923),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_957),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_937),
.Y(n_1060)
);

INVx8_ASAP7_75t_L g1061 ( 
.A(n_921),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_949),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_949),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_961),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_953),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_953),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_985),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_924),
.Y(n_1068)
);

BUFx10_ASAP7_75t_L g1069 ( 
.A(n_982),
.Y(n_1069)
);

AO22x2_ASAP7_75t_L g1070 ( 
.A1(n_924),
.A2(n_811),
.B1(n_847),
.B2(n_804),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_968),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_954),
.B(n_836),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_969),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_954),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_958),
.B(n_888),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_963),
.B(n_964),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_966),
.B(n_872),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_945),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_962),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_962),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_978),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_983),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_973),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_976),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_977),
.B(n_979),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_980),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_984),
.B(n_778),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_992),
.A2(n_791),
.B1(n_778),
.B2(n_646),
.Y(n_1088)
);

INVx4_ASAP7_75t_L g1089 ( 
.A(n_986),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_971),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_987),
.B(n_878),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_988),
.B(n_851),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_990),
.Y(n_1093)
);

INVx5_ASAP7_75t_L g1094 ( 
.A(n_971),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_991),
.A2(n_650),
.B1(n_728),
.B2(n_643),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_945),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_SL g1097 ( 
.A(n_925),
.B(n_650),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_952),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_947),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_993),
.B(n_791),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_916),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_996),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_996),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_996),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_918),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_972),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_952),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_918),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_993),
.B(n_883),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_972),
.Y(n_1110)
);

AND2x2_ASAP7_75t_SL g1111 ( 
.A(n_922),
.B(n_654),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_916),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_943),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_922),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_916),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_972),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_996),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_996),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_943),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_943),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_993),
.B(n_834),
.Y(n_1121)
);

INVx4_ASAP7_75t_L g1122 ( 
.A(n_952),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_972),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_918),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_L g1125 ( 
.A(n_947),
.B(n_896),
.C(n_891),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_993),
.B(n_885),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_916),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_959),
.B(n_654),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1102),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1121),
.B(n_913),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_1008),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1001),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1009),
.B(n_897),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1012),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1009),
.B(n_903),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1009),
.B(n_841),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1089),
.B(n_728),
.Y(n_1137)
);

NOR2xp67_ASAP7_75t_L g1138 ( 
.A(n_1053),
.B(n_768),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1009),
.B(n_846),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1000),
.B(n_848),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1100),
.B(n_804),
.Y(n_1141)
);

OAI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1095),
.A2(n_847),
.B1(n_811),
.B2(n_519),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1003),
.B(n_1006),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_1114),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1109),
.B(n_627),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1014),
.Y(n_1146)
);

NAND2x1_ASAP7_75t_L g1147 ( 
.A(n_1024),
.B(n_870),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_1099),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1126),
.B(n_683),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1103),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1017),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1104),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_998),
.Y(n_1153)
);

NOR3xp33_ASAP7_75t_L g1154 ( 
.A(n_1016),
.B(n_749),
.C(n_747),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1076),
.B(n_762),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1087),
.B(n_559),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1067),
.B(n_563),
.Y(n_1157)
);

INVxp67_ASAP7_75t_L g1158 ( 
.A(n_1058),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_1042),
.B(n_769),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1111),
.A2(n_530),
.B1(n_557),
.B2(n_725),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1089),
.B(n_573),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1023),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1040),
.B(n_576),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1027),
.B(n_580),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1010),
.B(n_763),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1013),
.A2(n_584),
.B1(n_587),
.B2(n_583),
.Y(n_1166)
);

NOR3xp33_ASAP7_75t_L g1167 ( 
.A(n_999),
.B(n_593),
.C(n_589),
.Y(n_1167)
);

AO221x1_ASAP7_75t_L g1168 ( 
.A1(n_1070),
.A2(n_743),
.B1(n_705),
.B2(n_603),
.C(n_611),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1117),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1033),
.B(n_594),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1031),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1020),
.B(n_787),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1061),
.B(n_771),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1118),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1061),
.B(n_774),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1098),
.B(n_1107),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1106),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1035),
.A2(n_612),
.B1(n_626),
.B2(n_610),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_1043),
.B(n_839),
.C(n_598),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1000),
.Y(n_1180)
);

OAI22x1_ASAP7_75t_R g1181 ( 
.A1(n_1105),
.A2(n_628),
.B1(n_639),
.B2(n_595),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1098),
.B(n_1107),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1055),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1002),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1033),
.B(n_640),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1002),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1033),
.B(n_641),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1025),
.B(n_775),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1075),
.B(n_649),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1072),
.B(n_1021),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1045),
.B(n_783),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1110),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1092),
.B(n_790),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1116),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_1026),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1033),
.B(n_653),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1122),
.B(n_659),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1004),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1007),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1046),
.A2(n_637),
.B1(n_644),
.B2(n_634),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1025),
.B(n_1075),
.Y(n_1201)
);

AND2x6_ASAP7_75t_L g1202 ( 
.A(n_1011),
.B(n_544),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1004),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1034),
.B(n_660),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1034),
.B(n_661),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_SL g1206 ( 
.A(n_1122),
.B(n_530),
.Y(n_1206)
);

INVx4_ASAP7_75t_L g1207 ( 
.A(n_1034),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1030),
.B(n_666),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1034),
.B(n_673),
.Y(n_1209)
);

NOR2xp67_ASAP7_75t_L g1210 ( 
.A(n_1041),
.B(n_648),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1007),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1007),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1108),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1018),
.A2(n_873),
.B(n_862),
.C(n_682),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1032),
.B(n_680),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1005),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1085),
.B(n_686),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1077),
.B(n_688),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1069),
.B(n_692),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1091),
.B(n_693),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1083),
.B(n_697),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1026),
.B(n_725),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1022),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1022),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1029),
.B(n_725),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1128),
.A2(n_530),
.B1(n_557),
.B2(n_647),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1084),
.B(n_702),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1069),
.B(n_704),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1093),
.B(n_711),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1052),
.B(n_717),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1086),
.B(n_724),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1123),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1005),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1101),
.B(n_729),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1101),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1112),
.B(n_730),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1019),
.A2(n_675),
.B1(n_698),
.B2(n_694),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1015),
.B(n_735),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1112),
.B(n_738),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1048),
.B(n_739),
.Y(n_1240)
);

NOR3xp33_ASAP7_75t_L g1241 ( 
.A(n_1125),
.B(n_759),
.C(n_742),
.Y(n_1241)
);

INVx4_ASAP7_75t_L g1242 ( 
.A(n_1022),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1036),
.A2(n_718),
.B1(n_733),
.B2(n_699),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1115),
.B(n_546),
.Y(n_1244)
);

NOR2x1p5_ASAP7_75t_L g1245 ( 
.A(n_1124),
.B(n_754),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1115),
.B(n_567),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1127),
.B(n_567),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1088),
.B(n_616),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1044),
.B(n_631),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1127),
.B(n_871),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1037),
.B(n_871),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1074),
.B(n_557),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1028),
.B(n_510),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1068),
.B(n_871),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1038),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1049),
.B(n_1113),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1051),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1096),
.B(n_514),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1057),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1049),
.B(n_518),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1057),
.B(n_871),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1050),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1059),
.A2(n_568),
.B1(n_604),
.B2(n_590),
.Y(n_1263)
);

OAI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1097),
.A2(n_622),
.B1(n_624),
.B2(n_516),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1064),
.B(n_520),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1078),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1071),
.B(n_875),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1113),
.B(n_522),
.Y(n_1268)
);

INVx4_ASAP7_75t_L g1269 ( 
.A(n_1113),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1073),
.B(n_523),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1081),
.B(n_875),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1082),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1050),
.B(n_525),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1119),
.B(n_537),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1070),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1039),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1063),
.B(n_875),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1047),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1056),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1065),
.A2(n_671),
.B1(n_590),
.B2(n_604),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1063),
.B(n_875),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1079),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1090),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1080),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1090),
.B(n_539),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1119),
.B(n_540),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1054),
.B(n_542),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1060),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1024),
.A2(n_614),
.B(n_568),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1094),
.B(n_1120),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1060),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1120),
.B(n_543),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1060),
.B(n_547),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1062),
.A2(n_669),
.B1(n_695),
.B2(n_614),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1062),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1062),
.B(n_551),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1119),
.A2(n_695),
.B1(n_669),
.B2(n_569),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1094),
.A2(n_570),
.B1(n_574),
.B2(n_566),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1066),
.B(n_575),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1066),
.A2(n_579),
.B1(n_591),
.B2(n_577),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1066),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1094),
.B(n_863),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1089),
.B(n_592),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_998),
.B(n_0),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_998),
.B(n_1),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1121),
.B(n_601),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1055),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1089),
.B(n_602),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1102),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1009),
.A2(n_606),
.B1(n_615),
.B2(n_605),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1009),
.B(n_599),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_998),
.B(n_1),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1121),
.B(n_617),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1121),
.B(n_618),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1183),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1143),
.B(n_2),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1164),
.A2(n_1184),
.B(n_1180),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1141),
.B(n_619),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1156),
.B(n_623),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1130),
.B(n_2),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1193),
.B(n_3),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1253),
.A2(n_633),
.B(n_625),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1153),
.B(n_3),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1289),
.A2(n_1198),
.B(n_1186),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1145),
.B(n_4),
.Y(n_1325)
);

AO21x1_ASAP7_75t_L g1326 ( 
.A1(n_1289),
.A2(n_866),
.B(n_708),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1158),
.B(n_635),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1206),
.B(n_638),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1149),
.B(n_5),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1206),
.B(n_645),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1131),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1203),
.A2(n_655),
.B(n_651),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1172),
.B(n_5),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1179),
.A2(n_658),
.B(n_662),
.C(n_657),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1306),
.B(n_6),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1190),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1216),
.A2(n_667),
.B(n_664),
.Y(n_1337)
);

O2A1O1Ixp5_ASAP7_75t_L g1338 ( 
.A1(n_1260),
.A2(n_1268),
.B(n_1286),
.C(n_1274),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1313),
.B(n_1314),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1307),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1233),
.A2(n_668),
.B1(n_674),
.B2(n_672),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1257),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1154),
.A2(n_9),
.B(n_6),
.C(n_7),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1163),
.B(n_7),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1235),
.A2(n_677),
.B(n_676),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1207),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1250),
.A2(n_684),
.B(n_678),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1304),
.B(n_9),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1305),
.B(n_1312),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1259),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1248),
.A2(n_603),
.B1(n_689),
.B2(n_685),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1155),
.B(n_10),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1138),
.B(n_690),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1179),
.A2(n_710),
.B(n_703),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1144),
.B(n_712),
.Y(n_1355)
);

INVx5_ASAP7_75t_L g1356 ( 
.A(n_1207),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1242),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1261),
.A2(n_720),
.B(n_714),
.Y(n_1358)
);

AOI21xp33_ASAP7_75t_L g1359 ( 
.A1(n_1240),
.A2(n_1142),
.B(n_1200),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1292),
.A2(n_732),
.B(n_727),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1287),
.A2(n_736),
.B(n_734),
.Y(n_1361)
);

OR2x6_ASAP7_75t_L g1362 ( 
.A(n_1201),
.B(n_721),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1148),
.B(n_737),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1140),
.B(n_11),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1277),
.A2(n_752),
.B(n_745),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1281),
.A2(n_758),
.B(n_753),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1201),
.B(n_761),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1218),
.A2(n_856),
.B(n_855),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1140),
.B(n_13),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1137),
.B(n_13),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1246),
.A2(n_856),
.B(n_855),
.Y(n_1371)
);

AO21x1_ASAP7_75t_L g1372 ( 
.A1(n_1246),
.A2(n_708),
.B(n_599),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1159),
.B(n_14),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1242),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1220),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_1375)
);

CKINVDCx10_ASAP7_75t_R g1376 ( 
.A(n_1181),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_R g1377 ( 
.A(n_1266),
.B(n_230),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1132),
.Y(n_1378)
);

O2A1O1Ixp5_ASAP7_75t_L g1379 ( 
.A1(n_1265),
.A2(n_18),
.B(n_15),
.C(n_17),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1195),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1129),
.B(n_17),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1225),
.B(n_19),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1150),
.B(n_19),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1152),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1169),
.B(n_20),
.Y(n_1385)
);

A2O1A1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1178),
.A2(n_856),
.B(n_857),
.C(n_855),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1174),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1256),
.A2(n_856),
.B(n_855),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1309),
.B(n_1136),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1214),
.A2(n_708),
.B(n_599),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1136),
.B(n_22),
.Y(n_1391)
);

BUFx4f_ASAP7_75t_L g1392 ( 
.A(n_1173),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1249),
.A2(n_861),
.B(n_857),
.C(n_708),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1222),
.B(n_25),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1134),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1255),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1247),
.A2(n_861),
.B(n_857),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1262),
.A2(n_708),
.B(n_599),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1167),
.B(n_857),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1247),
.A2(n_861),
.B(n_232),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1269),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1273),
.A2(n_861),
.B(n_233),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1139),
.B(n_25),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1210),
.B(n_708),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1217),
.A2(n_234),
.B(n_231),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1175),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1212),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_SL g1408 ( 
.A(n_1213),
.B(n_599),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1272),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1215),
.A2(n_239),
.B(n_236),
.Y(n_1410)
);

OAI21xp33_ASAP7_75t_L g1411 ( 
.A1(n_1219),
.A2(n_26),
.B(n_27),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1270),
.A2(n_246),
.B(n_240),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1271),
.A2(n_1251),
.B(n_1285),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1191),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1188),
.B(n_26),
.Y(n_1415)
);

INVxp33_ASAP7_75t_L g1416 ( 
.A(n_1189),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1147),
.A2(n_251),
.B(n_248),
.Y(n_1417)
);

OR2x6_ASAP7_75t_SL g1418 ( 
.A(n_1297),
.B(n_1166),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1234),
.A2(n_253),
.B(n_252),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1283),
.A2(n_708),
.B(n_599),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1212),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1139),
.B(n_28),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_1254),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1146),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1165),
.B(n_29),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1188),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1160),
.A2(n_32),
.B1(n_29),
.B2(n_30),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1151),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1236),
.A2(n_255),
.B(n_254),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_1245),
.Y(n_1430)
);

OAI21xp33_ASAP7_75t_L g1431 ( 
.A1(n_1228),
.A2(n_30),
.B(n_32),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1276),
.Y(n_1432)
);

OAI21xp33_ASAP7_75t_L g1433 ( 
.A1(n_1239),
.A2(n_33),
.B(n_34),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1157),
.B(n_33),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1298),
.B(n_1230),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1133),
.A2(n_258),
.B(n_257),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1269),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1135),
.A2(n_263),
.B(n_262),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1238),
.B(n_34),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1244),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1311),
.A2(n_37),
.B(n_39),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1311),
.A2(n_39),
.B(n_40),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1212),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1162),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1258),
.B(n_40),
.Y(n_1445)
);

CKINVDCx10_ASAP7_75t_R g1446 ( 
.A(n_1168),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1171),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1252),
.B(n_41),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1176),
.B(n_41),
.Y(n_1449)
);

NOR2xp67_ASAP7_75t_L g1450 ( 
.A(n_1296),
.B(n_267),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1223),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1298),
.B(n_42),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1177),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1182),
.B(n_42),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1243),
.B(n_45),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1221),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1223),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1275),
.B(n_45),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1223),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1192),
.Y(n_1460)
);

AND2x6_ASAP7_75t_L g1461 ( 
.A(n_1224),
.B(n_268),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1194),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1241),
.B(n_1310),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1293),
.A2(n_270),
.B(n_269),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1299),
.A2(n_272),
.B(n_271),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1290),
.A2(n_274),
.B(n_273),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1227),
.B(n_47),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1303),
.A2(n_276),
.B(n_275),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1224),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1308),
.A2(n_278),
.B(n_277),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_R g1471 ( 
.A(n_1224),
.B(n_280),
.Y(n_1471)
);

AOI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1288),
.A2(n_284),
.B(n_281),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1170),
.A2(n_286),
.B(n_285),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1231),
.B(n_48),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1229),
.B(n_49),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_1199),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1185),
.A2(n_288),
.B(n_287),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1208),
.B(n_49),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1226),
.B(n_50),
.Y(n_1479)
);

O2A1O1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1161),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1187),
.B(n_53),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1199),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1196),
.A2(n_291),
.B(n_290),
.Y(n_1483)
);

AO21x1_ASAP7_75t_L g1484 ( 
.A1(n_1263),
.A2(n_294),
.B(n_293),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1297),
.B(n_54),
.Y(n_1485)
);

AND2x4_ASAP7_75t_SL g1486 ( 
.A(n_1211),
.B(n_55),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1204),
.B(n_1205),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1237),
.A2(n_55),
.B(n_56),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1209),
.B(n_56),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1264),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1490)
);

BUFx4f_ASAP7_75t_L g1491 ( 
.A(n_1211),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1302),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1197),
.B(n_57),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1263),
.B(n_60),
.Y(n_1494)
);

A2O1A1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1278),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1279),
.A2(n_61),
.B(n_62),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1291),
.B(n_1295),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1339),
.A2(n_1301),
.B(n_1267),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1324),
.A2(n_1302),
.B(n_1284),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1359),
.A2(n_1232),
.B1(n_1282),
.B2(n_1280),
.Y(n_1500)
);

BUFx4f_ASAP7_75t_L g1501 ( 
.A(n_1492),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1392),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1414),
.Y(n_1503)
);

NOR2x1_ASAP7_75t_SL g1504 ( 
.A(n_1356),
.B(n_1202),
.Y(n_1504)
);

AOI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1371),
.A2(n_1202),
.B(n_1294),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1416),
.B(n_1300),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1317),
.A2(n_1202),
.B(n_301),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1319),
.B(n_1318),
.Y(n_1508)
);

O2A1O1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1316),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1344),
.A2(n_68),
.B1(n_63),
.B2(n_64),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1336),
.B(n_68),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1406),
.B(n_1456),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1434),
.B(n_69),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1492),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1315),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1373),
.B(n_70),
.Y(n_1516)
);

INVx4_ASAP7_75t_L g1517 ( 
.A(n_1356),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1384),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1413),
.A2(n_302),
.B(n_300),
.Y(n_1519)
);

BUFx2_ASAP7_75t_SL g1520 ( 
.A(n_1340),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1435),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1474),
.A2(n_74),
.B(n_71),
.C(n_73),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1320),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1396),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1370),
.A2(n_80),
.B1(n_75),
.B2(n_78),
.C(n_81),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1432),
.B(n_78),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1346),
.B(n_81),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1346),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1423),
.B(n_82),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1349),
.B(n_82),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1333),
.B(n_83),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1321),
.B(n_83),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1352),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1331),
.B(n_1418),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1445),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1449),
.B(n_87),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1368),
.A2(n_308),
.B(n_303),
.Y(n_1537)
);

NOR2x1_ASAP7_75t_L g1538 ( 
.A(n_1443),
.B(n_309),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1402),
.A2(n_312),
.B(n_311),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1342),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1350),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1380),
.B(n_87),
.Y(n_1542)
);

O2A1O1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1448),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1327),
.B(n_90),
.Y(n_1544)
);

A2O1A1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1335),
.A2(n_1431),
.B(n_1411),
.C(n_1488),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1492),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1409),
.B(n_91),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1449),
.B(n_92),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1426),
.B(n_93),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1389),
.B(n_95),
.Y(n_1550)
);

O2A1O1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1452),
.A2(n_97),
.B(n_95),
.C(n_96),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1430),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1325),
.B(n_96),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1454),
.B(n_97),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1400),
.A2(n_314),
.B(n_313),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1415),
.B(n_99),
.Y(n_1556)
);

A2O1A1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1467),
.A2(n_1425),
.B(n_1433),
.C(n_1329),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1454),
.B(n_99),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1491),
.B(n_100),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1364),
.B(n_100),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1397),
.A2(n_318),
.B(n_317),
.Y(n_1561)
);

O2A1O1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1343),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_1562)
);

O2A1O1Ixp5_ASAP7_75t_L g1563 ( 
.A1(n_1328),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1443),
.B(n_509),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1415),
.B(n_106),
.Y(n_1565)
);

OAI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1337),
.A2(n_107),
.B(n_108),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1348),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1491),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1369),
.B(n_110),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1427),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_1570)
);

A2O1A1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1475),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1412),
.A2(n_320),
.B(n_319),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1476),
.B(n_114),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1378),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1395),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1424),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1439),
.B(n_115),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1407),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1382),
.B(n_115),
.Y(n_1579)
);

INVx5_ASAP7_75t_L g1580 ( 
.A(n_1461),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1485),
.B(n_116),
.Y(n_1581)
);

INVxp33_ASAP7_75t_L g1582 ( 
.A(n_1394),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1460),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1428),
.Y(n_1584)
);

OR2x6_ASAP7_75t_L g1585 ( 
.A(n_1362),
.B(n_116),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1476),
.B(n_117),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_SL g1587 ( 
.A1(n_1441),
.A2(n_118),
.B(n_119),
.Y(n_1587)
);

O2A1O1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1478),
.A2(n_122),
.B(n_120),
.C(n_121),
.Y(n_1588)
);

OA22x2_ASAP7_75t_L g1589 ( 
.A1(n_1362),
.A2(n_123),
.B1(n_120),
.B2(n_121),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1330),
.B(n_124),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1444),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1351),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1487),
.A2(n_323),
.B(n_321),
.Y(n_1593)
);

CKINVDCx16_ASAP7_75t_R g1594 ( 
.A(n_1377),
.Y(n_1594)
);

OAI21xp33_ASAP7_75t_L g1595 ( 
.A1(n_1496),
.A2(n_125),
.B(n_126),
.Y(n_1595)
);

OAI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1391),
.A2(n_127),
.B(n_128),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1447),
.Y(n_1597)
);

INVx3_ASAP7_75t_SL g1598 ( 
.A(n_1486),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1453),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1494),
.B(n_129),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_L g1601 ( 
.A1(n_1463),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_1601)
);

A2O1A1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1493),
.A2(n_133),
.B(n_130),
.C(n_131),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1458),
.B(n_1323),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1381),
.B(n_133),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1363),
.B(n_1376),
.Y(n_1605)
);

INVx4_ASAP7_75t_L g1606 ( 
.A(n_1407),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1357),
.B(n_325),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1476),
.B(n_134),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1490),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1357),
.B(n_1374),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1383),
.B(n_136),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1455),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1407),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1403),
.B(n_138),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1422),
.B(n_139),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1421),
.Y(n_1616)
);

BUFx12f_ASAP7_75t_L g1617 ( 
.A(n_1421),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1347),
.A2(n_140),
.B(n_141),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1462),
.B(n_140),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1385),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_SL g1621 ( 
.A(n_1408),
.B(n_326),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1446),
.B(n_142),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1405),
.A2(n_329),
.B(n_327),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1497),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1481),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1482),
.B(n_142),
.Y(n_1626)
);

O2A1O1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1440),
.A2(n_146),
.B(n_143),
.C(n_145),
.Y(n_1627)
);

NAND3xp33_ASAP7_75t_SL g1628 ( 
.A(n_1375),
.B(n_143),
.C(n_145),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1479),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_1629)
);

INVx4_ASAP7_75t_L g1630 ( 
.A(n_1421),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1387),
.B(n_147),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1482),
.B(n_148),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_SL g1633 ( 
.A1(n_1480),
.A2(n_152),
.B(n_150),
.C(n_151),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1367),
.B(n_150),
.Y(n_1634)
);

OA21x2_ASAP7_75t_L g1635 ( 
.A1(n_1390),
.A2(n_333),
.B(n_332),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1482),
.B(n_151),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1457),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1451),
.B(n_153),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1457),
.B(n_154),
.Y(n_1639)
);

O2A1O1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1495),
.A2(n_156),
.B(n_154),
.C(n_155),
.Y(n_1640)
);

O2A1O1Ixp33_ASAP7_75t_L g1641 ( 
.A1(n_1442),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1341),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1459),
.Y(n_1643)
);

NAND3xp33_ASAP7_75t_SL g1644 ( 
.A(n_1354),
.B(n_158),
.C(n_159),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_R g1645 ( 
.A(n_1457),
.B(n_334),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1489),
.Y(n_1646)
);

O2A1O1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1379),
.A2(n_163),
.B(n_160),
.C(n_162),
.Y(n_1647)
);

OAI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1355),
.A2(n_1353),
.B1(n_1399),
.B2(n_1450),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1518),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1508),
.A2(n_1334),
.B(n_1338),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1507),
.A2(n_1420),
.B(n_1398),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1581),
.B(n_1459),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1624),
.B(n_1469),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1503),
.B(n_1469),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1545),
.A2(n_1484),
.B(n_1410),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1524),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1505),
.A2(n_1372),
.B(n_1326),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1499),
.A2(n_1537),
.B(n_1519),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1561),
.A2(n_1472),
.B(n_1388),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1513),
.B(n_1374),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1568),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1557),
.A2(n_1393),
.B(n_1419),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1618),
.A2(n_1361),
.B(n_1360),
.Y(n_1663)
);

AO31x2_ASAP7_75t_L g1664 ( 
.A1(n_1498),
.A2(n_1386),
.A3(n_1477),
.B(n_1473),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_L g1665 ( 
.A1(n_1555),
.A2(n_1483),
.B(n_1465),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1572),
.A2(n_1429),
.B(n_1466),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1603),
.B(n_1401),
.Y(n_1667)
);

OAI21x1_ASAP7_75t_L g1668 ( 
.A1(n_1539),
.A2(n_1464),
.B(n_1417),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1568),
.Y(n_1669)
);

NAND2x1p5_ASAP7_75t_L g1670 ( 
.A(n_1580),
.B(n_1401),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1520),
.Y(n_1671)
);

OAI21x1_ASAP7_75t_L g1672 ( 
.A1(n_1623),
.A2(n_1438),
.B(n_1436),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1576),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1583),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1544),
.A2(n_1332),
.B1(n_1345),
.B2(n_1437),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_R g1676 ( 
.A(n_1594),
.B(n_1437),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1577),
.A2(n_1468),
.B1(n_1470),
.B2(n_1404),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1635),
.A2(n_1358),
.B(n_1365),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1595),
.A2(n_1322),
.B(n_1366),
.C(n_1461),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1506),
.A2(n_1461),
.B1(n_1471),
.B2(n_165),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1635),
.A2(n_1461),
.B(n_162),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1566),
.A2(n_164),
.B(n_165),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1512),
.B(n_164),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1552),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1641),
.A2(n_166),
.B(n_167),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1584),
.Y(n_1686)
);

OAI21xp33_ASAP7_75t_L g1687 ( 
.A1(n_1596),
.A2(n_168),
.B(n_169),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1620),
.B(n_1550),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1617),
.Y(n_1689)
);

AOI211x1_ASAP7_75t_L g1690 ( 
.A1(n_1600),
.A2(n_1548),
.B(n_1554),
.C(n_1536),
.Y(n_1690)
);

OAI22x1_ASAP7_75t_L g1691 ( 
.A1(n_1534),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1593),
.A2(n_342),
.B(n_340),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1648),
.A2(n_172),
.B(n_173),
.Y(n_1693)
);

OAI21x1_ASAP7_75t_L g1694 ( 
.A1(n_1538),
.A2(n_346),
.B(n_344),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1580),
.A2(n_173),
.B(n_175),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1580),
.A2(n_175),
.B(n_176),
.Y(n_1696)
);

AOI211x1_ASAP7_75t_L g1697 ( 
.A1(n_1558),
.A2(n_1535),
.B(n_1567),
.C(n_1612),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1553),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_1698)
);

AO31x2_ASAP7_75t_L g1699 ( 
.A1(n_1625),
.A2(n_415),
.A3(n_505),
.B(n_504),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1644),
.A2(n_1522),
.B(n_1560),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1568),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1578),
.Y(n_1702)
);

NAND2x1p5_ASAP7_75t_L g1703 ( 
.A(n_1501),
.B(n_347),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1562),
.A2(n_178),
.B(n_179),
.Y(n_1704)
);

A2O1A1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1588),
.A2(n_180),
.B(n_182),
.C(n_183),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1556),
.B(n_180),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1646),
.B(n_184),
.Y(n_1707)
);

INVx4_ASAP7_75t_L g1708 ( 
.A(n_1598),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1530),
.B(n_184),
.Y(n_1709)
);

AOI21x1_ASAP7_75t_L g1710 ( 
.A1(n_1614),
.A2(n_349),
.B(n_348),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1569),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1501),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1621),
.A2(n_187),
.B(n_188),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1502),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1607),
.A2(n_189),
.B(n_190),
.Y(n_1715)
);

NAND2x1p5_ASAP7_75t_L g1716 ( 
.A(n_1517),
.B(n_350),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_SL g1717 ( 
.A1(n_1587),
.A2(n_190),
.B(n_191),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1597),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1607),
.A2(n_192),
.B(n_193),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1610),
.B(n_193),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1540),
.Y(n_1721)
);

OAI21x1_ASAP7_75t_L g1722 ( 
.A1(n_1528),
.A2(n_353),
.B(n_351),
.Y(n_1722)
);

OR2x6_ASAP7_75t_L g1723 ( 
.A(n_1585),
.B(n_354),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1615),
.A2(n_194),
.B(n_195),
.Y(n_1724)
);

A2O1A1Ixp33_ASAP7_75t_L g1725 ( 
.A1(n_1590),
.A2(n_194),
.B(n_195),
.C(n_197),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1541),
.Y(n_1726)
);

O2A1O1Ixp33_ASAP7_75t_SL g1727 ( 
.A1(n_1602),
.A2(n_197),
.B(n_198),
.C(n_199),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1631),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1514),
.B(n_200),
.Y(n_1729)
);

AO22x2_ASAP7_75t_L g1730 ( 
.A1(n_1628),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1613),
.Y(n_1731)
);

OAI21xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1642),
.A2(n_1525),
.B(n_1510),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1574),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1514),
.B(n_203),
.Y(n_1734)
);

OAI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1528),
.A2(n_356),
.B(n_355),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1604),
.B(n_1611),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1647),
.A2(n_358),
.B(n_357),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1575),
.Y(n_1738)
);

INVx4_ASAP7_75t_L g1739 ( 
.A(n_1613),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1571),
.A2(n_204),
.B(n_205),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1605),
.Y(n_1741)
);

NOR4xp25_ASAP7_75t_L g1742 ( 
.A(n_1543),
.B(n_206),
.C(n_207),
.D(n_208),
.Y(n_1742)
);

BUFx4_ASAP7_75t_SL g1743 ( 
.A(n_1585),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1514),
.B(n_206),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1515),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1565),
.B(n_209),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1589),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_1747)
);

BUFx4f_ASAP7_75t_SL g1748 ( 
.A(n_1613),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1582),
.B(n_210),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1532),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1504),
.A2(n_1610),
.B(n_1633),
.Y(n_1751)
);

XOR2xp5_ASAP7_75t_L g1752 ( 
.A(n_1546),
.B(n_361),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1616),
.Y(n_1753)
);

AO22x2_ASAP7_75t_L g1754 ( 
.A1(n_1591),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_1754)
);

O2A1O1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1627),
.A2(n_214),
.B(n_215),
.C(n_216),
.Y(n_1755)
);

O2A1O1Ixp33_ASAP7_75t_SL g1756 ( 
.A1(n_1559),
.A2(n_217),
.B(n_218),
.C(n_219),
.Y(n_1756)
);

INVxp67_ASAP7_75t_SL g1757 ( 
.A(n_1637),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1622),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1526),
.B(n_220),
.Y(n_1759)
);

OA21x2_ASAP7_75t_L g1760 ( 
.A1(n_1655),
.A2(n_1563),
.B(n_1547),
.Y(n_1760)
);

OA21x2_ASAP7_75t_L g1761 ( 
.A1(n_1657),
.A2(n_1586),
.B(n_1573),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1649),
.Y(n_1762)
);

NOR3xp33_ASAP7_75t_L g1763 ( 
.A(n_1732),
.B(n_1523),
.C(n_1533),
.Y(n_1763)
);

BUFx12f_ASAP7_75t_L g1764 ( 
.A(n_1741),
.Y(n_1764)
);

OAI222xp33_ASAP7_75t_L g1765 ( 
.A1(n_1747),
.A2(n_1680),
.B1(n_1728),
.B2(n_1758),
.C1(n_1723),
.C2(n_1736),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1656),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1687),
.A2(n_1609),
.B1(n_1570),
.B2(n_1592),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1697),
.A2(n_1629),
.B1(n_1521),
.B2(n_1531),
.Y(n_1768)
);

OR2x6_ASAP7_75t_L g1769 ( 
.A(n_1723),
.B(n_1564),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1712),
.B(n_1517),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1652),
.B(n_1638),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1682),
.A2(n_1601),
.B(n_1509),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_L g1773 ( 
.A(n_1725),
.B(n_1700),
.C(n_1650),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1688),
.B(n_1516),
.Y(n_1774)
);

OAI21x1_ASAP7_75t_SL g1775 ( 
.A1(n_1740),
.A2(n_1640),
.B(n_1551),
.Y(n_1775)
);

OA21x2_ASAP7_75t_L g1776 ( 
.A1(n_1681),
.A2(n_1636),
.B(n_1608),
.Y(n_1776)
);

AO21x2_ASAP7_75t_L g1777 ( 
.A1(n_1678),
.A2(n_1619),
.B(n_1645),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1685),
.A2(n_1599),
.B1(n_1500),
.B2(n_1634),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1673),
.Y(n_1779)
);

OAI21x1_ASAP7_75t_SL g1780 ( 
.A1(n_1755),
.A2(n_1632),
.B(n_1626),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1702),
.Y(n_1781)
);

OR2x6_ASAP7_75t_L g1782 ( 
.A(n_1693),
.B(n_1690),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1746),
.A2(n_1579),
.B1(n_1542),
.B2(n_1549),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1757),
.B(n_1606),
.Y(n_1784)
);

OAI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1658),
.A2(n_1643),
.B(n_1527),
.Y(n_1785)
);

INVxp67_ASAP7_75t_L g1786 ( 
.A(n_1654),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1674),
.Y(n_1787)
);

OA21x2_ASAP7_75t_L g1788 ( 
.A1(n_1662),
.A2(n_1639),
.B(n_1529),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1676),
.Y(n_1789)
);

OAI21x1_ASAP7_75t_SL g1790 ( 
.A1(n_1717),
.A2(n_1630),
.B(n_1606),
.Y(n_1790)
);

O2A1O1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1705),
.A2(n_1727),
.B(n_1759),
.C(n_1698),
.Y(n_1791)
);

OAI21x1_ASAP7_75t_L g1792 ( 
.A1(n_1659),
.A2(n_1511),
.B(n_1564),
.Y(n_1792)
);

NAND2xp33_ASAP7_75t_R g1793 ( 
.A(n_1689),
.B(n_220),
.Y(n_1793)
);

CKINVDCx20_ASAP7_75t_R g1794 ( 
.A(n_1684),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1686),
.Y(n_1795)
);

OAI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1742),
.A2(n_1704),
.B1(n_1709),
.B2(n_1724),
.C(n_1663),
.Y(n_1796)
);

INVx5_ASAP7_75t_L g1797 ( 
.A(n_1661),
.Y(n_1797)
);

BUFx2_ASAP7_75t_SL g1798 ( 
.A(n_1739),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1667),
.B(n_1616),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1754),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1718),
.Y(n_1801)
);

OAI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1713),
.A2(n_221),
.B(n_224),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1653),
.B(n_224),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1666),
.A2(n_225),
.B(n_226),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1721),
.Y(n_1805)
);

AO31x2_ASAP7_75t_L g1806 ( 
.A1(n_1651),
.A2(n_1677),
.A3(n_1679),
.B(n_1733),
.Y(n_1806)
);

BUFx6f_ASAP7_75t_L g1807 ( 
.A(n_1712),
.Y(n_1807)
);

OAI21x1_ASAP7_75t_L g1808 ( 
.A1(n_1668),
.A2(n_468),
.B(n_365),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1660),
.B(n_226),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_SL g1810 ( 
.A1(n_1754),
.A2(n_366),
.B1(n_369),
.B2(n_370),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1731),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1671),
.B(n_1729),
.Y(n_1812)
);

NAND2x1p5_ASAP7_75t_L g1813 ( 
.A(n_1712),
.B(n_371),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_SL g1814 ( 
.A1(n_1730),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_SL g1815 ( 
.A1(n_1743),
.A2(n_376),
.B1(n_377),
.B2(n_378),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1726),
.Y(n_1816)
);

OAI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1715),
.A2(n_381),
.B(n_382),
.Y(n_1817)
);

OAI21x1_ASAP7_75t_L g1818 ( 
.A1(n_1665),
.A2(n_383),
.B(n_386),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1672),
.A2(n_389),
.B(n_390),
.Y(n_1819)
);

OAI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1719),
.A2(n_1751),
.B(n_1696),
.Y(n_1820)
);

NAND2x1p5_ASAP7_75t_L g1821 ( 
.A(n_1661),
.B(n_391),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1707),
.B(n_393),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1738),
.Y(n_1823)
);

OAI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1695),
.A2(n_394),
.B(n_395),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1699),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1773),
.A2(n_1730),
.B1(n_1711),
.B2(n_1750),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1769),
.A2(n_1675),
.B(n_1737),
.Y(n_1827)
);

OAI21x1_ASAP7_75t_L g1828 ( 
.A1(n_1785),
.A2(n_1710),
.B(n_1694),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1762),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1781),
.B(n_1749),
.Y(n_1830)
);

OA21x2_ASAP7_75t_L g1831 ( 
.A1(n_1825),
.A2(n_1792),
.B(n_1820),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1762),
.B(n_1706),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1769),
.A2(n_1692),
.B(n_1670),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1763),
.A2(n_1691),
.B1(n_1752),
.B2(n_1734),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1779),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1779),
.B(n_1729),
.Y(n_1836)
);

OA21x2_ASAP7_75t_L g1837 ( 
.A1(n_1804),
.A2(n_1808),
.B(n_1818),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1795),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1823),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1806),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1786),
.Y(n_1841)
);

AO21x2_ASAP7_75t_L g1842 ( 
.A1(n_1777),
.A2(n_1722),
.B(n_1735),
.Y(n_1842)
);

OA21x2_ASAP7_75t_L g1843 ( 
.A1(n_1819),
.A2(n_1720),
.B(n_1683),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1796),
.A2(n_1756),
.B(n_1716),
.Y(n_1844)
);

OA21x2_ASAP7_75t_L g1845 ( 
.A1(n_1766),
.A2(n_1734),
.B(n_1744),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1787),
.B(n_1745),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1801),
.B(n_1744),
.Y(n_1847)
);

OAI21x1_ASAP7_75t_L g1848 ( 
.A1(n_1824),
.A2(n_1703),
.B(n_1753),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1806),
.Y(n_1849)
);

NOR2x1_ASAP7_75t_R g1850 ( 
.A(n_1764),
.B(n_1708),
.Y(n_1850)
);

AO21x1_ASAP7_75t_L g1851 ( 
.A1(n_1791),
.A2(n_1699),
.B(n_1664),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1772),
.A2(n_1714),
.B(n_1701),
.Y(n_1852)
);

OA21x2_ASAP7_75t_L g1853 ( 
.A1(n_1805),
.A2(n_1699),
.B(n_1664),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1816),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1775),
.A2(n_1669),
.B1(n_1661),
.B2(n_1748),
.Y(n_1855)
);

A2O1A1Ixp33_ASAP7_75t_L g1856 ( 
.A1(n_1802),
.A2(n_1669),
.B(n_1664),
.C(n_398),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1771),
.B(n_1669),
.Y(n_1857)
);

AOI21x1_ASAP7_75t_L g1858 ( 
.A1(n_1788),
.A2(n_396),
.B(n_397),
.Y(n_1858)
);

OAI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1814),
.A2(n_400),
.B(n_402),
.Y(n_1859)
);

CKINVDCx11_ASAP7_75t_R g1860 ( 
.A(n_1794),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1831),
.B(n_1806),
.Y(n_1861)
);

INVx3_ASAP7_75t_L g1862 ( 
.A(n_1831),
.Y(n_1862)
);

OR2x6_ASAP7_75t_L g1863 ( 
.A(n_1845),
.B(n_1827),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1831),
.Y(n_1864)
);

INVx3_ASAP7_75t_L g1865 ( 
.A(n_1831),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1829),
.Y(n_1866)
);

HB1xp67_ASAP7_75t_L g1867 ( 
.A(n_1829),
.Y(n_1867)
);

BUFx6f_ASAP7_75t_L g1868 ( 
.A(n_1858),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1835),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1835),
.Y(n_1870)
);

OAI21x1_ASAP7_75t_L g1871 ( 
.A1(n_1840),
.A2(n_1760),
.B(n_1817),
.Y(n_1871)
);

INVx2_ASAP7_75t_SL g1872 ( 
.A(n_1846),
.Y(n_1872)
);

AO21x2_ASAP7_75t_L g1873 ( 
.A1(n_1851),
.A2(n_1780),
.B(n_1765),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1852),
.B(n_1809),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1841),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1839),
.Y(n_1876)
);

AO21x2_ASAP7_75t_L g1877 ( 
.A1(n_1851),
.A2(n_1767),
.B(n_1768),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1838),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1838),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1853),
.Y(n_1880)
);

INVx2_ASAP7_75t_SL g1881 ( 
.A(n_1846),
.Y(n_1881)
);

INVx3_ASAP7_75t_L g1882 ( 
.A(n_1840),
.Y(n_1882)
);

OAI211xp5_ASAP7_75t_L g1883 ( 
.A1(n_1874),
.A2(n_1844),
.B(n_1826),
.C(n_1834),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1877),
.A2(n_1873),
.B1(n_1874),
.B2(n_1859),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1863),
.A2(n_1782),
.B1(n_1800),
.B2(n_1856),
.Y(n_1885)
);

BUFx2_ASAP7_75t_L g1886 ( 
.A(n_1875),
.Y(n_1886)
);

OAI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1863),
.A2(n_1782),
.B1(n_1793),
.B2(n_1845),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1875),
.B(n_1830),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1872),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1872),
.B(n_1881),
.Y(n_1890)
);

HB1xp67_ASAP7_75t_L g1891 ( 
.A(n_1866),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1878),
.Y(n_1892)
);

OAI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1863),
.A2(n_1845),
.B1(n_1847),
.B2(n_1843),
.Y(n_1893)
);

OAI21xp33_ASAP7_75t_L g1894 ( 
.A1(n_1863),
.A2(n_1830),
.B(n_1832),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1878),
.Y(n_1895)
);

AOI221xp5_ASAP7_75t_L g1896 ( 
.A1(n_1877),
.A2(n_1783),
.B1(n_1854),
.B2(n_1774),
.C(n_1832),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1863),
.A2(n_1855),
.B1(n_1833),
.B2(n_1810),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1872),
.B(n_1854),
.Y(n_1898)
);

OAI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1871),
.A2(n_1848),
.B(n_1788),
.Y(n_1899)
);

INVx3_ASAP7_75t_L g1900 ( 
.A(n_1892),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1891),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1891),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1898),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1890),
.B(n_1881),
.Y(n_1904)
);

NOR2x1_ASAP7_75t_L g1905 ( 
.A(n_1886),
.B(n_1789),
.Y(n_1905)
);

INVx3_ASAP7_75t_L g1906 ( 
.A(n_1888),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1889),
.B(n_1881),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1903),
.B(n_1877),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1901),
.Y(n_1909)
);

INVxp67_ASAP7_75t_SL g1910 ( 
.A(n_1905),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1906),
.B(n_1877),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1906),
.B(n_1896),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1909),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1910),
.B(n_1900),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1908),
.Y(n_1915)
);

OAI31xp33_ASAP7_75t_L g1916 ( 
.A1(n_1912),
.A2(n_1883),
.A3(n_1887),
.B(n_1884),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1911),
.B(n_1900),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1910),
.B(n_1900),
.Y(n_1918)
);

NOR2x1p5_ASAP7_75t_L g1919 ( 
.A(n_1913),
.B(n_1850),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1914),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1915),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1921),
.Y(n_1922)
);

BUFx2_ASAP7_75t_L g1923 ( 
.A(n_1920),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1923),
.Y(n_1924)
);

CKINVDCx14_ASAP7_75t_R g1925 ( 
.A(n_1924),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1925),
.Y(n_1926)
);

OAI21xp33_ASAP7_75t_L g1927 ( 
.A1(n_1925),
.A2(n_1920),
.B(n_1922),
.Y(n_1927)
);

AOI222xp33_ASAP7_75t_L g1928 ( 
.A1(n_1927),
.A2(n_1923),
.B1(n_1926),
.B2(n_1914),
.C1(n_1918),
.C2(n_1917),
.Y(n_1928)
);

NAND3xp33_ASAP7_75t_L g1929 ( 
.A(n_1926),
.B(n_1916),
.C(n_1918),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1928),
.Y(n_1930)
);

AOI322xp5_ASAP7_75t_L g1931 ( 
.A1(n_1929),
.A2(n_1917),
.A3(n_1893),
.B1(n_1894),
.B2(n_1864),
.C1(n_1861),
.C2(n_1865),
.Y(n_1931)
);

AOI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1929),
.A2(n_1893),
.B1(n_1885),
.B2(n_1864),
.C(n_1899),
.Y(n_1932)
);

INVx1_ASAP7_75t_SL g1933 ( 
.A(n_1930),
.Y(n_1933)
);

NOR3xp33_ASAP7_75t_L g1934 ( 
.A(n_1932),
.B(n_1850),
.C(n_1860),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1931),
.A2(n_1919),
.B1(n_1897),
.B2(n_1901),
.Y(n_1935)
);

XOR2x2_ASAP7_75t_L g1936 ( 
.A(n_1933),
.B(n_1815),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1934),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1935),
.Y(n_1938)
);

INVxp67_ASAP7_75t_SL g1939 ( 
.A(n_1933),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1933),
.A2(n_1873),
.B1(n_1865),
.B2(n_1862),
.Y(n_1940)
);

OAI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1935),
.A2(n_1902),
.B1(n_1907),
.B2(n_1904),
.Y(n_1941)
);

BUFx2_ASAP7_75t_L g1942 ( 
.A(n_1933),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1942),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1939),
.Y(n_1944)
);

NOR2x1_ASAP7_75t_L g1945 ( 
.A(n_1938),
.B(n_1941),
.Y(n_1945)
);

INVx2_ASAP7_75t_SL g1946 ( 
.A(n_1936),
.Y(n_1946)
);

NOR2xp67_ASAP7_75t_L g1947 ( 
.A(n_1937),
.B(n_1940),
.Y(n_1947)
);

AO22x1_ASAP7_75t_L g1948 ( 
.A1(n_1939),
.A2(n_1902),
.B1(n_1895),
.B2(n_1812),
.Y(n_1948)
);

NOR2x1_ASAP7_75t_L g1949 ( 
.A(n_1942),
.B(n_1803),
.Y(n_1949)
);

NOR2x1_ASAP7_75t_L g1950 ( 
.A(n_1942),
.B(n_1822),
.Y(n_1950)
);

OAI22x1_ASAP7_75t_L g1951 ( 
.A1(n_1942),
.A2(n_1813),
.B1(n_1812),
.B2(n_1821),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1942),
.Y(n_1952)
);

INVxp67_ASAP7_75t_SL g1953 ( 
.A(n_1952),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1949),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1943),
.B(n_1862),
.Y(n_1955)
);

INVxp67_ASAP7_75t_L g1956 ( 
.A(n_1945),
.Y(n_1956)
);

NAND2x1p5_ASAP7_75t_L g1957 ( 
.A(n_1944),
.B(n_1807),
.Y(n_1957)
);

NAND4xp75_ASAP7_75t_L g1958 ( 
.A(n_1947),
.B(n_1843),
.C(n_1760),
.D(n_1857),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1950),
.Y(n_1959)
);

AOI22xp5_ASAP7_75t_SL g1960 ( 
.A1(n_1946),
.A2(n_1798),
.B1(n_1807),
.B2(n_1843),
.Y(n_1960)
);

HB1xp67_ASAP7_75t_L g1961 ( 
.A(n_1948),
.Y(n_1961)
);

NOR2x1_ASAP7_75t_L g1962 ( 
.A(n_1951),
.B(n_1798),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1952),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1952),
.Y(n_1964)
);

NOR3xp33_ASAP7_75t_L g1965 ( 
.A(n_1952),
.B(n_1858),
.C(n_1862),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1952),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1952),
.Y(n_1967)
);

XNOR2x1_ASAP7_75t_L g1968 ( 
.A(n_1945),
.B(n_1770),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1952),
.B(n_1857),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1952),
.B(n_1866),
.Y(n_1970)
);

AND2x2_ASAP7_75t_SL g1971 ( 
.A(n_1943),
.B(n_1807),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1952),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1952),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1944),
.B(n_1862),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1952),
.Y(n_1975)
);

AND3x4_ASAP7_75t_L g1976 ( 
.A(n_1945),
.B(n_1784),
.C(n_1836),
.Y(n_1976)
);

NOR2x1_ASAP7_75t_SL g1977 ( 
.A(n_1952),
.B(n_1873),
.Y(n_1977)
);

NOR2x1_ASAP7_75t_L g1978 ( 
.A(n_1943),
.B(n_1873),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1956),
.Y(n_1979)
);

NOR2x1_ASAP7_75t_L g1980 ( 
.A(n_1966),
.B(n_1863),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1953),
.Y(n_1981)
);

AOI221xp5_ASAP7_75t_L g1982 ( 
.A1(n_1961),
.A2(n_1868),
.B1(n_1865),
.B2(n_1862),
.C(n_1861),
.Y(n_1982)
);

AOI221xp5_ASAP7_75t_L g1983 ( 
.A1(n_1959),
.A2(n_1868),
.B1(n_1865),
.B2(n_1861),
.C(n_1880),
.Y(n_1983)
);

AOI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1954),
.A2(n_1843),
.B1(n_1868),
.B2(n_1865),
.Y(n_1984)
);

OAI21xp33_ASAP7_75t_L g1985 ( 
.A1(n_1963),
.A2(n_1882),
.B(n_1879),
.Y(n_1985)
);

AOI21xp33_ASAP7_75t_L g1986 ( 
.A1(n_1971),
.A2(n_405),
.B(n_408),
.Y(n_1986)
);

AOI211x1_ASAP7_75t_L g1987 ( 
.A1(n_1964),
.A2(n_1879),
.B(n_1870),
.C(n_1869),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1975),
.A2(n_1868),
.B(n_1837),
.Y(n_1988)
);

AOI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1965),
.A2(n_1868),
.B1(n_1880),
.B2(n_1840),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1968),
.B(n_1868),
.Y(n_1990)
);

OAI22xp33_ASAP7_75t_L g1991 ( 
.A1(n_1955),
.A2(n_1868),
.B1(n_1797),
.B2(n_1837),
.Y(n_1991)
);

NOR4xp75_ASAP7_75t_L g1992 ( 
.A(n_1970),
.B(n_1790),
.C(n_1882),
.D(n_1799),
.Y(n_1992)
);

AOI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1976),
.A2(n_1880),
.B1(n_1840),
.B2(n_1842),
.Y(n_1993)
);

AOI21xp5_ASAP7_75t_L g1994 ( 
.A1(n_1967),
.A2(n_1837),
.B(n_1867),
.Y(n_1994)
);

NOR4xp25_ASAP7_75t_L g1995 ( 
.A(n_1972),
.B(n_1973),
.C(n_1974),
.D(n_1957),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1969),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1977),
.B(n_1842),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1969),
.A2(n_1837),
.B(n_1867),
.Y(n_1998)
);

XOR2xp5_ASAP7_75t_L g1999 ( 
.A(n_1962),
.B(n_409),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1978),
.B(n_1797),
.Y(n_2000)
);

AO22x2_ASAP7_75t_L g2001 ( 
.A1(n_1958),
.A2(n_1847),
.B1(n_1784),
.B2(n_1836),
.Y(n_2001)
);

OAI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1960),
.A2(n_1778),
.B1(n_1870),
.B2(n_1869),
.Y(n_2002)
);

AOI211xp5_ASAP7_75t_SL g2003 ( 
.A1(n_1956),
.A2(n_1882),
.B(n_1811),
.C(n_1836),
.Y(n_2003)
);

AOI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1961),
.A2(n_1776),
.B1(n_1842),
.B2(n_1848),
.Y(n_2004)
);

INVxp67_ASAP7_75t_SL g2005 ( 
.A(n_1981),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1979),
.Y(n_2006)
);

NAND3x1_ASAP7_75t_L g2007 ( 
.A(n_1996),
.B(n_1995),
.C(n_2000),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1999),
.Y(n_2008)
);

BUFx3_ASAP7_75t_L g2009 ( 
.A(n_1990),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1980),
.B(n_1849),
.Y(n_2010)
);

NOR2x1p5_ASAP7_75t_L g2011 ( 
.A(n_1997),
.B(n_1882),
.Y(n_2011)
);

INVx4_ASAP7_75t_L g2012 ( 
.A(n_2001),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1987),
.Y(n_2013)
);

CKINVDCx20_ASAP7_75t_R g2014 ( 
.A(n_1986),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1993),
.B(n_410),
.Y(n_2015)
);

INVx5_ASAP7_75t_L g2016 ( 
.A(n_1992),
.Y(n_2016)
);

AOI211xp5_ASAP7_75t_L g2017 ( 
.A1(n_1985),
.A2(n_1871),
.B(n_1828),
.C(n_1849),
.Y(n_2017)
);

XNOR2x1_ASAP7_75t_L g2018 ( 
.A(n_2001),
.B(n_2002),
.Y(n_2018)
);

XOR2x1_ASAP7_75t_L g2019 ( 
.A(n_1991),
.B(n_1776),
.Y(n_2019)
);

INVx3_ASAP7_75t_L g2020 ( 
.A(n_2003),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1988),
.Y(n_2021)
);

OAI22xp5_ASAP7_75t_SL g2022 ( 
.A1(n_2004),
.A2(n_1797),
.B1(n_1845),
.B2(n_1836),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1994),
.B(n_1849),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1984),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_2005),
.B(n_1982),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2006),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2012),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_2007),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_2014),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_2013),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_2020),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2018),
.Y(n_2032)
);

AOI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_2008),
.A2(n_1983),
.B1(n_1998),
.B2(n_1989),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_2021),
.A2(n_1828),
.B(n_1871),
.Y(n_2034)
);

AND3x2_ASAP7_75t_L g2035 ( 
.A(n_2024),
.B(n_411),
.C(n_416),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_2016),
.Y(n_2036)
);

OR3x2_ASAP7_75t_L g2037 ( 
.A(n_2027),
.B(n_2009),
.C(n_2016),
.Y(n_2037)
);

OAI22xp5_ASAP7_75t_SL g2038 ( 
.A1(n_2036),
.A2(n_2015),
.B1(n_2023),
.B2(n_2010),
.Y(n_2038)
);

INVx2_ASAP7_75t_SL g2039 ( 
.A(n_2028),
.Y(n_2039)
);

XNOR2xp5_ASAP7_75t_L g2040 ( 
.A(n_2032),
.B(n_2029),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_2028),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_2031),
.B(n_2026),
.Y(n_2042)
);

OAI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_2030),
.A2(n_2017),
.B(n_2019),
.Y(n_2043)
);

XOR2xp5_ASAP7_75t_L g2044 ( 
.A(n_2033),
.B(n_2011),
.Y(n_2044)
);

AOI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_2040),
.A2(n_2025),
.B(n_2034),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_2037),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2039),
.B(n_2035),
.Y(n_2047)
);

NAND3xp33_ASAP7_75t_L g2048 ( 
.A(n_2041),
.B(n_2022),
.C(n_418),
.Y(n_2048)
);

OAI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_2044),
.A2(n_1882),
.B1(n_1761),
.B2(n_1876),
.Y(n_2049)
);

OAI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_2046),
.A2(n_2042),
.B1(n_2043),
.B2(n_2038),
.Y(n_2050)
);

OAI21x1_ASAP7_75t_SL g2051 ( 
.A1(n_2045),
.A2(n_2047),
.B(n_2048),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2049),
.Y(n_2052)
);

AO22x2_ASAP7_75t_L g2053 ( 
.A1(n_2046),
.A2(n_417),
.B1(n_421),
.B2(n_422),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_2050),
.B(n_423),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_SL g2055 ( 
.A1(n_2052),
.A2(n_424),
.B1(n_425),
.B2(n_429),
.Y(n_2055)
);

AOI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_2054),
.A2(n_2053),
.B1(n_2051),
.B2(n_1761),
.Y(n_2056)
);

AOI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_2055),
.A2(n_430),
.B(n_431),
.Y(n_2057)
);

AOI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_2057),
.A2(n_432),
.B(n_435),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2056),
.Y(n_2059)
);

AOI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_2057),
.A2(n_438),
.B(n_440),
.Y(n_2060)
);

AOI22xp5_ASAP7_75t_SL g2061 ( 
.A1(n_2059),
.A2(n_444),
.B1(n_448),
.B2(n_450),
.Y(n_2061)
);

AOI222xp33_ASAP7_75t_L g2062 ( 
.A1(n_2058),
.A2(n_452),
.B1(n_453),
.B2(n_454),
.C1(n_456),
.C2(n_460),
.Y(n_2062)
);

OR2x6_ASAP7_75t_L g2063 ( 
.A(n_2061),
.B(n_2060),
.Y(n_2063)
);

NAND4xp75_ASAP7_75t_L g2064 ( 
.A(n_2063),
.B(n_2062),
.C(n_463),
.D(n_465),
.Y(n_2064)
);

AOI211xp5_ASAP7_75t_L g2065 ( 
.A1(n_2064),
.A2(n_461),
.B(n_466),
.C(n_467),
.Y(n_2065)
);


endmodule