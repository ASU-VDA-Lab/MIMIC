module fake_jpeg_14703_n_297 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_155;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_34),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_51),
.Y(n_63)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_29),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_58),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_25),
.B1(n_28),
.B2(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_56),
.B1(n_62),
.B2(n_26),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_25),
.B1(n_32),
.B2(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_25),
.B1(n_32),
.B2(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_71),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_66),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_20),
.C(n_39),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_68),
.B(n_92),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_76),
.Y(n_99)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_35),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_54),
.C(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_86),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_41),
.B(n_17),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_74),
.B(n_22),
.C(n_30),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_20),
.C(n_39),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_36),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_20),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_0),
.Y(n_123)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_85),
.Y(n_104)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_32),
.B1(n_28),
.B2(n_21),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_84),
.A2(n_97),
.B1(n_22),
.B2(n_30),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_35),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_94),
.Y(n_105)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_21),
.B1(n_26),
.B2(n_34),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_89),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_18),
.B1(n_36),
.B2(n_12),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_22),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_44),
.B(n_17),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_48),
.A2(n_30),
.B1(n_34),
.B2(n_33),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_18),
.B(n_26),
.C(n_33),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_106),
.A2(n_115),
.B(n_123),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_39),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_36),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_108),
.B(n_31),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_33),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_19),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_112),
.B(n_118),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_78),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_98),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_122),
.B1(n_93),
.B2(n_70),
.Y(n_132)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_31),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_86),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_71),
.B1(n_72),
.B2(n_67),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_127),
.A2(n_140),
.B1(n_148),
.B2(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_64),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_138),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_136),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_126),
.A2(n_82),
.B1(n_65),
.B2(n_75),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_135),
.A2(n_110),
.B1(n_116),
.B2(n_114),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_81),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_77),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_142),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_69),
.B1(n_88),
.B2(n_83),
.Y(n_140)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_66),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_145),
.B(n_155),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_75),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_85),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_106),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_95),
.C(n_79),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_127),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_100),
.B(n_23),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_146),
.B(n_109),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_147),
.B(n_153),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_99),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_79),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_152),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_19),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_119),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_0),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_123),
.B(n_100),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_157),
.B(n_160),
.Y(n_208)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_99),
.B1(n_102),
.B2(n_111),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_159),
.A2(n_164),
.B1(n_128),
.B2(n_155),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_143),
.A2(n_115),
.B1(n_120),
.B2(n_116),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_170),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_149),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_173),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_174),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_136),
.B(n_109),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_179),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_139),
.B(n_146),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_141),
.B(n_121),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_114),
.B(n_110),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_182),
.B(n_183),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_0),
.B(n_1),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_142),
.B(n_24),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_121),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_185),
.Y(n_201)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_187),
.Y(n_192)
);

AOI22x1_ASAP7_75t_SL g188 ( 
.A1(n_185),
.A2(n_141),
.B1(n_154),
.B2(n_156),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_188),
.A2(n_202),
.B(n_207),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_178),
.B1(n_186),
.B2(n_174),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_197),
.B1(n_206),
.B2(n_210),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_150),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_195),
.B(n_209),
.Y(n_220)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_156),
.B1(n_141),
.B2(n_128),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_164),
.Y(n_225)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_133),
.B1(n_131),
.B2(n_154),
.Y(n_206)
);

XOR2x2_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_145),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_181),
.A2(n_121),
.B1(n_119),
.B2(n_24),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_161),
.A2(n_0),
.B(n_1),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_183),
.B(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_212),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_175),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_203),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_168),
.B1(n_162),
.B2(n_169),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_201),
.B1(n_190),
.B2(n_189),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_176),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_222),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_170),
.C(n_159),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_224),
.C(n_228),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_172),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_162),
.C(n_166),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_230),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_208),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_192),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_161),
.C(n_182),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_171),
.Y(n_229)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_179),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_231),
.A2(n_201),
.B1(n_200),
.B2(n_199),
.Y(n_234)
);

OAI322xp33_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_184),
.A3(n_160),
.B1(n_157),
.B2(n_163),
.C1(n_19),
.C2(n_7),
.Y(n_232)
);

NOR3xp33_ASAP7_75t_SL g233 ( 
.A(n_232),
.B(n_10),
.C(n_13),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_239),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_223),
.B(n_230),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_235),
.B(n_236),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_217),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_237),
.A2(n_214),
.B1(n_191),
.B2(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_218),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_241),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_242),
.B(n_248),
.Y(n_251)
);

O2A1O1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_244),
.A2(n_213),
.B(n_211),
.C(n_241),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_198),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_210),
.C(n_2),
.Y(n_260)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_246),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_233),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_234),
.A2(n_231),
.B(n_202),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_252),
.A2(n_254),
.B(n_261),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_272)
);

AOI322xp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_226),
.A3(n_223),
.B1(n_225),
.B2(n_189),
.C1(n_222),
.C2(n_224),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_243),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_244),
.A2(n_228),
.B1(n_184),
.B2(n_219),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_257),
.A2(n_254),
.B1(n_260),
.B2(n_261),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_259),
.C(n_252),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_1),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_266),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_262),
.C(n_257),
.Y(n_274)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_243),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_268),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_245),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_245),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_270),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_9),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_261),
.A2(n_9),
.B1(n_14),
.B2(n_4),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_255),
.B1(n_10),
.B2(n_6),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_264),
.C(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_279),
.B1(n_14),
.B2(n_15),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_265),
.Y(n_283)
);

NOR2x1_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_6),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_7),
.B(n_13),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_271),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_283),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_270),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_275),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_SL g292 ( 
.A(n_286),
.B(n_287),
.C(n_288),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_286),
.A2(n_279),
.B(n_280),
.C(n_282),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_2),
.B(n_3),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_L g293 ( 
.A1(n_291),
.A2(n_287),
.B(n_274),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_294),
.C(n_295),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g294 ( 
.A(n_289),
.B(n_15),
.CI(n_2),
.CON(n_294),
.SN(n_294)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_292),
.Y(n_297)
);


endmodule