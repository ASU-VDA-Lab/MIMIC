module fake_jpeg_8969_n_191 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_191);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_SL g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_30),
.Y(n_47)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_13),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_34),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_14),
.B1(n_13),
.B2(n_23),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_45),
.B1(n_21),
.B2(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_48),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_14),
.B1(n_18),
.B2(n_12),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_44),
.B1(n_33),
.B2(n_32),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_32),
.B(n_26),
.C(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_30),
.A2(n_18),
.B1(n_12),
.B2(n_15),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_24),
.B1(n_21),
.B2(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_65),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_20),
.B1(n_35),
.B2(n_6),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_27),
.B1(n_26),
.B2(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_27),
.B1(n_1),
.B2(n_3),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_11),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_25),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_11),
.B1(n_1),
.B2(n_5),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_28),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_25),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_43),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_0),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_35),
.C(n_37),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_79),
.C(n_60),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_40),
.B1(n_39),
.B2(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_53),
.Y(n_85)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_38),
.B1(n_37),
.B2(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_81),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_25),
.C(n_29),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_50),
.A2(n_46),
.B1(n_49),
.B2(n_6),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_54),
.B(n_5),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_95),
.B(n_99),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_98),
.C(n_66),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_55),
.B(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_75),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_70),
.C(n_79),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_93),
.A2(n_76),
.B1(n_69),
.B2(n_74),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_93),
.B1(n_84),
.B2(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_109),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_78),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_66),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_114),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_77),
.C(n_71),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_95),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_71),
.B(n_65),
.C(n_77),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_125),
.B1(n_106),
.B2(n_100),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_120),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_122),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_87),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_124),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_99),
.CI(n_84),
.CON(n_124),
.SN(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_94),
.B(n_19),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_6),
.Y(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_83),
.B1(n_88),
.B2(n_92),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_100),
.B1(n_111),
.B2(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_136),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_137),
.B1(n_139),
.B2(n_142),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_128),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_110),
.B1(n_102),
.B2(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_65),
.B1(n_46),
.B2(n_49),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_125),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_140),
.B(n_130),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_83),
.B1(n_29),
.B2(n_28),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_136),
.A2(n_129),
.B1(n_117),
.B2(n_124),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_149),
.B1(n_16),
.B2(n_29),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_130),
.C(n_122),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_141),
.C(n_132),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_124),
.B1(n_120),
.B2(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_154),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_126),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_139),
.Y(n_158)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_83),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_0),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_160),
.C(n_162),
.Y(n_166)
);

FAx1_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_144),
.CI(n_142),
.CON(n_157),
.SN(n_157)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_159),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_19),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_152),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_147),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_28),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_147),
.C(n_148),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_171),
.C(n_157),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_170),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_153),
.C(n_150),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_153),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_157),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_176),
.A2(n_178),
.B(n_7),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_16),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_166),
.B(n_7),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_179),
.B(n_181),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_182),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_174),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_34),
.C(n_8),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_187),
.B1(n_184),
.B2(n_10),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_188),
.B(n_183),
.Y(n_189)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_0),
.B(n_34),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_16),
.Y(n_191)
);


endmodule