module fake_jpeg_30811_n_154 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_35),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_23),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_71),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_0),
.CON(n_71),
.SN(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_72),
.B(n_53),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_76),
.B1(n_80),
.B2(n_86),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_85),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_50),
.B1(n_55),
.B2(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_64),
.B1(n_57),
.B2(n_47),
.Y(n_80)
);

CKINVDCx9p33_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_65),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_58),
.B1(n_47),
.B2(n_48),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_68),
.B(n_77),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_2),
.B(n_4),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_67),
.B1(n_48),
.B2(n_49),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_116)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_82),
.B1(n_54),
.B2(n_61),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_97),
.A2(n_52),
.B1(n_3),
.B2(n_4),
.Y(n_103)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_1),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_5),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_107),
.B1(n_109),
.B2(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_7),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_95),
.B1(n_93),
.B2(n_101),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_22),
.B1(n_41),
.B2(n_40),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_114),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_19),
.B1(n_39),
.B2(n_38),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_9),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_117),
.B1(n_9),
.B2(n_10),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_42),
.B1(n_16),
.B2(n_24),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_87),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_8),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_99),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_121),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_123),
.B(n_127),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_132),
.B1(n_113),
.B2(n_112),
.Y(n_136)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_131),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_10),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_129),
.B(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_11),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_11),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_118),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_137),
.C(n_125),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_122),
.C(n_123),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_27),
.B(n_36),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_124),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_141),
.B(n_143),
.Y(n_146)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_134),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_146),
.B(n_139),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_138),
.B1(n_145),
.B2(n_140),
.Y(n_148)
);

OAI321xp33_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_142),
.A3(n_144),
.B1(n_133),
.B2(n_15),
.C(n_25),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_30),
.B(n_31),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g152 ( 
.A(n_151),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_32),
.C1(n_37),
.C2(n_150),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_12),
.Y(n_154)
);


endmodule