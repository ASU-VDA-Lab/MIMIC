module fake_jpeg_29577_n_219 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_1),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_19),
.Y(n_67)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_27),
.B1(n_16),
.B2(n_23),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_64),
.B1(n_18),
.B2(n_26),
.Y(n_83)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_21),
.B1(n_16),
.B2(n_23),
.Y(n_76)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_66),
.Y(n_73)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_24),
.B1(n_18),
.B2(n_22),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_22),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_67),
.B(n_71),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_68),
.B(n_86),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_77),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_48),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_29),
.B1(n_26),
.B2(n_20),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_82),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_24),
.C(n_29),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_87),
.C(n_92),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_76),
.A2(n_83),
.B1(n_88),
.B2(n_94),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_19),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_27),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_27),
.B1(n_23),
.B2(n_21),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_85),
.A2(n_91),
.B(n_87),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_23),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_21),
.C(n_16),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_30),
.B1(n_21),
.B2(n_16),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_16),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_60),
.B(n_30),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_59),
.C(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_54),
.A2(n_59),
.B1(n_63),
.B2(n_5),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_2),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_4),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_4),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_15),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_15),
.C(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_4),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_82),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_123),
.Y(n_137)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_121),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_99),
.B(n_97),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_132),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_74),
.B(n_86),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_113),
.B(n_117),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_76),
.B1(n_82),
.B2(n_91),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_146),
.B1(n_118),
.B2(n_116),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_99),
.B(n_75),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_92),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_134),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_90),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_90),
.B1(n_78),
.B2(n_95),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_115),
.C(n_113),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_152),
.C(n_157),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_129),
.B(n_125),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_101),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_153),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_135),
.B1(n_145),
.B2(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_111),
.C(n_100),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_98),
.A3(n_103),
.B1(n_112),
.B2(n_78),
.C1(n_105),
.C2(n_110),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_120),
.C(n_98),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_121),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_158),
.B(n_159),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_5),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_96),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_6),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_164),
.B(n_6),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_142),
.B(n_130),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_128),
.B(n_7),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_178),
.B1(n_138),
.B2(n_141),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_173),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_131),
.B1(n_146),
.B2(n_125),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_138),
.B1(n_141),
.B2(n_128),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_164),
.B(n_134),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_176),
.A2(n_148),
.B(n_160),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_137),
.B1(n_129),
.B2(n_145),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_179),
.A2(n_156),
.B1(n_150),
.B2(n_155),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_189),
.B(n_184),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_167),
.A2(n_157),
.B(n_161),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_186),
.B(n_191),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_183),
.Y(n_195)
);

OAI322xp33_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_155),
.A3(n_152),
.B1(n_136),
.B2(n_154),
.C1(n_163),
.C2(n_151),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_166),
.B1(n_179),
.B2(n_174),
.Y(n_193)
);

INVxp33_ASAP7_75t_SL g186 ( 
.A(n_177),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_170),
.B(n_139),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_175),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_176),
.C(n_171),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_175),
.C(n_165),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_190),
.B1(n_6),
.B2(n_7),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_193),
.A2(n_185),
.B1(n_188),
.B2(n_191),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_168),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_13),
.C(n_10),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_180),
.A2(n_174),
.B(n_165),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_197),
.A2(n_200),
.B1(n_7),
.B2(n_8),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_198),
.B(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_204),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_203),
.A2(n_196),
.B1(n_199),
.B2(n_197),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_195),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_192),
.B(n_13),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_206),
.B(n_207),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_194),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_211),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_205),
.A2(n_9),
.B(n_11),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_212),
.B(n_210),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_213),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_201),
.B(n_207),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_217),
.B1(n_203),
.B2(n_11),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_12),
.Y(n_219)
);


endmodule