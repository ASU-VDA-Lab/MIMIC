module fake_jpeg_31741_n_192 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_192);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_30),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_55),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_18),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_62),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_18),
.B1(n_31),
.B2(n_29),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_19),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_32),
.C(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_16),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_68),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_41),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_71),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_51),
.B1(n_45),
.B2(n_34),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_69),
.A2(n_17),
.B1(n_5),
.B2(n_4),
.Y(n_115)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_32),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_73),
.B(n_87),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_22),
.B1(n_31),
.B2(n_25),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_80),
.B1(n_83),
.B2(n_84),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_22),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_92),
.B1(n_0),
.B2(n_1),
.Y(n_103)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_81),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_26),
.B1(n_16),
.B2(n_2),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_8),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_16),
.B1(n_17),
.B2(n_3),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_10),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_17),
.B1(n_1),
.B2(n_3),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_46),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_56),
.B1(n_59),
.B2(n_65),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_90),
.B1(n_75),
.B2(n_70),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_65),
.B1(n_17),
.B2(n_3),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_71),
.B1(n_66),
.B2(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_0),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_0),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_17),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_111),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_83),
.B1(n_74),
.B2(n_80),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_116),
.B(n_119),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_66),
.B(n_76),
.C(n_68),
.D(n_67),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_104),
.B(n_115),
.C(n_105),
.D(n_93),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_107),
.B(n_106),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_131),
.B(n_97),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_133),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_66),
.B(n_71),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_67),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_134),
.B(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_139),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_140),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_100),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_121),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_144),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_106),
.B(n_113),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_148),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_113),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_104),
.B1(n_127),
.B2(n_124),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_161),
.B1(n_145),
.B2(n_143),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_130),
.C(n_131),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_159),
.C(n_144),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_117),
.A3(n_132),
.B1(n_133),
.B2(n_129),
.C1(n_122),
.C2(n_120),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_148),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_132),
.C(n_120),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_142),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_163),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_136),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_136),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_166),
.C(n_168),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_153),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_169),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_142),
.C(n_143),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_145),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_168),
.A2(n_152),
.B(n_157),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_161),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_154),
.B(n_155),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_177),
.Y(n_180)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_164),
.C(n_151),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_179),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_94),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_182),
.B(n_13),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_174),
.B(n_15),
.Y(n_182)
);

AOI21x1_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_13),
.B(n_14),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_174),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_185),
.B(n_186),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_173),
.B1(n_94),
.B2(n_82),
.Y(n_186)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_4),
.B(n_5),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_185),
.C(n_183),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_190),
.B(n_4),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_90),
.B(n_173),
.Y(n_192)
);


endmodule