module fake_ibex_2019_n_1101 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1101);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1101;

wire n_1084;
wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_177;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_1080;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_991;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1044;
wire n_1018;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_1077;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_317;
wire n_280;
wire n_340;
wire n_708;
wire n_375;
wire n_901;
wire n_1096;
wire n_187;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_1056;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_158;
wire n_1029;
wire n_859;
wire n_259;
wire n_276;
wire n_470;
wire n_339;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1053;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_1055;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1057;
wire n_1068;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_694;
wire n_523;
wire n_787;
wire n_977;
wire n_1075;
wire n_719;
wire n_370;
wire n_614;
wire n_431;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_1081;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_1001;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_1020;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_580;
wire n_483;
wire n_420;
wire n_487;
wire n_769;
wire n_1082;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_1089;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_167;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_1038;
wire n_999;
wire n_1092;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1062;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_433;
wire n_299;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_1063;
wire n_351;
wire n_456;
wire n_368;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1100;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_554;
wire n_553;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_1049;
wire n_1086;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_444;
wire n_562;
wire n_564;
wire n_506;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_706;
wire n_624;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_615;
wire n_512;
wire n_950;
wire n_685;
wire n_1026;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_894;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_712;
wire n_702;
wire n_451;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_817;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_1073;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_379;
wire n_320;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_172;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_1085;
wire n_361;
wire n_1095;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_195;
wire n_885;
wire n_588;
wire n_212;
wire n_513;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_912;
wire n_921;
wire n_874;
wire n_890;
wire n_1058;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_159;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_1035;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

INVxp67_ASAP7_75t_SL g157 ( 
.A(n_117),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_97),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_78),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_41),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_26),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_13),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_64),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_82),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_69),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_66),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_14),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g173 ( 
.A(n_48),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_76),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_84),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_52),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_6),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_63),
.Y(n_181)
);

INVxp33_ASAP7_75t_SL g182 ( 
.A(n_98),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_65),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_14),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_32),
.Y(n_187)
);

INVxp33_ASAP7_75t_SL g188 ( 
.A(n_6),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_16),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_25),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_39),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_7),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_3),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_47),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g198 ( 
.A(n_61),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_56),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_40),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_15),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_141),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_38),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_21),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_17),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_79),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_45),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_67),
.Y(n_210)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_94),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_20),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_4),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_25),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_58),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_124),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_22),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_116),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_93),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_70),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_44),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_118),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_42),
.Y(n_227)
);

INVxp33_ASAP7_75t_SL g228 ( 
.A(n_33),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_54),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_0),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_125),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_72),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_145),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_123),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_73),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_121),
.Y(n_236)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_13),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_15),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_7),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_120),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_0),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_107),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_86),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_23),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_9),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_136),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_35),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_142),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_149),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_62),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_37),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_20),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_24),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_4),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_132),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_130),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_59),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_85),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_9),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_5),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_129),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_31),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_102),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_57),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_95),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_74),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_5),
.B(n_110),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_91),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_81),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_213),
.B(n_1),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_161),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_177),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_213),
.B(n_1),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_2),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_177),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_206),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_164),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_165),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_168),
.Y(n_280)
);

OA21x2_ASAP7_75t_L g281 ( 
.A1(n_183),
.A2(n_71),
.B(n_154),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_169),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_174),
.Y(n_283)
);

AND2x4_ASAP7_75t_L g284 ( 
.A(n_170),
.B(n_199),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_195),
.A2(n_3),
.B1(n_8),
.B2(n_10),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_183),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_165),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_165),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_176),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_165),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_259),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_184),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_241),
.B(n_8),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_193),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_184),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_259),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_170),
.B(n_10),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_199),
.B(n_11),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_220),
.B(n_11),
.Y(n_302)
);

NAND2xp33_ASAP7_75t_L g303 ( 
.A(n_185),
.B(n_156),
.Y(n_303)
);

NAND2xp33_ASAP7_75t_SL g304 ( 
.A(n_185),
.B(n_12),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_215),
.B(n_12),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_197),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_235),
.B(n_16),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_197),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_216),
.B(n_17),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_233),
.B(n_18),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_233),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_204),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_178),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_233),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_220),
.B(n_18),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_204),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_235),
.B(n_196),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_226),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_225),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_259),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_162),
.Y(n_321)
);

NAND2x1_ASAP7_75t_L g322 ( 
.A(n_259),
.B(n_19),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_166),
.B(n_19),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_226),
.B(n_21),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_163),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_179),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_225),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_181),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_189),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_191),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_172),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_194),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_200),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_263),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_269),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_203),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_208),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_167),
.B(n_22),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_209),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_212),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_263),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_180),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_186),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_267),
.B(n_23),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_217),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_218),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_219),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_192),
.B(n_244),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_221),
.Y(n_349)
);

AND2x6_ASAP7_75t_L g350 ( 
.A(n_222),
.B(n_223),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_227),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_232),
.Y(n_352)
);

CKINVDCx8_ASAP7_75t_R g353 ( 
.A(n_243),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_187),
.B(n_24),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_248),
.B(n_26),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_187),
.B(n_27),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_269),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_302),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_276),
.Y(n_359)
);

NAND2xp33_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_159),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_302),
.Y(n_361)
);

INVx4_ASAP7_75t_SL g362 ( 
.A(n_350),
.Y(n_362)
);

AND2x6_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_234),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_284),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_302),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_357),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_284),
.B(n_240),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_307),
.A2(n_238),
.B1(n_214),
.B2(n_252),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_277),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_284),
.B(n_202),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_317),
.Y(n_371)
);

NOR2x1p5_ASAP7_75t_L g372 ( 
.A(n_317),
.B(n_239),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_357),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_276),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_357),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_277),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_304),
.A2(n_237),
.B1(n_188),
.B2(n_236),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_315),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_276),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_323),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_291),
.B(n_207),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_278),
.B(n_246),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_348),
.B(n_230),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_324),
.B(n_245),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_307),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_297),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_159),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_325),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_271),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_331),
.B(n_239),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_278),
.B(n_247),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_325),
.Y(n_393)
);

NAND2x1p5_ASAP7_75t_L g394 ( 
.A(n_323),
.B(n_253),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_271),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_280),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_338),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_353),
.B(n_158),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_270),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_335),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_353),
.B(n_260),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_280),
.B(n_201),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_282),
.B(n_190),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_356),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_282),
.B(n_249),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_327),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_279),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_272),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_272),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_357),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_283),
.B(n_254),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_283),
.B(n_182),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_335),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_338),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_275),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_285),
.B(n_262),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_318),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_357),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_335),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_285),
.B(n_211),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_275),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_350),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_322),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_273),
.A2(n_188),
.B1(n_237),
.B2(n_228),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_290),
.B(n_190),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_287),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_355),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_279),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_279),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_279),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_290),
.B(n_182),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_318),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_350),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_287),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_295),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_313),
.B(n_228),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_322),
.Y(n_439)
);

NAND3xp33_ASAP7_75t_SL g440 ( 
.A(n_354),
.B(n_260),
.C(n_224),
.Y(n_440)
);

NAND2x1p5_ASAP7_75t_L g441 ( 
.A(n_355),
.B(n_250),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_295),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_298),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_356),
.B(n_224),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_298),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_306),
.Y(n_446)
);

INVx5_ASAP7_75t_L g447 ( 
.A(n_293),
.Y(n_447)
);

NAND2x1_ASAP7_75t_L g448 ( 
.A(n_350),
.B(n_313),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_279),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_350),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_286),
.A2(n_296),
.B1(n_160),
.B2(n_171),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_321),
.B(n_158),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_306),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_326),
.B(n_251),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_342),
.B(n_255),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_308),
.Y(n_456)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_293),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_308),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_326),
.B(n_256),
.Y(n_459)
);

AO21x2_ASAP7_75t_L g460 ( 
.A1(n_310),
.A2(n_257),
.B(n_268),
.Y(n_460)
);

OAI21xp33_ASAP7_75t_L g461 ( 
.A1(n_343),
.A2(n_261),
.B(n_266),
.Y(n_461)
);

INVx5_ASAP7_75t_L g462 ( 
.A(n_293),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_328),
.B(n_329),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_312),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_312),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_328),
.B(n_229),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_329),
.B(n_229),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_316),
.Y(n_468)
);

OAI221xp5_ASAP7_75t_L g469 ( 
.A1(n_305),
.A2(n_210),
.B1(n_173),
.B2(n_198),
.C(n_157),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_330),
.B(n_236),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_281),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_316),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_319),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_330),
.B(n_265),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_332),
.B(n_264),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_319),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_334),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_334),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_341),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_274),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_341),
.Y(n_481)
);

AO22x2_ASAP7_75t_L g482 ( 
.A1(n_274),
.A2(n_242),
.B1(n_160),
.B2(n_258),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_300),
.A2(n_258),
.B1(n_231),
.B2(n_205),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_301),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_288),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_332),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_333),
.B(n_269),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_345),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_484),
.B(n_333),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_396),
.Y(n_490)
);

OR2x6_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_309),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_396),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_389),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_471),
.A2(n_281),
.B(n_351),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_448),
.Y(n_495)
);

OR2x6_ASAP7_75t_L g496 ( 
.A(n_470),
.B(n_344),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_425),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_390),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_389),
.Y(n_499)
);

NAND2x1p5_ASAP7_75t_L g500 ( 
.A(n_463),
.B(n_281),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

BUFx4f_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_393),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_387),
.B(n_344),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_359),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_400),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_424),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_374),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_452),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_379),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_391),
.B(n_336),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_424),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_484),
.B(n_336),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_399),
.B(n_337),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_399),
.B(n_337),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_358),
.A2(n_346),
.B1(n_351),
.B2(n_349),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_471),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_437),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_378),
.B(n_339),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_384),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_395),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_453),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_465),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_405),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_405),
.B(n_339),
.Y(n_525)
);

CKINVDCx8_ASAP7_75t_R g526 ( 
.A(n_416),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_463),
.B(n_340),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_413),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_380),
.B(n_340),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_384),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_407),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_435),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_467),
.B(n_171),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_413),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_425),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_367),
.B(n_346),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_439),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_483),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_367),
.B(n_349),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_386),
.B(n_418),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_439),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_435),
.B(n_347),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_408),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_362),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_464),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_473),
.Y(n_546)
);

AND2x4_ASAP7_75t_SL g547 ( 
.A(n_402),
.B(n_205),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_363),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_363),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_418),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_468),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_362),
.Y(n_552)
);

INVx5_ASAP7_75t_L g553 ( 
.A(n_363),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_381),
.B(n_347),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_380),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_486),
.B(n_352),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_450),
.B(n_361),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_467),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_450),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_410),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_444),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_365),
.A2(n_352),
.B1(n_345),
.B2(n_303),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_456),
.Y(n_563)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_363),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_398),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_R g566 ( 
.A(n_398),
.B(n_440),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_488),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_414),
.B(n_281),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_381),
.B(n_397),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_433),
.B(n_231),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_456),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_419),
.Y(n_572)
);

AOI22x1_ASAP7_75t_L g573 ( 
.A1(n_369),
.A2(n_269),
.B1(n_314),
.B2(n_311),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_397),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_474),
.A2(n_422),
.B1(n_376),
.B2(n_383),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_371),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_411),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_417),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_423),
.Y(n_579)
);

AND2x4_ASAP7_75t_SL g580 ( 
.A(n_483),
.B(n_320),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_428),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_394),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_436),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_385),
.B(n_294),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_422),
.B(n_27),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_442),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_443),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_474),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_438),
.B(n_320),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_385),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_383),
.B(n_320),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_441),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_404),
.B(n_299),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_446),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_458),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_472),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_434),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_474),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_476),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_427),
.B(n_299),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_441),
.Y(n_602)
);

O2A1O1Ixp33_ASAP7_75t_L g603 ( 
.A1(n_469),
.A2(n_299),
.B(n_29),
.C(n_30),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_403),
.B(n_311),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_477),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_401),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_370),
.B(n_311),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_478),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_490),
.B(n_372),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_520),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_490),
.Y(n_611)
);

BUFx2_ASAP7_75t_SL g612 ( 
.A(n_492),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_492),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_588),
.Y(n_614)
);

INVx6_ASAP7_75t_L g615 ( 
.A(n_606),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_502),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_520),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_568),
.A2(n_494),
.B(n_517),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_514),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_588),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_515),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_582),
.B(n_593),
.Y(n_622)
);

BUFx4f_ASAP7_75t_L g623 ( 
.A(n_585),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_549),
.B(n_429),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_498),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_520),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_575),
.A2(n_368),
.B1(n_406),
.B2(n_382),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_519),
.Y(n_628)
);

BUFx2_ASAP7_75t_SL g629 ( 
.A(n_526),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_540),
.B(n_528),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_592),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_502),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_540),
.Y(n_633)
);

CKINVDCx8_ASAP7_75t_R g634 ( 
.A(n_498),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_530),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_540),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_549),
.B(n_364),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_530),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_517),
.A2(n_360),
.B(n_388),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_536),
.A2(n_474),
.B1(n_370),
.B2(n_440),
.Y(n_640)
);

NAND2x1p5_ASAP7_75t_L g641 ( 
.A(n_549),
.B(n_479),
.Y(n_641)
);

AOI21xp33_ASAP7_75t_L g642 ( 
.A1(n_603),
.A2(n_460),
.B(n_469),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_574),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_588),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_588),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_528),
.B(n_455),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_530),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_599),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_536),
.B(n_426),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_555),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_539),
.B(n_475),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_577),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_539),
.B(n_382),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_569),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_585),
.A2(n_461),
.B1(n_454),
.B2(n_392),
.Y(n_655)
);

A2O1A1Ixp33_ASAP7_75t_SL g656 ( 
.A1(n_594),
.A2(n_481),
.B(n_406),
.C(n_459),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_599),
.Y(n_657)
);

BUFx4f_ASAP7_75t_SL g658 ( 
.A(n_602),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_521),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_534),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_606),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_534),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_550),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_577),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_547),
.B(n_480),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_549),
.B(n_401),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_606),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_577),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_529),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_578),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_547),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_578),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_578),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_606),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_489),
.B(n_392),
.Y(n_675)
);

OAI22xp33_ASAP7_75t_L g676 ( 
.A1(n_533),
.A2(n_451),
.B1(n_377),
.B2(n_454),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_585),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_521),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_496),
.B(n_482),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_550),
.Y(n_680)
);

AOI222xp33_ASAP7_75t_L g681 ( 
.A1(n_538),
.A2(n_482),
.B1(n_459),
.B2(n_461),
.C1(n_451),
.C2(n_377),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_500),
.A2(n_460),
.B(n_415),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_526),
.Y(n_683)
);

BUFx4_ASAP7_75t_SL g684 ( 
.A(n_496),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_491),
.A2(n_421),
.B1(n_487),
.B2(n_401),
.Y(n_685)
);

AOI221xp5_ASAP7_75t_L g686 ( 
.A1(n_525),
.A2(n_288),
.B1(n_311),
.B2(n_294),
.C(n_289),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_570),
.B(n_28),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_561),
.B(n_491),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_513),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_531),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_516),
.B(n_447),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_543),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_509),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_556),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_561),
.A2(n_447),
.B1(n_462),
.B2(n_457),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_535),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_579),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_566),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_599),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_491),
.A2(n_447),
.B1(n_462),
.B2(n_457),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_554),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_579),
.Y(n_702)
);

CKINVDCx11_ASAP7_75t_R g703 ( 
.A(n_496),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_524),
.B(n_511),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_535),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_527),
.A2(n_288),
.B(n_314),
.C(n_311),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_579),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_566),
.Y(n_708)
);

CKINVDCx6p67_ASAP7_75t_R g709 ( 
.A(n_572),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_591),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_500),
.A2(n_485),
.B(n_366),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_535),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_504),
.B(n_28),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_599),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_591),
.B(n_29),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_516),
.B(n_462),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_537),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_575),
.B(n_457),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_581),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_L g720 ( 
.A(n_507),
.B(n_288),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_581),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_576),
.B(n_580),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_618),
.A2(n_542),
.B(n_557),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_628),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_643),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_669),
.A2(n_538),
.B1(n_558),
.B2(n_565),
.Y(n_726)
);

INVxp33_ASAP7_75t_L g727 ( 
.A(n_665),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_654),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_650),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_622),
.B(n_693),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_655),
.A2(n_562),
.B1(n_560),
.B2(n_583),
.Y(n_731)
);

AND2x6_ASAP7_75t_SL g732 ( 
.A(n_679),
.B(n_594),
.Y(n_732)
);

AOI21x1_ASAP7_75t_L g733 ( 
.A1(n_618),
.A2(n_604),
.B(n_589),
.Y(n_733)
);

NAND2x1p5_ASAP7_75t_L g734 ( 
.A(n_611),
.B(n_553),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_619),
.Y(n_735)
);

AND2x2_ASAP7_75t_SL g736 ( 
.A(n_623),
.B(n_580),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_621),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_654),
.Y(n_738)
);

O2A1O1Ixp33_ASAP7_75t_SL g739 ( 
.A1(n_656),
.A2(n_583),
.B(n_560),
.C(n_567),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_690),
.Y(n_740)
);

BUFx2_ASAP7_75t_SL g741 ( 
.A(n_616),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_623),
.A2(n_548),
.B1(n_553),
.B2(n_564),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_692),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_611),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_689),
.B(n_572),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_675),
.B(n_653),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_622),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_613),
.B(n_598),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_635),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_704),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_679),
.A2(n_681),
.B1(n_676),
.B2(n_701),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_694),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_658),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_611),
.B(n_553),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_682),
.A2(n_653),
.B(n_639),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_715),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_679),
.A2(n_541),
.B1(n_497),
.B2(n_537),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_715),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_675),
.B(n_506),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_658),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_655),
.A2(n_677),
.B1(n_651),
.B2(n_627),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_661),
.Y(n_762)
);

BUFx8_ASAP7_75t_SL g763 ( 
.A(n_625),
.Y(n_763)
);

AOI221xp5_ASAP7_75t_L g764 ( 
.A1(n_676),
.A2(n_608),
.B1(n_595),
.B2(n_605),
.C(n_586),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_613),
.B(n_598),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_681),
.A2(n_713),
.B1(n_649),
.B2(n_630),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_633),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_649),
.A2(n_630),
.B1(n_688),
.B2(n_677),
.Y(n_768)
);

NOR2x1_ASAP7_75t_SL g769 ( 
.A(n_612),
.B(n_553),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_622),
.Y(n_770)
);

AOI221xp5_ASAP7_75t_L g771 ( 
.A1(n_627),
.A2(n_590),
.B1(n_596),
.B2(n_600),
.C(n_597),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_634),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_635),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_632),
.B(n_548),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_671),
.A2(n_562),
.B1(n_557),
.B2(n_541),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_636),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_646),
.A2(n_671),
.B1(n_703),
.B2(n_642),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_646),
.A2(n_497),
.B1(n_537),
.B2(n_546),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_659),
.A2(n_564),
.B1(n_587),
.B2(n_581),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_631),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_709),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_684),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_651),
.B(n_587),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_682),
.A2(n_542),
.B(n_584),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_640),
.B(n_587),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_710),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_710),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_640),
.A2(n_564),
.B1(n_518),
.B2(n_522),
.Y(n_788)
);

O2A1O1Ixp5_ASAP7_75t_L g789 ( 
.A1(n_687),
.A2(n_584),
.B(n_607),
.C(n_601),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_684),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_642),
.A2(n_545),
.B1(n_499),
.B2(n_571),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_678),
.B(n_563),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_SL g793 ( 
.A1(n_629),
.A2(n_564),
.B1(n_499),
.B2(n_571),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_609),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_698),
.A2(n_523),
.B1(n_522),
.B2(n_518),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_638),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_683),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_668),
.B(n_499),
.Y(n_798)
);

BUFx4_ASAP7_75t_R g799 ( 
.A(n_667),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_708),
.A2(n_551),
.B1(n_523),
.B2(n_563),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_SL g801 ( 
.A1(n_722),
.A2(n_571),
.B1(n_563),
.B2(n_493),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_609),
.B(n_495),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_661),
.B(n_551),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_660),
.A2(n_601),
.B1(n_501),
.B2(n_503),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_615),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_674),
.B(n_662),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_668),
.A2(n_510),
.B1(n_505),
.B2(n_508),
.Y(n_807)
);

AO31x2_ASAP7_75t_L g808 ( 
.A1(n_706),
.A2(n_510),
.A3(n_505),
.B(n_508),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_663),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_697),
.B(n_495),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_615),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_674),
.B(n_30),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_680),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_639),
.A2(n_507),
.B(n_559),
.Y(n_814)
);

AO31x2_ASAP7_75t_L g815 ( 
.A1(n_711),
.A2(n_552),
.A3(n_544),
.B(n_288),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_638),
.Y(n_816)
);

OR2x6_ASAP7_75t_L g817 ( 
.A(n_641),
.B(n_544),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_696),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_644),
.B(n_544),
.Y(n_819)
);

AO21x2_ASAP7_75t_L g820 ( 
.A1(n_711),
.A2(n_289),
.B(n_292),
.Y(n_820)
);

CKINVDCx12_ASAP7_75t_R g821 ( 
.A(n_610),
.Y(n_821)
);

AO31x2_ASAP7_75t_L g822 ( 
.A1(n_691),
.A2(n_716),
.A3(n_718),
.B(n_664),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_705),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_644),
.B(n_552),
.Y(n_824)
);

BUFx2_ASAP7_75t_SL g825 ( 
.A(n_644),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_712),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_617),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_697),
.B(n_31),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_719),
.A2(n_512),
.B1(n_559),
.B2(n_532),
.Y(n_829)
);

CKINVDCx11_ASAP7_75t_R g830 ( 
.A(n_614),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_615),
.Y(n_831)
);

CKINVDCx8_ASAP7_75t_R g832 ( 
.A(n_644),
.Y(n_832)
);

NAND2x1p5_ASAP7_75t_L g833 ( 
.A(n_614),
.B(n_552),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_719),
.A2(n_507),
.B1(n_559),
.B2(n_532),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_652),
.A2(n_670),
.B1(n_672),
.B2(n_673),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_717),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_718),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_702),
.A2(n_507),
.B1(n_559),
.B2(n_532),
.Y(n_838)
);

AOI221xp5_ASAP7_75t_L g839 ( 
.A1(n_691),
.A2(n_289),
.B1(n_292),
.B2(n_294),
.C(n_314),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_SL g840 ( 
.A1(n_707),
.A2(n_532),
.B1(n_512),
.B2(n_32),
.Y(n_840)
);

OAI21x1_ASAP7_75t_L g841 ( 
.A1(n_641),
.A2(n_573),
.B(n_512),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_614),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_700),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_626),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_647),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_721),
.A2(n_512),
.B1(n_289),
.B2(n_292),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_716),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_685),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_624),
.B(n_314),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_637),
.A2(n_289),
.B1(n_292),
.B2(n_294),
.Y(n_850)
);

AOI221xp5_ASAP7_75t_L g851 ( 
.A1(n_751),
.A2(n_686),
.B1(n_695),
.B2(n_720),
.C(n_666),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_746),
.A2(n_686),
.B1(n_699),
.B2(n_714),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_766),
.A2(n_714),
.B1(n_699),
.B2(n_657),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_735),
.B(n_714),
.Y(n_854)
);

NOR2x1_ASAP7_75t_L g855 ( 
.A(n_753),
.B(n_699),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_763),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_736),
.A2(n_657),
.B1(n_648),
.B2(n_645),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_737),
.B(n_724),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_755),
.A2(n_657),
.B(n_648),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_752),
.B(n_648),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_759),
.B(n_645),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_761),
.A2(n_645),
.B1(n_620),
.B2(n_292),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_730),
.B(n_620),
.Y(n_863)
);

BUFx12f_ASAP7_75t_L g864 ( 
.A(n_790),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_750),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_SL g866 ( 
.A1(n_770),
.A2(n_620),
.B1(n_294),
.B2(n_314),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_759),
.A2(n_420),
.B(n_449),
.C(n_432),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_725),
.B(n_34),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_777),
.A2(n_485),
.B1(n_449),
.B2(n_432),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_726),
.A2(n_843),
.B1(n_761),
.B2(n_745),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_SL g871 ( 
.A1(n_770),
.A2(n_485),
.B1(n_449),
.B2(n_432),
.Y(n_871)
);

BUFx12f_ASAP7_75t_L g872 ( 
.A(n_772),
.Y(n_872)
);

OAI211xp5_ASAP7_75t_SL g873 ( 
.A1(n_794),
.A2(n_36),
.B(n_43),
.C(n_46),
.Y(n_873)
);

AOI21xp33_ASAP7_75t_L g874 ( 
.A1(n_795),
.A2(n_431),
.B(n_430),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_SL g875 ( 
.A1(n_782),
.A2(n_431),
.B1(n_430),
.B2(n_420),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_745),
.B(n_49),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_783),
.A2(n_431),
.B1(n_430),
.B2(n_420),
.Y(n_877)
);

OAI221xp5_ASAP7_75t_L g878 ( 
.A1(n_768),
.A2(n_412),
.B1(n_409),
.B2(n_375),
.C(n_373),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_780),
.B(n_50),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_785),
.A2(n_412),
.B1(n_409),
.B2(n_375),
.Y(n_880)
);

OAI21x1_ASAP7_75t_L g881 ( 
.A1(n_733),
.A2(n_409),
.B(n_375),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_739),
.A2(n_412),
.B(n_373),
.Y(n_882)
);

OAI22xp33_ASAP7_75t_L g883 ( 
.A1(n_727),
.A2(n_373),
.B1(n_366),
.B2(n_55),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_814),
.A2(n_366),
.B(n_53),
.Y(n_884)
);

OAI21xp33_ASAP7_75t_L g885 ( 
.A1(n_764),
.A2(n_51),
.B(n_60),
.Y(n_885)
);

AOI211xp5_ASAP7_75t_L g886 ( 
.A1(n_792),
.A2(n_68),
.B(n_75),
.C(n_77),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_830),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_847),
.A2(n_848),
.B1(n_837),
.B2(n_728),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_740),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_738),
.A2(n_80),
.B1(n_83),
.B2(n_87),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_757),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_743),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_785),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_756),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_758),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_786),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_771),
.A2(n_119),
.B1(n_122),
.B2(n_126),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_787),
.B(n_147),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_817),
.B(n_127),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_729),
.A2(n_128),
.B1(n_135),
.B2(n_138),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_767),
.B(n_140),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_799),
.Y(n_902)
);

AOI21xp33_ASAP7_75t_L g903 ( 
.A1(n_795),
.A2(n_146),
.B(n_143),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_809),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_747),
.B(n_144),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_812),
.A2(n_828),
.B1(n_800),
.B2(n_731),
.Y(n_906)
);

AOI221xp5_ASAP7_75t_L g907 ( 
.A1(n_731),
.A2(n_776),
.B1(n_813),
.B2(n_791),
.C(n_800),
.Y(n_907)
);

INVx4_ASAP7_75t_L g908 ( 
.A(n_781),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_741),
.B(n_760),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_805),
.B(n_802),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_788),
.A2(n_807),
.B1(n_840),
.B2(n_801),
.Y(n_911)
);

OAI221xp5_ASAP7_75t_L g912 ( 
.A1(n_778),
.A2(n_775),
.B1(n_804),
.B2(n_789),
.C(n_788),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_802),
.B(n_774),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_806),
.A2(n_762),
.B1(n_765),
.B2(n_748),
.Y(n_914)
);

NAND3xp33_ASAP7_75t_L g915 ( 
.A(n_839),
.B(n_784),
.C(n_850),
.Y(n_915)
);

OAI221xp5_ASAP7_75t_L g916 ( 
.A1(n_793),
.A2(n_823),
.B1(n_818),
.B2(n_826),
.C(n_836),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_797),
.A2(n_821),
.B1(n_807),
.B2(n_765),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_832),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_845),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_835),
.A2(n_817),
.B1(n_762),
.B2(n_779),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_835),
.A2(n_817),
.B1(n_811),
.B2(n_810),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_827),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_811),
.A2(n_810),
.B1(n_838),
.B2(n_825),
.Y(n_923)
);

INVxp67_ASAP7_75t_SL g924 ( 
.A(n_769),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_774),
.B(n_744),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_803),
.Y(n_926)
);

NAND2x1_ASAP7_75t_L g927 ( 
.A(n_819),
.B(n_824),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_SL g928 ( 
.A1(n_732),
.A2(n_748),
.B1(n_834),
.B2(n_838),
.Y(n_928)
);

OAI211xp5_ASAP7_75t_L g929 ( 
.A1(n_831),
.A2(n_816),
.B(n_749),
.C(n_796),
.Y(n_929)
);

OAI221xp5_ASAP7_75t_SL g930 ( 
.A1(n_723),
.A2(n_798),
.B1(n_773),
.B2(n_844),
.C(n_849),
.Y(n_930)
);

OAI22xp33_ASAP7_75t_L g931 ( 
.A1(n_798),
.A2(n_744),
.B1(n_834),
.B2(n_742),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_822),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_819),
.A2(n_824),
.B1(n_754),
.B2(n_829),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_822),
.B(n_734),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_822),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_808),
.Y(n_936)
);

AO221x1_ASAP7_75t_L g937 ( 
.A1(n_846),
.A2(n_842),
.B1(n_833),
.B2(n_815),
.C(n_734),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_808),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_808),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_833),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_861),
.Y(n_941)
);

AOI33xp33_ASAP7_75t_L g942 ( 
.A1(n_865),
.A2(n_892),
.A3(n_888),
.B1(n_928),
.B2(n_858),
.B3(n_870),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_889),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_L g944 ( 
.A(n_886),
.B(n_846),
.C(n_842),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_911),
.A2(n_820),
.B1(n_842),
.B2(n_841),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_911),
.A2(n_815),
.B1(n_820),
.B2(n_902),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_926),
.B(n_815),
.Y(n_947)
);

OAI221xp5_ASAP7_75t_L g948 ( 
.A1(n_906),
.A2(n_917),
.B1(n_914),
.B2(n_907),
.C(n_912),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_902),
.A2(n_916),
.B1(n_921),
.B2(n_899),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_896),
.B(n_904),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_861),
.Y(n_951)
);

OAI221xp5_ASAP7_75t_L g952 ( 
.A1(n_933),
.A2(n_851),
.B1(n_913),
.B2(n_885),
.C(n_868),
.Y(n_952)
);

OAI222xp33_ASAP7_75t_L g953 ( 
.A1(n_921),
.A2(n_920),
.B1(n_923),
.B2(n_899),
.C1(n_893),
.C2(n_934),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_932),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_919),
.Y(n_955)
);

OAI221xp5_ASAP7_75t_L g956 ( 
.A1(n_853),
.A2(n_930),
.B1(n_910),
.B2(n_869),
.C(n_920),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_876),
.A2(n_924),
.B1(n_879),
.B2(n_909),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_918),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_935),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_881),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_922),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_908),
.B(n_918),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_876),
.A2(n_923),
.B1(n_852),
.B2(n_931),
.Y(n_963)
);

AOI221xp5_ASAP7_75t_SL g964 ( 
.A1(n_893),
.A2(n_905),
.B1(n_898),
.B2(n_901),
.C(n_863),
.Y(n_964)
);

OA21x2_ASAP7_75t_L g965 ( 
.A1(n_936),
.A2(n_938),
.B(n_939),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_860),
.A2(n_937),
.B1(n_918),
.B2(n_903),
.Y(n_966)
);

AOI221xp5_ASAP7_75t_L g967 ( 
.A1(n_903),
.A2(n_908),
.B1(n_874),
.B2(n_887),
.C(n_873),
.Y(n_967)
);

INVxp67_ASAP7_75t_SL g968 ( 
.A(n_854),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_862),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_855),
.Y(n_970)
);

AOI221xp5_ASAP7_75t_L g971 ( 
.A1(n_874),
.A2(n_887),
.B1(n_862),
.B2(n_929),
.C(n_915),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_927),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_940),
.Y(n_973)
);

NAND3xp33_ASAP7_75t_L g974 ( 
.A(n_897),
.B(n_900),
.C(n_890),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_877),
.A2(n_880),
.B(n_867),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_925),
.B(n_940),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_880),
.Y(n_977)
);

OAI222xp33_ASAP7_75t_L g978 ( 
.A1(n_856),
.A2(n_925),
.B1(n_866),
.B2(n_878),
.C1(n_891),
.C2(n_877),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_925),
.A2(n_887),
.B1(n_883),
.B2(n_857),
.Y(n_979)
);

OAI33xp33_ASAP7_75t_L g980 ( 
.A1(n_864),
.A2(n_872),
.A3(n_895),
.B1(n_894),
.B2(n_884),
.B3(n_875),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_859),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_882),
.B(n_871),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_926),
.B(n_751),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_858),
.B(n_889),
.Y(n_984)
);

NAND3xp33_ASAP7_75t_L g985 ( 
.A(n_928),
.B(n_533),
.C(n_467),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_858),
.B(n_889),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_928),
.A2(n_679),
.B1(n_751),
.B2(n_681),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_858),
.B(n_889),
.Y(n_988)
);

OAI221xp5_ASAP7_75t_L g989 ( 
.A1(n_870),
.A2(n_751),
.B1(n_679),
.B2(n_746),
.C(n_777),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_932),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_906),
.A2(n_483),
.B1(n_751),
.B2(n_623),
.Y(n_991)
);

OA21x2_ASAP7_75t_L g992 ( 
.A1(n_936),
.A2(n_938),
.B(n_939),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_954),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_954),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_990),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_941),
.B(n_951),
.Y(n_996)
);

AOI221xp5_ASAP7_75t_L g997 ( 
.A1(n_991),
.A2(n_987),
.B1(n_948),
.B2(n_989),
.C(n_953),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_947),
.Y(n_998)
);

NAND2x1_ASAP7_75t_L g999 ( 
.A(n_959),
.B(n_990),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_972),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_984),
.B(n_988),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_965),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_984),
.B(n_988),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_986),
.B(n_962),
.Y(n_1004)
);

AOI211x1_ASAP7_75t_L g1005 ( 
.A1(n_985),
.A2(n_952),
.B(n_956),
.C(n_986),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_992),
.B(n_965),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_955),
.B(n_943),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_981),
.B(n_977),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_983),
.B(n_968),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_942),
.B(n_983),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_992),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_961),
.B(n_946),
.Y(n_1012)
);

OAI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_957),
.A2(n_963),
.B1(n_950),
.B2(n_976),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_969),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_977),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_976),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_969),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_949),
.B(n_945),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_942),
.B(n_964),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_973),
.B(n_981),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1001),
.B(n_966),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1001),
.B(n_960),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_1002),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1003),
.B(n_960),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_998),
.B(n_958),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1003),
.B(n_960),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_1008),
.B(n_960),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_1014),
.B(n_971),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_1006),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_993),
.B(n_970),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_997),
.A2(n_980),
.B1(n_967),
.B2(n_974),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_998),
.B(n_979),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_993),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_1009),
.B(n_975),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1030),
.B(n_1007),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1023),
.Y(n_1036)
);

OAI221xp5_ASAP7_75t_L g1037 ( 
.A1(n_1031),
.A2(n_997),
.B1(n_1019),
.B2(n_1010),
.C(n_1004),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1030),
.B(n_1007),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1022),
.B(n_1006),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1033),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1022),
.B(n_1006),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1024),
.B(n_1014),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_1021),
.B(n_1010),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1024),
.B(n_1026),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1026),
.B(n_1008),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1021),
.B(n_1012),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1033),
.B(n_1012),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1043),
.B(n_1029),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_1044),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1046),
.B(n_1029),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1042),
.B(n_1029),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_1036),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1040),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1042),
.B(n_1034),
.Y(n_1054)
);

NOR2x1_ASAP7_75t_L g1055 ( 
.A(n_1037),
.B(n_1000),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1035),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1036),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1038),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_1054),
.B(n_1039),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_1049),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1053),
.Y(n_1061)
);

XOR2x2_ASAP7_75t_L g1062 ( 
.A(n_1055),
.B(n_1005),
.Y(n_1062)
);

AOI211xp5_ASAP7_75t_L g1063 ( 
.A1(n_1048),
.A2(n_1013),
.B(n_1034),
.C(n_1019),
.Y(n_1063)
);

OAI211xp5_ASAP7_75t_L g1064 ( 
.A1(n_1056),
.A2(n_1031),
.B(n_1005),
.C(n_1058),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_1050),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1051),
.Y(n_1066)
);

NAND3xp33_ASAP7_75t_L g1067 ( 
.A(n_1052),
.B(n_1028),
.C(n_1025),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1052),
.B(n_1039),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_SL g1069 ( 
.A1(n_1057),
.A2(n_1032),
.B1(n_1025),
.B2(n_1000),
.Y(n_1069)
);

OAI221xp5_ASAP7_75t_L g1070 ( 
.A1(n_1062),
.A2(n_1032),
.B1(n_1047),
.B2(n_1028),
.C(n_1009),
.Y(n_1070)
);

NOR3x1_ASAP7_75t_L g1071 ( 
.A(n_1064),
.B(n_1015),
.C(n_1013),
.Y(n_1071)
);

OAI21xp33_ASAP7_75t_L g1072 ( 
.A1(n_1062),
.A2(n_1018),
.B(n_1044),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1061),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1068),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_1060),
.B(n_1045),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_1065),
.Y(n_1076)
);

XNOR2xp5_ASAP7_75t_L g1077 ( 
.A(n_1065),
.B(n_1041),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1072),
.A2(n_1063),
.B1(n_1069),
.B2(n_1067),
.Y(n_1078)
);

AOI221xp5_ASAP7_75t_L g1079 ( 
.A1(n_1072),
.A2(n_1066),
.B1(n_1068),
.B2(n_1059),
.C(n_1041),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1073),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_1076),
.B(n_1057),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1077),
.A2(n_978),
.B(n_1018),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_SL g1083 ( 
.A(n_1071),
.B(n_944),
.C(n_1015),
.Y(n_1083)
);

NOR3xp33_ASAP7_75t_L g1084 ( 
.A(n_1083),
.B(n_1070),
.C(n_1074),
.Y(n_1084)
);

NAND3xp33_ASAP7_75t_SL g1085 ( 
.A(n_1078),
.B(n_999),
.C(n_1045),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1080),
.Y(n_1086)
);

AOI22x1_ASAP7_75t_L g1087 ( 
.A1(n_1082),
.A2(n_1075),
.B1(n_982),
.B2(n_1020),
.Y(n_1087)
);

NOR4xp25_ASAP7_75t_L g1088 ( 
.A(n_1079),
.B(n_994),
.C(n_995),
.D(n_1020),
.Y(n_1088)
);

OR4x2_ASAP7_75t_L g1089 ( 
.A(n_1085),
.B(n_1081),
.C(n_1075),
.D(n_1016),
.Y(n_1089)
);

OAI211xp5_ASAP7_75t_L g1090 ( 
.A1(n_1087),
.A2(n_1000),
.B(n_994),
.C(n_995),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1086),
.Y(n_1091)
);

OR3x2_ASAP7_75t_L g1092 ( 
.A(n_1084),
.B(n_1088),
.C(n_1011),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_1086),
.Y(n_1093)
);

XNOR2xp5_ASAP7_75t_L g1094 ( 
.A(n_1091),
.B(n_1090),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1093),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1092),
.A2(n_1016),
.B1(n_1027),
.B2(n_996),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_1093),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_SL g1098 ( 
.A1(n_1097),
.A2(n_1089),
.B1(n_982),
.B2(n_1016),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_1098),
.Y(n_1099)
);

AOI22x1_ASAP7_75t_L g1100 ( 
.A1(n_1099),
.A2(n_1095),
.B1(n_1094),
.B2(n_1096),
.Y(n_1100)
);

AOI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_1100),
.A2(n_999),
.B(n_1017),
.Y(n_1101)
);


endmodule