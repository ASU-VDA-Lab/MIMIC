module fake_jpeg_21277_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_8),
.C(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_47),
.B(n_54),
.Y(n_112)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_50),
.B(n_59),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_19),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_55),
.Y(n_72)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_0),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_33),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_20),
.B(n_9),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_66),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_32),
.B1(n_23),
.B2(n_17),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_68),
.A2(n_102),
.B1(n_105),
.B2(n_109),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_80),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_34),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_78),
.B(n_79),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_34),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_53),
.B(n_32),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_83),
.B(n_29),
.C(n_31),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_84),
.B(n_92),
.Y(n_153)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_55),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_29),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_23),
.B1(n_17),
.B2(n_24),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_41),
.B1(n_44),
.B2(n_27),
.Y(n_127)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_94),
.Y(n_132)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_20),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_63),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_101),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_23),
.B1(n_17),
.B2(n_30),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_111),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_57),
.A2(n_35),
.B1(n_40),
.B2(n_26),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_45),
.B(n_26),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_57),
.A2(n_35),
.B1(n_40),
.B2(n_38),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_37),
.B1(n_22),
.B2(n_24),
.Y(n_151)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_29),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_62),
.B1(n_43),
.B2(n_46),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_118),
.A2(n_138),
.B1(n_151),
.B2(n_152),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

NAND2x1_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_49),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_SL g157 ( 
.A(n_122),
.B(n_68),
.C(n_102),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_127),
.A2(n_154),
.B1(n_82),
.B2(n_107),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_74),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_18),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_133),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_28),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_28),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_150),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_76),
.B(n_117),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_31),
.B1(n_24),
.B2(n_36),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_93),
.A2(n_36),
.B1(n_37),
.B2(n_22),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_29),
.B(n_28),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_0),
.B(n_1),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_99),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_130),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_70),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_105),
.A2(n_31),
.B1(n_24),
.B2(n_22),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_113),
.A2(n_31),
.B1(n_37),
.B2(n_2),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_157),
.A2(n_161),
.B(n_162),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_107),
.B1(n_97),
.B2(n_88),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_122),
.A2(n_76),
.B(n_100),
.C(n_69),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_96),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_138),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_167),
.A2(n_177),
.B(n_178),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_96),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_181),
.Y(n_209)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_97),
.B1(n_104),
.B2(n_108),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_153),
.B(n_14),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_174),
.B(n_175),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_153),
.B(n_12),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_132),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_176),
.B(n_184),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_104),
.B(n_77),
.C(n_82),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_71),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_118),
.A2(n_77),
.B1(n_81),
.B2(n_71),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_134),
.B(n_10),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_134),
.B(n_136),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_187),
.Y(n_201)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_128),
.B(n_116),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_116),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_191),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_146),
.A2(n_81),
.B1(n_2),
.B2(n_3),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_189),
.A2(n_149),
.B1(n_131),
.B2(n_142),
.Y(n_204)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_129),
.B(n_10),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_73),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_120),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_122),
.C(n_144),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_199),
.C(n_207),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_160),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_213),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_131),
.Y(n_200)
);

AOI221xp5_ASAP7_75t_L g247 ( 
.A1(n_200),
.A2(n_189),
.B1(n_184),
.B2(n_191),
.C(n_174),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_204),
.A2(n_205),
.B1(n_211),
.B2(n_183),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_182),
.A2(n_126),
.B1(n_145),
.B2(n_141),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_148),
.C(n_126),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_148),
.C(n_123),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_210),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_123),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_182),
.A2(n_121),
.B1(n_125),
.B2(n_119),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_1),
.B(n_3),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_164),
.B(n_161),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_215),
.B(n_219),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_125),
.C(n_119),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_218),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_162),
.B(n_120),
.C(n_73),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_162),
.B(n_120),
.C(n_7),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_1),
.Y(n_220)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_162),
.B(n_7),
.C(n_11),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_219),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_171),
.Y(n_223)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_156),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_228),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_15),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_227),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_229),
.B(n_232),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_201),
.B(n_175),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_236),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_200),
.A2(n_177),
.B1(n_157),
.B2(n_158),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_238),
.B1(n_245),
.B2(n_253),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_222),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_246),
.B(n_248),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_210),
.A2(n_159),
.B1(n_164),
.B2(n_171),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_249),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_209),
.B1(n_215),
.B2(n_202),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_197),
.A2(n_172),
.B1(n_192),
.B2(n_173),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_217),
.A2(n_192),
.B(n_186),
.Y(n_246)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_202),
.C(n_220),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_217),
.A2(n_173),
.B(n_190),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_197),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_252),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_226),
.A2(n_169),
.B(n_165),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_251),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_226),
.A2(n_169),
.B(n_165),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_223),
.A2(n_180),
.B1(n_194),
.B2(n_156),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_261),
.A2(n_274),
.B(n_248),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_244),
.A2(n_207),
.B1(n_208),
.B2(n_216),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_270),
.B1(n_238),
.B2(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_195),
.C(n_199),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_267),
.C(n_240),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_209),
.C(n_218),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_231),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_249),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_212),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_272),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_231),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_230),
.B(n_254),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_275),
.Y(n_288)
);

AOI32xp33_ASAP7_75t_L g274 ( 
.A1(n_237),
.A2(n_203),
.A3(n_214),
.B1(n_196),
.B2(n_228),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_229),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_246),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_284),
.Y(n_294)
);

AOI21x1_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_248),
.B(n_252),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_SL g297 ( 
.A(n_281),
.B(n_256),
.Y(n_297)
);

BUFx12f_ASAP7_75t_SL g282 ( 
.A(n_274),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_285),
.B(n_290),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_240),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_259),
.C(n_276),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_235),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_292),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_260),
.A2(n_268),
.B(n_264),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_258),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_259),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_283),
.B(n_232),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_301),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_290),
.B(n_256),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_303),
.C(n_306),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_257),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_278),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_242),
.C(n_257),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_272),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_305),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_258),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_242),
.C(n_273),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_282),
.B(n_269),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_315),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_292),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_285),
.C(n_291),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_281),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_316),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_311),
.A2(n_297),
.B(n_288),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_302),
.A3(n_265),
.B1(n_306),
.B2(n_241),
.C1(n_294),
.C2(n_233),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_307),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_241),
.B(n_294),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_243),
.B(n_224),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_323),
.A2(n_243),
.B(n_307),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_315),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_324),
.B(n_326),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_314),
.B1(n_322),
.B2(n_321),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_327),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_317),
.A2(n_310),
.B(n_221),
.C(n_227),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_329),
.A2(n_328),
.B1(n_4),
.B2(n_5),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_331),
.Y(n_332)
);

MAJx2_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_330),
.C(n_331),
.Y(n_333)
);


endmodule