module fake_ibex_1328_n_4110 (n_151, n_85, n_599, n_778, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_738, n_475, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_785, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_768, n_338, n_173, n_696, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_592, n_495, n_762, n_410, n_308, n_675, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_217, n_324, n_391, n_537, n_728, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_232, n_380, n_749, n_281, n_559, n_425, n_4110);

input n_151;
input n_85;
input n_599;
input n_778;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_738;
input n_475;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_785;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_768;
input n_338;
input n_173;
input n_696;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4110;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_2607;
wire n_1382;
wire n_3548;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_845;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_802;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3440;
wire n_3135;
wire n_3904;
wire n_850;
wire n_3729;
wire n_3175;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_3984;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_1766;
wire n_3566;
wire n_3184;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_824;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3884;
wire n_3949;
wire n_3507;
wire n_3881;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2846;
wire n_2685;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2413;
wire n_2249;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_3973;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_3097;
wire n_2906;
wire n_3030;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2806;
wire n_2283;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_1637;
wire n_3858;
wire n_841;
wire n_2900;
wire n_3310;
wire n_810;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_1620;
wire n_869;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3874;
wire n_1281;
wire n_3094;
wire n_3217;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_4079;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4103;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_819;
wire n_3950;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3733;
wire n_3626;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2573;
wire n_2423;
wire n_859;
wire n_3849;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4092;
wire n_3003;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_3331;
wire n_2910;
wire n_3119;
wire n_2590;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2991;
wire n_2234;
wire n_847;
wire n_2699;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3797;
wire n_3441;
wire n_1395;
wire n_998;
wire n_1729;
wire n_1115;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_4047;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_814;
wire n_3829;
wire n_1864;
wire n_943;
wire n_3087;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_803;
wire n_2570;
wire n_4051;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3719;
wire n_3390;
wire n_3948;
wire n_1400;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_3070;
wire n_3477;
wire n_3646;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_1439;
wire n_2263;
wire n_2352;
wire n_2212;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2654;
wire n_2463;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_1185;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2875;
wire n_2684;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_991;
wire n_1331;
wire n_961;
wire n_1223;
wire n_2127;
wire n_3747;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_4071;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3673;
wire n_3476;
wire n_2842;
wire n_3990;
wire n_2994;
wire n_2011;
wire n_4066;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_4085;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_798;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_838;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4099;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_3930;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2320;
wire n_2237;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_4022;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_3162;
wire n_2984;
wire n_2732;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_3044;
wire n_3493;
wire n_2447;
wire n_2868;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3538;
wire n_1261;
wire n_2299;
wire n_3393;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3647;
wire n_3623;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3604;
wire n_1838;
wire n_3649;
wire n_833;
wire n_3540;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_3059;
wire n_2567;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_4058;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_4017;
wire n_1547;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1542;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_956;
wire n_3561;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3942;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_3102;
wire n_2872;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4049;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3343;
wire n_3163;
wire n_3752;
wire n_3786;
wire n_4061;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_4045;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1992;
wire n_1685;
wire n_1784;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1488;
wire n_849;
wire n_1193;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3380;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_4038;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1516;
wire n_1027;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2303;
wire n_949;
wire n_2357;
wire n_2104;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_3938;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_4088;
wire n_2136;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_2802;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3689;
wire n_3582;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_3527;
wire n_2754;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_799;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2917;
wire n_2726;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4106;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_4075;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2349;
wire n_2100;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

INVx1_ASAP7_75t_L g793 ( 
.A(n_658),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_633),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_714),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_704),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_766),
.Y(n_797)
);

CKINVDCx16_ASAP7_75t_R g798 ( 
.A(n_507),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_93),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_692),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_767),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_513),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_442),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_490),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_281),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_284),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_468),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_436),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_75),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_66),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_579),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_476),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_230),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_92),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_357),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_440),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_296),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_557),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_746),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_760),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_342),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_282),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_347),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_210),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_779),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_747),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_256),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_594),
.Y(n_828)
);

CKINVDCx14_ASAP7_75t_R g829 ( 
.A(n_290),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_109),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_757),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_532),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_334),
.B(n_584),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_240),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_792),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_368),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_632),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_64),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_578),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_398),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_465),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_706),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_692),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_589),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_417),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_41),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_305),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_153),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_159),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_154),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_256),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_375),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_680),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_102),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_787),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_693),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_584),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_143),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_435),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_216),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_650),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_652),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_95),
.B(n_449),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_275),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_130),
.Y(n_865)
);

BUFx10_ASAP7_75t_L g866 ( 
.A(n_639),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_29),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_699),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_3),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_667),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_480),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_144),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_289),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_24),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_206),
.Y(n_875)
);

BUFx10_ASAP7_75t_L g876 ( 
.A(n_7),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_254),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_645),
.B(n_356),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_594),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_492),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_152),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_349),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_522),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_764),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_619),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_643),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_68),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_11),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_312),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_43),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_211),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_151),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_72),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_667),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_40),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_L g896 ( 
.A(n_270),
.B(n_315),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_213),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_506),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_47),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_547),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_63),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_618),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_547),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_533),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_554),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_527),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_622),
.Y(n_907)
);

CKINVDCx20_ASAP7_75t_R g908 ( 
.A(n_645),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_287),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_23),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_414),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_739),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_127),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_373),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_722),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_631),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_710),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_636),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_320),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_600),
.Y(n_920)
);

CKINVDCx16_ASAP7_75t_R g921 ( 
.A(n_769),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_238),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_770),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_400),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_247),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_790),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_499),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_65),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_608),
.Y(n_929)
);

BUFx5_ASAP7_75t_L g930 ( 
.A(n_751),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_637),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_251),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_221),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_307),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_397),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_106),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_225),
.Y(n_937)
);

CKINVDCx16_ASAP7_75t_R g938 ( 
.A(n_124),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_774),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_250),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_633),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_445),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_9),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_604),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_519),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_96),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_660),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_555),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_175),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_118),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_738),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_158),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_112),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_340),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_452),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_146),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_227),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_186),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_244),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_697),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_78),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_590),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_368),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_521),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_367),
.B(n_234),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_517),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_715),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_249),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_407),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_236),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_239),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_359),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_775),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_118),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_354),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_456),
.B(n_107),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_516),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_4),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_647),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_336),
.B(n_250),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_321),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_506),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_309),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_791),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_622),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_579),
.Y(n_986)
);

BUFx10_ASAP7_75t_L g987 ( 
.A(n_311),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_301),
.Y(n_988)
);

BUFx10_ASAP7_75t_L g989 ( 
.A(n_778),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_329),
.Y(n_990)
);

BUFx5_ASAP7_75t_L g991 ( 
.A(n_394),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_9),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_718),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_317),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_16),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_285),
.Y(n_996)
);

INVxp67_ASAP7_75t_SL g997 ( 
.A(n_785),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_468),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_524),
.Y(n_999)
);

CKINVDCx16_ASAP7_75t_R g1000 ( 
.A(n_739),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_736),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_451),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_117),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_77),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_689),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_641),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_213),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_32),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_13),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_488),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_306),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_326),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_401),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_76),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_711),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_345),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_260),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_761),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_128),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_285),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_738),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_581),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_95),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_651),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_414),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_220),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_187),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_92),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_449),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_725),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_98),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_286),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_157),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_271),
.Y(n_1034)
);

BUFx5_ASAP7_75t_L g1035 ( 
.A(n_789),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_600),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_280),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_87),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_140),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_93),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_505),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_525),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_272),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_77),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_72),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_715),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_527),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_76),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_245),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_362),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_313),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_263),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_55),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_765),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_324),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_181),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_424),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_230),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_90),
.Y(n_1059)
);

BUFx5_ASAP7_75t_L g1060 ( 
.A(n_23),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_25),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_67),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_154),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_542),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_514),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_123),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_189),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_374),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_534),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_613),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_610),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_514),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_593),
.Y(n_1073)
);

CKINVDCx16_ASAP7_75t_R g1074 ( 
.A(n_100),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_536),
.Y(n_1075)
);

BUFx10_ASAP7_75t_L g1076 ( 
.A(n_642),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_172),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_648),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_582),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_403),
.Y(n_1080)
);

NOR2xp67_ASAP7_75t_L g1081 ( 
.A(n_513),
.B(n_710),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_587),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_477),
.Y(n_1083)
);

CKINVDCx14_ASAP7_75t_R g1084 ( 
.A(n_385),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_783),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_48),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_238),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_244),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_782),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_322),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_721),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_114),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_304),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_84),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_366),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_669),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_502),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_529),
.Y(n_1098)
);

CKINVDCx16_ASAP7_75t_R g1099 ( 
.A(n_161),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_730),
.Y(n_1100)
);

CKINVDCx16_ASAP7_75t_R g1101 ( 
.A(n_722),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_695),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_407),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_585),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_8),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_478),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_697),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_362),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_355),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_538),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_198),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_777),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_712),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_538),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_330),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_691),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_192),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_303),
.Y(n_1118)
);

CKINVDCx14_ASAP7_75t_R g1119 ( 
.A(n_371),
.Y(n_1119)
);

BUFx8_ASAP7_75t_SL g1120 ( 
.A(n_726),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_683),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_15),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_619),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_444),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_106),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_446),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_781),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_483),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_224),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_466),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_618),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_609),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_237),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_254),
.B(n_426),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_65),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_713),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_99),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_263),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_204),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_482),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_345),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_654),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_411),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_158),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_473),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_708),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_719),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_7),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_545),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_435),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_287),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_723),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_295),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_400),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_139),
.Y(n_1155)
);

CKINVDCx14_ASAP7_75t_R g1156 ( 
.A(n_84),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_459),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_674),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_536),
.Y(n_1159)
);

BUFx8_ASAP7_75t_SL g1160 ( 
.A(n_203),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_378),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_720),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_744),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_301),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_716),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_436),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_36),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_24),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_17),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_433),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_204),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_571),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_705),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_626),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_729),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_261),
.Y(n_1176)
);

INVxp33_ASAP7_75t_L g1177 ( 
.A(n_310),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_773),
.Y(n_1178)
);

INVxp67_ASAP7_75t_SL g1179 ( 
.A(n_398),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_788),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_717),
.Y(n_1181)
);

BUFx10_ASAP7_75t_L g1182 ( 
.A(n_728),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_81),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_86),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_726),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_293),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_511),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_119),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_235),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_296),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_232),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_258),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_709),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_528),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_111),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_580),
.Y(n_1196)
);

BUFx5_ASAP7_75t_L g1197 ( 
.A(n_580),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_554),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_479),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_239),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_179),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_412),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_385),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_763),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_640),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_218),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_40),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_286),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_505),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_366),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_211),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_137),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_569),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_664),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_78),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_470),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_724),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_161),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_674),
.Y(n_1219)
);

BUFx10_ASAP7_75t_L g1220 ( 
.A(n_156),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_754),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_752),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_393),
.Y(n_1223)
);

BUFx5_ASAP7_75t_L g1224 ( 
.A(n_228),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_707),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_604),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_934),
.B(n_0),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_829),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_991),
.Y(n_1229)
);

BUFx8_ASAP7_75t_SL g1230 ( 
.A(n_1120),
.Y(n_1230)
);

INVx6_ASAP7_75t_L g1231 ( 
.A(n_989),
.Y(n_1231)
);

BUFx8_ASAP7_75t_SL g1232 ( 
.A(n_1120),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_934),
.B(n_1),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_807),
.B(n_3),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1177),
.B(n_2),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_991),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_991),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_919),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_991),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_991),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_991),
.Y(n_1241)
);

OAI22x1_ASAP7_75t_R g1242 ( 
.A1(n_815),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_919),
.Y(n_1243)
);

BUFx12f_ASAP7_75t_L g1244 ( 
.A(n_866),
.Y(n_1244)
);

INVx5_ASAP7_75t_L g1245 ( 
.A(n_989),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_814),
.B(n_6),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_991),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1060),
.Y(n_1248)
);

BUFx8_ASAP7_75t_SL g1249 ( 
.A(n_1160),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1060),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_919),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_943),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_943),
.B(n_5),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1060),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_819),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1018),
.B(n_8),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1060),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_847),
.B(n_978),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1060),
.Y(n_1259)
);

OA21x2_ASAP7_75t_L g1260 ( 
.A1(n_855),
.A2(n_749),
.B(n_748),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1060),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_866),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1060),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1197),
.Y(n_1264)
);

INVx5_ASAP7_75t_L g1265 ( 
.A(n_989),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1197),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1197),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_840),
.B(n_11),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_803),
.B(n_10),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_919),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1197),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_829),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1197),
.Y(n_1273)
);

BUFx8_ASAP7_75t_L g1274 ( 
.A(n_971),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1177),
.B(n_10),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1033),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1084),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_803),
.B(n_12),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1033),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1084),
.B(n_12),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1197),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1224),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_866),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_824),
.B(n_13),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_859),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1224),
.Y(n_1286)
);

INVx6_ASAP7_75t_L g1287 ( 
.A(n_876),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_825),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_855),
.A2(n_753),
.B(n_750),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_831),
.A2(n_756),
.B(n_755),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_835),
.B(n_14),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1033),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1119),
.B(n_14),
.Y(n_1293)
);

OAI22x1_ASAP7_75t_SL g1294 ( 
.A1(n_815),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1294)
);

BUFx8_ASAP7_75t_L g1295 ( 
.A(n_1224),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_797),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1033),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_926),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1224),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1047),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1047),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1047),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1047),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1119),
.A2(n_1156),
.B1(n_938),
.B2(n_1000),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1156),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1305)
);

INVxp33_ASAP7_75t_SL g1306 ( 
.A(n_861),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_876),
.Y(n_1307)
);

INVx5_ASAP7_75t_L g1308 ( 
.A(n_1067),
.Y(n_1308)
);

INVx5_ASAP7_75t_L g1309 ( 
.A(n_1067),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_824),
.B(n_19),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_876),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1224),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1224),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1067),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1224),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_798),
.B(n_20),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_895),
.B(n_21),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1067),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_895),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1074),
.B(n_1099),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1204),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1093),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_973),
.A2(n_759),
.B(n_758),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1093),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_830),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1190),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_830),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_916),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1306),
.A2(n_1285),
.B1(n_1304),
.B2(n_1320),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1319),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1227),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1230),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1232),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1272),
.B(n_1101),
.Y(n_1334)
);

BUFx4f_ASAP7_75t_L g1335 ( 
.A(n_1244),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1249),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1277),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1227),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1288),
.Y(n_1339)
);

AOI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1236),
.A2(n_1112),
.B(n_1089),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1304),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1298),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1283),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1311),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1274),
.Y(n_1345)
);

NAND2xp33_ASAP7_75t_R g1346 ( 
.A(n_1316),
.B(n_794),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1274),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1296),
.Y(n_1348)
);

NOR2xp67_ASAP7_75t_L g1349 ( 
.A(n_1245),
.B(n_992),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1255),
.A2(n_1056),
.B1(n_1135),
.B2(n_1041),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1296),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1287),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1231),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1287),
.Y(n_1354)
);

CKINVDCx16_ASAP7_75t_R g1355 ( 
.A(n_1326),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1295),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1231),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1245),
.B(n_1221),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1295),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1280),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1238),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1233),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_1293),
.Y(n_1363)
);

CKINVDCx16_ASAP7_75t_R g1364 ( 
.A(n_1235),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1275),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_R g1366 ( 
.A(n_1262),
.B(n_984),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1328),
.Y(n_1367)
);

BUFx10_ASAP7_75t_L g1368 ( 
.A(n_1253),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1253),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1245),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_R g1371 ( 
.A(n_1307),
.B(n_1265),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_1242),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1265),
.Y(n_1373)
);

AND2x6_ASAP7_75t_L g1374 ( 
.A(n_1269),
.B(n_1204),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1265),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1294),
.Y(n_1376)
);

INVx11_ASAP7_75t_L g1377 ( 
.A(n_1242),
.Y(n_1377)
);

NOR2xp67_ASAP7_75t_L g1378 ( 
.A(n_1252),
.B(n_1144),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1294),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1269),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1278),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1278),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1228),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1321),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1258),
.Y(n_1385)
);

NOR2xp67_ASAP7_75t_L g1386 ( 
.A(n_1252),
.B(n_1174),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1258),
.B(n_921),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1284),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_1228),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1310),
.Y(n_1390)
);

NOR2xp67_ASAP7_75t_L g1391 ( 
.A(n_1325),
.B(n_882),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1308),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1308),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1317),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1234),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1246),
.B(n_1049),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1308),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1305),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1236),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1305),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1256),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1239),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1268),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1325),
.B(n_1219),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1291),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1327),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1238),
.Y(n_1407)
);

NOR2xp67_ASAP7_75t_L g1408 ( 
.A(n_1327),
.B(n_1309),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_R g1409 ( 
.A(n_1239),
.B(n_984),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1324),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1247),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1247),
.B(n_898),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1248),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1248),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1260),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1260),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1259),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1289),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1289),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1259),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1229),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1271),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1271),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1324),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1282),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1282),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1286),
.Y(n_1427)
);

NAND2xp33_ASAP7_75t_R g1428 ( 
.A(n_1323),
.B(n_795),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1286),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1299),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1299),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1313),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1313),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1237),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1240),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1241),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1250),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1254),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1257),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1261),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1263),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1264),
.Y(n_1442)
);

AND3x2_ASAP7_75t_L g1443 ( 
.A(n_1266),
.B(n_1179),
.C(n_1086),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_R g1444 ( 
.A(n_1309),
.B(n_1085),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1267),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1273),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1281),
.Y(n_1447)
);

CKINVDCx16_ASAP7_75t_R g1448 ( 
.A(n_1312),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_R g1449 ( 
.A(n_1315),
.B(n_1222),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1238),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1290),
.Y(n_1451)
);

CKINVDCx20_ASAP7_75t_R g1452 ( 
.A(n_1323),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1243),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1243),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1251),
.Y(n_1455)
);

CKINVDCx6p67_ASAP7_75t_R g1456 ( 
.A(n_1251),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1251),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_R g1458 ( 
.A(n_1270),
.B(n_801),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1270),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1270),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1276),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1276),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1276),
.Y(n_1463)
);

NOR2xp67_ASAP7_75t_L g1464 ( 
.A(n_1279),
.B(n_878),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1279),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1292),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1292),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1292),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1297),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1297),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1297),
.Y(n_1471)
);

CKINVDCx6p67_ASAP7_75t_R g1472 ( 
.A(n_1300),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1300),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1301),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_R g1475 ( 
.A(n_1301),
.B(n_820),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1301),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1302),
.B(n_826),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1302),
.B(n_898),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1302),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1303),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1303),
.Y(n_1481)
);

BUFx10_ASAP7_75t_L g1482 ( 
.A(n_1303),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1314),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1314),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1318),
.Y(n_1485)
);

NOR2xp67_ASAP7_75t_L g1486 ( 
.A(n_1324),
.B(n_976),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1318),
.Y(n_1487)
);

CKINVDCx16_ASAP7_75t_R g1488 ( 
.A(n_1322),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1322),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1230),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1319),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1296),
.B(n_1215),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_R g1493 ( 
.A(n_1244),
.B(n_923),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1230),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_R g1495 ( 
.A(n_1244),
.B(n_939),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1230),
.Y(n_1496)
);

NOR2xp67_ASAP7_75t_L g1497 ( 
.A(n_1245),
.B(n_980),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1230),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1230),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1238),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1230),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1319),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1272),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1227),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1385),
.B(n_1054),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1338),
.Y(n_1506)
);

NOR2xp67_ASAP7_75t_SL g1507 ( 
.A(n_1348),
.B(n_1178),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1351),
.B(n_1127),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1428),
.B(n_863),
.C(n_833),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1355),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1412),
.B(n_1180),
.Y(n_1511)
);

NOR2xp67_ASAP7_75t_L g1512 ( 
.A(n_1382),
.B(n_762),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_SL g1513 ( 
.A(n_1415),
.B(n_997),
.Y(n_1513)
);

BUFx5_ASAP7_75t_L g1514 ( 
.A(n_1451),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1387),
.B(n_884),
.Y(n_1515)
);

INVx4_ASAP7_75t_L g1516 ( 
.A(n_1488),
.Y(n_1516)
);

NOR3xp33_ASAP7_75t_L g1517 ( 
.A(n_1364),
.B(n_823),
.C(n_804),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_SL g1518 ( 
.A(n_1416),
.B(n_930),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1330),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1353),
.B(n_799),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1338),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1492),
.B(n_800),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1365),
.B(n_945),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1382),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1448),
.B(n_996),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1395),
.B(n_1002),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1331),
.B(n_896),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_1342),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1334),
.B(n_898),
.Y(n_1529)
);

XNOR2xp5_ASAP7_75t_L g1530 ( 
.A(n_1356),
.B(n_816),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1367),
.Y(n_1531)
);

INVxp67_ASAP7_75t_L g1532 ( 
.A(n_1503),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1491),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1368),
.B(n_1093),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1503),
.B(n_987),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1362),
.B(n_1002),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1502),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1478),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1369),
.B(n_1014),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1388),
.B(n_1093),
.Y(n_1540)
);

NAND2xp33_ASAP7_75t_SL g1541 ( 
.A(n_1409),
.B(n_816),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1504),
.B(n_1019),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1381),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1400),
.A2(n_796),
.B1(n_802),
.B2(n_793),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1390),
.B(n_1019),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1392),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1406),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1396),
.B(n_827),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1405),
.B(n_805),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1393),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1378),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1397),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1435),
.B(n_1080),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1394),
.B(n_1337),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1436),
.B(n_1080),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1386),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1437),
.B(n_1158),
.Y(n_1557)
);

OR2x6_ASAP7_75t_L g1558 ( 
.A(n_1343),
.B(n_965),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1438),
.B(n_1158),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1464),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_SL g1561 ( 
.A(n_1374),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1440),
.B(n_806),
.Y(n_1562)
);

NAND2xp33_ASAP7_75t_L g1563 ( 
.A(n_1374),
.B(n_930),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1434),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1357),
.B(n_808),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1486),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1441),
.B(n_811),
.Y(n_1567)
);

OR2x6_ASAP7_75t_L g1568 ( 
.A(n_1391),
.B(n_1081),
.Y(n_1568)
);

NAND2xp33_ASAP7_75t_L g1569 ( 
.A(n_1374),
.B(n_930),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1434),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1366),
.Y(n_1571)
);

INVxp67_ASAP7_75t_L g1572 ( 
.A(n_1346),
.Y(n_1572)
);

INVx8_ASAP7_75t_L g1573 ( 
.A(n_1374),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1340),
.A2(n_810),
.B(n_809),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1404),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1384),
.B(n_1130),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1442),
.B(n_812),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1421),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1335),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1408),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1349),
.Y(n_1581)
);

INVxp33_ASAP7_75t_L g1582 ( 
.A(n_1493),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1447),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1413),
.B(n_1130),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1497),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_L g1586 ( 
.A(n_1414),
.B(n_1134),
.C(n_851),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1445),
.B(n_813),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1417),
.B(n_1133),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1449),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1420),
.B(n_817),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1425),
.A2(n_897),
.B(n_843),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1426),
.B(n_1427),
.Y(n_1592)
);

NOR3xp33_ASAP7_75t_L g1593 ( 
.A(n_1329),
.B(n_880),
.C(n_874),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1429),
.B(n_818),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_SL g1595 ( 
.A(n_1377),
.Y(n_1595)
);

NOR2xp67_ASAP7_75t_L g1596 ( 
.A(n_1358),
.B(n_768),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1430),
.B(n_821),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1432),
.B(n_822),
.Y(n_1598)
);

NOR3xp33_ASAP7_75t_L g1599 ( 
.A(n_1376),
.B(n_1015),
.C(n_942),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1433),
.B(n_1443),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1352),
.B(n_1354),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1350),
.B(n_1401),
.Y(n_1602)
);

BUFx12f_ASAP7_75t_L g1603 ( 
.A(n_1332),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1443),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1358),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1359),
.B(n_1133),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1447),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1371),
.B(n_1133),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1370),
.B(n_828),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1335),
.B(n_987),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1373),
.B(n_832),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1339),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1375),
.B(n_834),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1482),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1399),
.B(n_1411),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1439),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1403),
.B(n_836),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1360),
.B(n_838),
.Y(n_1618)
);

INVx2_ASAP7_75t_SL g1619 ( 
.A(n_1495),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1402),
.B(n_839),
.Y(n_1620)
);

NAND2xp33_ASAP7_75t_L g1621 ( 
.A(n_1418),
.B(n_930),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1446),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1344),
.B(n_987),
.Y(n_1623)
);

AOI221xp5_ASAP7_75t_L g1624 ( 
.A1(n_1363),
.A2(n_862),
.B1(n_868),
.B2(n_857),
.C(n_850),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1482),
.Y(n_1625)
);

INVx2_ASAP7_75t_SL g1626 ( 
.A(n_1444),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1422),
.B(n_841),
.Y(n_1627)
);

NAND3xp33_ASAP7_75t_L g1628 ( 
.A(n_1423),
.B(n_875),
.C(n_871),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1431),
.B(n_842),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1477),
.B(n_1458),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_1484),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1345),
.B(n_1076),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_L g1633 ( 
.A(n_1456),
.Y(n_1633)
);

NAND3xp33_ASAP7_75t_L g1634 ( 
.A(n_1419),
.B(n_900),
.C(n_885),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1475),
.B(n_845),
.Y(n_1635)
);

AND2x2_ASAP7_75t_SL g1636 ( 
.A(n_1347),
.B(n_843),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1452),
.A2(n_901),
.B1(n_905),
.B2(n_903),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1472),
.Y(n_1638)
);

NOR2x1p5_ASAP7_75t_L g1639 ( 
.A(n_1333),
.B(n_846),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1454),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1455),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1336),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1462),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1463),
.B(n_848),
.Y(n_1644)
);

AND2x6_ASAP7_75t_L g1645 ( 
.A(n_1474),
.B(n_897),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1465),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1466),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1383),
.A2(n_910),
.B1(n_918),
.B2(n_909),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1467),
.B(n_852),
.Y(n_1649)
);

NOR3xp33_ASAP7_75t_L g1650 ( 
.A(n_1379),
.B(n_1050),
.C(n_1024),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1468),
.B(n_853),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1469),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1470),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1471),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1341),
.B(n_854),
.Y(n_1655)
);

NOR3xp33_ASAP7_75t_L g1656 ( 
.A(n_1490),
.B(n_1113),
.C(n_1100),
.Y(n_1656)
);

CKINVDCx20_ASAP7_75t_R g1657 ( 
.A(n_1372),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1480),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1494),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1483),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1389),
.B(n_856),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_SL g1662 ( 
.A(n_1496),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1485),
.B(n_858),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1498),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_SL g1665 ( 
.A(n_1499),
.B(n_930),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1487),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1398),
.B(n_860),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1489),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1476),
.Y(n_1669)
);

BUFx6f_ASAP7_75t_L g1670 ( 
.A(n_1361),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1501),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1457),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1457),
.B(n_864),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1453),
.B(n_1171),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1460),
.B(n_865),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1461),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1361),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1473),
.B(n_867),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1479),
.B(n_869),
.Y(n_1679)
);

NOR3xp33_ASAP7_75t_L g1680 ( 
.A(n_1481),
.B(n_1187),
.C(n_1173),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1450),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1459),
.B(n_870),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1407),
.B(n_872),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1407),
.B(n_873),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1407),
.B(n_877),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1410),
.B(n_879),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1410),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1410),
.B(n_881),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_SL g1689 ( 
.A(n_1424),
.B(n_1189),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1424),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1424),
.B(n_883),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1500),
.B(n_886),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1500),
.Y(n_1693)
);

NOR3xp33_ASAP7_75t_L g1694 ( 
.A(n_1500),
.B(n_888),
.C(n_887),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1385),
.B(n_889),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1380),
.A2(n_931),
.B1(n_935),
.B2(n_933),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1387),
.B(n_890),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1387),
.B(n_891),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1385),
.B(n_892),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1385),
.B(n_893),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1385),
.B(n_894),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1503),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1385),
.B(n_1076),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1385),
.B(n_899),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1385),
.B(n_1206),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1385),
.B(n_902),
.Y(n_1706)
);

A2O1A1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1380),
.A2(n_936),
.B(n_946),
.C(n_944),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1385),
.B(n_904),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1385),
.B(n_906),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_SL g1710 ( 
.A(n_1415),
.B(n_930),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1330),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1385),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1385),
.B(n_907),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1503),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1385),
.B(n_911),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1330),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1385),
.B(n_1206),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1385),
.B(n_1076),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1503),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1338),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1385),
.B(n_913),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1385),
.B(n_915),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1385),
.B(n_917),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1330),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1385),
.B(n_1182),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1338),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1385),
.B(n_920),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1330),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1385),
.B(n_922),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1330),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1387),
.B(n_925),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1385),
.B(n_927),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1385),
.B(n_929),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1355),
.B(n_1226),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_SL g1735 ( 
.A(n_1415),
.B(n_1035),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1338),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1385),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1387),
.B(n_932),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1387),
.B(n_937),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1385),
.B(n_1206),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1338),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1385),
.B(n_940),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1330),
.Y(n_1743)
);

INVx2_ASAP7_75t_SL g1744 ( 
.A(n_1385),
.Y(n_1744)
);

OR2x6_ASAP7_75t_L g1745 ( 
.A(n_1343),
.B(n_914),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1387),
.B(n_941),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1338),
.Y(n_1747)
);

NOR3xp33_ASAP7_75t_L g1748 ( 
.A(n_1355),
.B(n_948),
.C(n_947),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1712),
.B(n_951),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1564),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1570),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1633),
.B(n_949),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1575),
.B(n_950),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1532),
.B(n_837),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1702),
.B(n_844),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1510),
.Y(n_1756)
);

INVx5_ASAP7_75t_L g1757 ( 
.A(n_1633),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1521),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1633),
.B(n_1737),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1744),
.B(n_1592),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1516),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1543),
.B(n_954),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1745),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1528),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1573),
.Y(n_1765)
);

NOR2x2_ASAP7_75t_L g1766 ( 
.A(n_1745),
.B(n_951),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1714),
.B(n_956),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1719),
.B(n_955),
.Y(n_1768)
);

INVx2_ASAP7_75t_SL g1769 ( 
.A(n_1745),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1573),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1516),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1548),
.B(n_958),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1697),
.B(n_961),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1603),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1662),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1698),
.B(n_962),
.Y(n_1776)
);

INVx2_ASAP7_75t_SL g1777 ( 
.A(n_1631),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1642),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1731),
.B(n_964),
.Y(n_1779)
);

NOR2x1_ASAP7_75t_R g1780 ( 
.A(n_1671),
.B(n_966),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1529),
.A2(n_968),
.B1(n_969),
.B2(n_967),
.Y(n_1781)
);

AO22x1_ASAP7_75t_L g1782 ( 
.A1(n_1571),
.A2(n_959),
.B1(n_970),
.B2(n_955),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1602),
.B(n_849),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1720),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1738),
.B(n_979),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1538),
.B(n_952),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1513),
.A2(n_985),
.B1(n_986),
.B2(n_981),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1547),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1739),
.B(n_988),
.Y(n_1789)
);

BUFx6f_ASAP7_75t_L g1790 ( 
.A(n_1573),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1726),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1736),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1645),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1741),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1746),
.B(n_990),
.Y(n_1795)
);

NOR3xp33_ASAP7_75t_SL g1796 ( 
.A(n_1661),
.B(n_995),
.C(n_993),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1525),
.B(n_1515),
.Y(n_1797)
);

BUFx3_ASAP7_75t_L g1798 ( 
.A(n_1664),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1747),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1511),
.B(n_998),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1506),
.B(n_999),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1524),
.Y(n_1802)
);

AOI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1513),
.A2(n_1008),
.B1(n_1010),
.B2(n_1001),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1589),
.B(n_1011),
.Y(n_1804)
);

BUFx2_ASAP7_75t_L g1805 ( 
.A(n_1734),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1695),
.B(n_1012),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1703),
.B(n_908),
.Y(n_1807)
);

INVxp67_ASAP7_75t_L g1808 ( 
.A(n_1718),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1725),
.B(n_959),
.Y(n_1809)
);

BUFx3_ASAP7_75t_L g1810 ( 
.A(n_1579),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1637),
.A2(n_982),
.B1(n_994),
.B2(n_970),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1604),
.B(n_953),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1616),
.Y(n_1813)
);

INVx2_ASAP7_75t_SL g1814 ( 
.A(n_1610),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1638),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1643),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1699),
.B(n_1700),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1634),
.A2(n_994),
.B1(n_1006),
.B2(n_982),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1541),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1622),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1505),
.B(n_1016),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_1645),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1585),
.B(n_957),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_SL g1824 ( 
.A1(n_1636),
.A2(n_1218),
.B1(n_1007),
.B2(n_1104),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1530),
.A2(n_1007),
.B1(n_1104),
.B2(n_1006),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1519),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1531),
.Y(n_1827)
);

BUFx5_ASAP7_75t_L g1828 ( 
.A(n_1645),
.Y(n_1828)
);

INVx2_ASAP7_75t_SL g1829 ( 
.A(n_1652),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1701),
.B(n_1023),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_R g1831 ( 
.A(n_1619),
.B(n_1123),
.Y(n_1831)
);

BUFx8_ASAP7_75t_L g1832 ( 
.A(n_1662),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1533),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1634),
.A2(n_963),
.B1(n_972),
.B2(n_960),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1704),
.B(n_1025),
.Y(n_1835)
);

INVx2_ASAP7_75t_SL g1836 ( 
.A(n_1653),
.Y(n_1836)
);

AND2x4_ASAP7_75t_SL g1837 ( 
.A(n_1535),
.B(n_1182),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1593),
.A2(n_974),
.B1(n_977),
.B2(n_975),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1549),
.B(n_1212),
.Y(n_1839)
);

NAND2x1p5_ASAP7_75t_L g1840 ( 
.A(n_1601),
.B(n_1003),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1537),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1706),
.A2(n_1029),
.B1(n_1030),
.B2(n_1028),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1612),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1595),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1708),
.B(n_1031),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1709),
.B(n_1034),
.Y(n_1846)
);

OR2x6_ASAP7_75t_L g1847 ( 
.A(n_1659),
.B(n_983),
.Y(n_1847)
);

AND2x6_ASAP7_75t_SL g1848 ( 
.A(n_1667),
.B(n_1004),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1711),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1713),
.B(n_1038),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1716),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1670),
.Y(n_1852)
);

BUFx8_ASAP7_75t_L g1853 ( 
.A(n_1595),
.Y(n_1853)
);

INVx3_ASAP7_75t_L g1854 ( 
.A(n_1653),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1715),
.B(n_912),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1600),
.B(n_1040),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1590),
.B(n_1044),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1721),
.B(n_1045),
.Y(n_1858)
);

INVx5_ASAP7_75t_L g1859 ( 
.A(n_1626),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1724),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_SL g1861 ( 
.A1(n_1561),
.A2(n_928),
.B1(n_1027),
.B2(n_924),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1581),
.B(n_1005),
.Y(n_1862)
);

NAND3xp33_ASAP7_75t_SL g1863 ( 
.A(n_1656),
.B(n_1064),
.C(n_1046),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1728),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1509),
.A2(n_1586),
.B1(n_1605),
.B2(n_1628),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1617),
.B(n_1182),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1730),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_R g1868 ( 
.A(n_1657),
.B(n_1103),
.Y(n_1868)
);

BUFx3_ASAP7_75t_L g1869 ( 
.A(n_1614),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1722),
.B(n_1090),
.Y(n_1870)
);

O2A1O1Ixp5_ASAP7_75t_L g1871 ( 
.A1(n_1584),
.A2(n_1070),
.B(n_1082),
.C(n_983),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1723),
.B(n_1098),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1623),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1743),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1594),
.B(n_1048),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1578),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_1632),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1554),
.B(n_1220),
.Y(n_1878)
);

INVx2_ASAP7_75t_SL g1879 ( 
.A(n_1674),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1583),
.Y(n_1880)
);

NAND2xp33_ASAP7_75t_L g1881 ( 
.A(n_1514),
.B(n_1035),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_SL g1882 ( 
.A1(n_1655),
.A2(n_1183),
.B1(n_1195),
.B2(n_1149),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1526),
.Y(n_1883)
);

INVx5_ASAP7_75t_L g1884 ( 
.A(n_1625),
.Y(n_1884)
);

INVx5_ASAP7_75t_L g1885 ( 
.A(n_1568),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1646),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1536),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1727),
.B(n_1052),
.Y(n_1888)
);

INVx3_ASAP7_75t_L g1889 ( 
.A(n_1607),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1615),
.A2(n_1013),
.B1(n_1017),
.B2(n_1009),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1546),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1539),
.Y(n_1892)
);

BUFx2_ASAP7_75t_L g1893 ( 
.A(n_1729),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1509),
.A2(n_1021),
.B1(n_1022),
.B2(n_1020),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1542),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1732),
.B(n_1053),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1550),
.Y(n_1897)
);

BUFx6f_ASAP7_75t_L g1898 ( 
.A(n_1670),
.Y(n_1898)
);

INVx2_ASAP7_75t_SL g1899 ( 
.A(n_1647),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1552),
.Y(n_1900)
);

CKINVDCx11_ASAP7_75t_R g1901 ( 
.A(n_1558),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1670),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1572),
.B(n_1026),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1733),
.B(n_1055),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1545),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1523),
.Y(n_1906)
);

CKINVDCx20_ASAP7_75t_R g1907 ( 
.A(n_1618),
.Y(n_1907)
);

OAI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1544),
.A2(n_1742),
.B1(n_1710),
.B2(n_1735),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1620),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1591),
.B(n_1627),
.Y(n_1910)
);

AOI21x1_ASAP7_75t_L g1911 ( 
.A1(n_1512),
.A2(n_1036),
.B(n_1032),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1544),
.B(n_1220),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1629),
.B(n_1522),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1560),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1566),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1580),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1574),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1648),
.B(n_1220),
.Y(n_1918)
);

NAND3xp33_ASAP7_75t_SL g1919 ( 
.A(n_1624),
.B(n_1209),
.C(n_1208),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1683),
.Y(n_1920)
);

AND2x6_ASAP7_75t_L g1921 ( 
.A(n_1561),
.B(n_1070),
.Y(n_1921)
);

AOI22xp33_ASAP7_75t_L g1922 ( 
.A1(n_1586),
.A2(n_1037),
.B1(n_1042),
.B2(n_1039),
.Y(n_1922)
);

OR2x2_ASAP7_75t_SL g1923 ( 
.A(n_1639),
.B(n_1043),
.Y(n_1923)
);

INVx4_ASAP7_75t_L g1924 ( 
.A(n_1558),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1684),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1686),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1597),
.B(n_1057),
.Y(n_1927)
);

INVx3_ASAP7_75t_L g1928 ( 
.A(n_1527),
.Y(n_1928)
);

INVx5_ASAP7_75t_L g1929 ( 
.A(n_1568),
.Y(n_1929)
);

OR2x4_ASAP7_75t_L g1930 ( 
.A(n_1565),
.B(n_1051),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1691),
.Y(n_1931)
);

BUFx6f_ASAP7_75t_L g1932 ( 
.A(n_1677),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1598),
.B(n_1058),
.Y(n_1933)
);

BUFx3_ASAP7_75t_L g1934 ( 
.A(n_1654),
.Y(n_1934)
);

BUFx6f_ASAP7_75t_L g1935 ( 
.A(n_1677),
.Y(n_1935)
);

BUFx6f_ASAP7_75t_L g1936 ( 
.A(n_1677),
.Y(n_1936)
);

OR2x6_ASAP7_75t_L g1937 ( 
.A(n_1558),
.B(n_1082),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1562),
.B(n_1059),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1527),
.Y(n_1939)
);

BUFx2_ASAP7_75t_L g1940 ( 
.A(n_1567),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1692),
.Y(n_1941)
);

NOR3xp33_ASAP7_75t_SL g1942 ( 
.A(n_1707),
.B(n_1062),
.C(n_1061),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1628),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1512),
.B(n_1577),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1551),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1556),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1673),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1696),
.B(n_1065),
.Y(n_1948)
);

INVx5_ASAP7_75t_L g1949 ( 
.A(n_1568),
.Y(n_1949)
);

NAND2xp33_ASAP7_75t_SL g1950 ( 
.A(n_1582),
.B(n_1211),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1668),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1517),
.A2(n_1071),
.B1(n_1072),
.B2(n_1066),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1587),
.B(n_1073),
.Y(n_1953)
);

BUFx6f_ASAP7_75t_L g1954 ( 
.A(n_1669),
.Y(n_1954)
);

AOI22xp33_ASAP7_75t_L g1955 ( 
.A1(n_1748),
.A2(n_1063),
.B1(n_1069),
.B2(n_1068),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1640),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1665),
.B(n_1514),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1534),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1553),
.B(n_1555),
.Y(n_1959)
);

BUFx12f_ASAP7_75t_L g1960 ( 
.A(n_1665),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1689),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1611),
.B(n_1079),
.Y(n_1962)
);

INVx3_ASAP7_75t_L g1963 ( 
.A(n_1641),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1694),
.A2(n_1075),
.B1(n_1078),
.B2(n_1077),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1609),
.B(n_1613),
.Y(n_1965)
);

AOI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1563),
.A2(n_1569),
.B(n_1559),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1675),
.Y(n_1967)
);

INVx1_ASAP7_75t_SL g1968 ( 
.A(n_1644),
.Y(n_1968)
);

BUFx3_ASAP7_75t_L g1969 ( 
.A(n_1658),
.Y(n_1969)
);

INVx3_ASAP7_75t_L g1970 ( 
.A(n_1660),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1514),
.B(n_1083),
.Y(n_1971)
);

AND2x6_ASAP7_75t_L g1972 ( 
.A(n_1666),
.B(n_1117),
.Y(n_1972)
);

INVx3_ASAP7_75t_L g1973 ( 
.A(n_1649),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1557),
.B(n_1088),
.Y(n_1974)
);

AOI22xp33_ASAP7_75t_L g1975 ( 
.A1(n_1680),
.A2(n_1087),
.B1(n_1096),
.B2(n_1095),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1520),
.B(n_1091),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1740),
.B(n_1092),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1599),
.B(n_1094),
.Y(n_1978)
);

OR2x6_ASAP7_75t_L g1979 ( 
.A(n_1606),
.B(n_1117),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1540),
.B(n_1097),
.Y(n_1980)
);

NOR2x1_ASAP7_75t_R g1981 ( 
.A(n_1635),
.B(n_1102),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1705),
.B(n_1105),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1717),
.A2(n_1109),
.B1(n_1110),
.B2(n_1108),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1507),
.B(n_1106),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1651),
.B(n_1107),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1621),
.A2(n_1114),
.B1(n_1115),
.B2(n_1111),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1676),
.Y(n_1987)
);

AOI22xp33_ASAP7_75t_L g1988 ( 
.A1(n_1588),
.A2(n_1735),
.B1(n_1518),
.B2(n_1710),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1685),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1688),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1682),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1663),
.A2(n_1122),
.B1(n_1124),
.B2(n_1121),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1508),
.B(n_1116),
.Y(n_1993)
);

AOI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1576),
.A2(n_1678),
.B1(n_1679),
.B2(n_1650),
.Y(n_1994)
);

INVx3_ASAP7_75t_L g1995 ( 
.A(n_1681),
.Y(n_1995)
);

INVxp67_ASAP7_75t_L g1996 ( 
.A(n_1608),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1596),
.B(n_1118),
.Y(n_1997)
);

INVx2_ASAP7_75t_SL g1998 ( 
.A(n_1630),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1672),
.B(n_1125),
.Y(n_1999)
);

BUFx4f_ASAP7_75t_L g2000 ( 
.A(n_1690),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1687),
.Y(n_2001)
);

BUFx3_ASAP7_75t_L g2002 ( 
.A(n_1693),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1564),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1564),
.B(n_1128),
.Y(n_2004)
);

AND2x6_ASAP7_75t_L g2005 ( 
.A(n_1573),
.B(n_1132),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1510),
.Y(n_2006)
);

NOR2xp67_ASAP7_75t_L g2007 ( 
.A(n_1579),
.B(n_22),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1564),
.B(n_1129),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1532),
.B(n_1131),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1564),
.B(n_1137),
.Y(n_2010)
);

BUFx6f_ASAP7_75t_L g2011 ( 
.A(n_1573),
.Y(n_2011)
);

OR2x6_ASAP7_75t_L g2012 ( 
.A(n_1510),
.B(n_1132),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1564),
.B(n_1142),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1564),
.B(n_1143),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1510),
.Y(n_2015)
);

INVx5_ASAP7_75t_L g2016 ( 
.A(n_1633),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1564),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_1575),
.B(n_1126),
.Y(n_2018)
);

INVxp67_ASAP7_75t_SL g2019 ( 
.A(n_1510),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1633),
.B(n_1146),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1712),
.B(n_1147),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_1633),
.B(n_1148),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1506),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1712),
.B(n_1150),
.Y(n_2024)
);

BUFx3_ASAP7_75t_L g2025 ( 
.A(n_1633),
.Y(n_2025)
);

NOR2x1p5_ASAP7_75t_L g2026 ( 
.A(n_1603),
.B(n_1157),
.Y(n_2026)
);

AOI22xp5_ASAP7_75t_L g2027 ( 
.A1(n_2018),
.A2(n_1154),
.B1(n_1155),
.B2(n_1152),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1756),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1757),
.B(n_1216),
.Y(n_2029)
);

A2O1A1Ixp33_ASAP7_75t_L g2030 ( 
.A1(n_1910),
.A2(n_1136),
.B(n_1139),
.C(n_1138),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1912),
.B(n_1161),
.Y(n_2031)
);

A2O1A1Ixp33_ASAP7_75t_L g2032 ( 
.A1(n_1913),
.A2(n_1140),
.B(n_1145),
.C(n_1141),
.Y(n_2032)
);

BUFx12f_ASAP7_75t_L g2033 ( 
.A(n_1832),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1750),
.Y(n_2034)
);

INVx3_ASAP7_75t_L g2035 ( 
.A(n_1765),
.Y(n_2035)
);

INVx2_ASAP7_75t_SL g2036 ( 
.A(n_1757),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1808),
.B(n_1162),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1757),
.B(n_1205),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1813),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1797),
.B(n_1164),
.Y(n_2040)
);

AOI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_1817),
.A2(n_1153),
.B(n_1151),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1959),
.A2(n_1163),
.B(n_1159),
.Y(n_2042)
);

AOI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_1881),
.A2(n_1167),
.B(n_1165),
.Y(n_2043)
);

INVx5_ASAP7_75t_L g2044 ( 
.A(n_2005),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1909),
.B(n_1166),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1751),
.B(n_1168),
.Y(n_2046)
);

OAI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_2018),
.A2(n_1908),
.B1(n_1879),
.B2(n_1986),
.Y(n_2047)
);

NOR3xp33_ASAP7_75t_L g2048 ( 
.A(n_1863),
.B(n_1225),
.C(n_1223),
.Y(n_2048)
);

O2A1O1Ixp33_ASAP7_75t_L g2049 ( 
.A1(n_1992),
.A2(n_1176),
.B(n_1186),
.C(n_1175),
.Y(n_2049)
);

AOI21xp5_ASAP7_75t_L g2050 ( 
.A1(n_1966),
.A2(n_1200),
.B(n_1194),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_1811),
.B(n_1169),
.Y(n_2051)
);

AOI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_1957),
.A2(n_1202),
.B(n_1201),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1852),
.Y(n_2053)
);

NOR2x1_ASAP7_75t_R g2054 ( 
.A(n_1901),
.B(n_1170),
.Y(n_2054)
);

NOR2xp67_ASAP7_75t_L g2055 ( 
.A(n_2016),
.B(n_771),
.Y(n_2055)
);

BUFx8_ASAP7_75t_L g2056 ( 
.A(n_1774),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1768),
.B(n_1172),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_1906),
.B(n_1973),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2003),
.B(n_1181),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_2017),
.B(n_1820),
.Y(n_2060)
);

BUFx2_ASAP7_75t_L g2061 ( 
.A(n_2006),
.Y(n_2061)
);

NOR3xp33_ASAP7_75t_SL g2062 ( 
.A(n_1775),
.B(n_1185),
.C(n_1184),
.Y(n_2062)
);

BUFx12f_ASAP7_75t_L g2063 ( 
.A(n_1832),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1826),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_SL g2065 ( 
.A(n_1780),
.B(n_1188),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1997),
.A2(n_1210),
.B(n_1207),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1827),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1833),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1841),
.Y(n_2069)
);

A2O1A1Ixp33_ASAP7_75t_SL g2070 ( 
.A1(n_1976),
.A2(n_1213),
.B(n_1203),
.C(n_1191),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1987),
.Y(n_2071)
);

NOR2x1_ASAP7_75t_L g2072 ( 
.A(n_1883),
.B(n_1203),
.Y(n_2072)
);

INVx5_ASAP7_75t_L g2073 ( 
.A(n_2005),
.Y(n_2073)
);

BUFx4f_ASAP7_75t_L g2074 ( 
.A(n_2005),
.Y(n_2074)
);

OR2x6_ASAP7_75t_L g2075 ( 
.A(n_1782),
.B(n_1213),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1753),
.A2(n_1193),
.B(n_1192),
.Y(n_2076)
);

NOR2xp33_ASAP7_75t_L g2077 ( 
.A(n_1807),
.B(n_1196),
.Y(n_2077)
);

INVxp67_ASAP7_75t_L g2078 ( 
.A(n_1843),
.Y(n_2078)
);

INVxp67_ASAP7_75t_L g2079 ( 
.A(n_2019),
.Y(n_2079)
);

O2A1O1Ixp33_ASAP7_75t_L g2080 ( 
.A1(n_1919),
.A2(n_1772),
.B(n_1818),
.C(n_1890),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_R g2081 ( 
.A(n_1764),
.B(n_1198),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_1853),
.Y(n_2082)
);

INVx5_ASAP7_75t_L g2083 ( 
.A(n_2005),
.Y(n_2083)
);

O2A1O1Ixp33_ASAP7_75t_L g2084 ( 
.A1(n_1991),
.A2(n_1217),
.B(n_1199),
.C(n_1214),
.Y(n_2084)
);

AOI21xp5_ASAP7_75t_L g2085 ( 
.A1(n_1967),
.A2(n_1214),
.B(n_1206),
.Y(n_2085)
);

BUFx12f_ASAP7_75t_L g2086 ( 
.A(n_1853),
.Y(n_2086)
);

CKINVDCx20_ASAP7_75t_R g2087 ( 
.A(n_1868),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1894),
.B(n_1214),
.Y(n_2088)
);

O2A1O1Ixp33_ASAP7_75t_L g2089 ( 
.A1(n_1989),
.A2(n_1990),
.B(n_1918),
.C(n_1776),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1849),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1968),
.B(n_25),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_1831),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_1947),
.B(n_26),
.Y(n_2093)
);

AOI221xp5_ASAP7_75t_L g2094 ( 
.A1(n_1838),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.C(n_30),
.Y(n_2094)
);

BUFx12f_ASAP7_75t_L g2095 ( 
.A(n_1844),
.Y(n_2095)
);

O2A1O1Ixp33_ASAP7_75t_L g2096 ( 
.A1(n_1773),
.A2(n_30),
.B(n_27),
.C(n_28),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1851),
.Y(n_2097)
);

HB1xp67_ASAP7_75t_L g2098 ( 
.A(n_1798),
.Y(n_2098)
);

BUFx6f_ASAP7_75t_L g2099 ( 
.A(n_1852),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_L g2100 ( 
.A(n_1855),
.B(n_31),
.Y(n_2100)
);

NOR3xp33_ASAP7_75t_SL g2101 ( 
.A(n_1825),
.B(n_32),
.C(n_33),
.Y(n_2101)
);

HB1xp67_ASAP7_75t_L g2102 ( 
.A(n_2015),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1893),
.B(n_33),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_1783),
.A2(n_1035),
.B1(n_36),
.B2(n_34),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_1870),
.B(n_35),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_1749),
.B(n_37),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1940),
.B(n_37),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_1763),
.B(n_38),
.Y(n_2108)
);

AOI21xp5_ASAP7_75t_L g2109 ( 
.A1(n_1971),
.A2(n_776),
.B(n_772),
.Y(n_2109)
);

NOR2xp33_ASAP7_75t_R g2110 ( 
.A(n_1950),
.B(n_38),
.Y(n_2110)
);

BUFx3_ASAP7_75t_L g2111 ( 
.A(n_2025),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1887),
.B(n_1892),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1769),
.B(n_39),
.Y(n_2113)
);

O2A1O1Ixp33_ASAP7_75t_L g2114 ( 
.A1(n_1779),
.A2(n_45),
.B(n_42),
.C(n_44),
.Y(n_2114)
);

INVx1_ASAP7_75t_SL g2115 ( 
.A(n_1766),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1809),
.B(n_46),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1895),
.B(n_1905),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1922),
.B(n_46),
.Y(n_2118)
);

INVxp67_ASAP7_75t_L g2119 ( 
.A(n_2012),
.Y(n_2119)
);

BUFx4f_ASAP7_75t_SL g2120 ( 
.A(n_1778),
.Y(n_2120)
);

O2A1O1Ixp33_ASAP7_75t_L g2121 ( 
.A1(n_1785),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1860),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_1872),
.B(n_49),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1786),
.B(n_50),
.Y(n_2124)
);

BUFx8_ASAP7_75t_SL g2125 ( 
.A(n_2012),
.Y(n_2125)
);

INVx3_ASAP7_75t_L g2126 ( 
.A(n_1765),
.Y(n_2126)
);

BUFx2_ASAP7_75t_L g2127 ( 
.A(n_1788),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1786),
.B(n_50),
.Y(n_2128)
);

OAI22x1_ASAP7_75t_L g2129 ( 
.A1(n_2026),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_2129)
);

OR2x6_ASAP7_75t_L g2130 ( 
.A(n_1924),
.B(n_51),
.Y(n_2130)
);

O2A1O1Ixp33_ASAP7_75t_L g2131 ( 
.A1(n_1789),
.A2(n_1795),
.B(n_1800),
.C(n_1948),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1864),
.Y(n_2132)
);

NOR3xp33_ASAP7_75t_SL g2133 ( 
.A(n_1882),
.B(n_52),
.C(n_53),
.Y(n_2133)
);

NAND2x1_ASAP7_75t_SL g2134 ( 
.A(n_1754),
.B(n_54),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_1898),
.Y(n_2135)
);

NAND2x1p5_ASAP7_75t_L g2136 ( 
.A(n_1761),
.B(n_1771),
.Y(n_2136)
);

A2O1A1Ixp33_ASAP7_75t_SL g2137 ( 
.A1(n_1896),
.A2(n_784),
.B(n_786),
.C(n_780),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1824),
.B(n_55),
.Y(n_2138)
);

O2A1O1Ixp33_ASAP7_75t_L g2139 ( 
.A1(n_1920),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_2139)
);

NOR2xp33_ASAP7_75t_L g2140 ( 
.A(n_1755),
.B(n_56),
.Y(n_2140)
);

AOI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_1834),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_SL g2142 ( 
.A(n_1960),
.B(n_59),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1812),
.B(n_60),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1812),
.B(n_61),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_1814),
.B(n_745),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1925),
.B(n_62),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1926),
.B(n_62),
.Y(n_2147)
);

AND2x4_ASAP7_75t_L g2148 ( 
.A(n_1969),
.B(n_63),
.Y(n_2148)
);

NOR2xp33_ASAP7_75t_L g2149 ( 
.A(n_1805),
.B(n_64),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1931),
.B(n_66),
.Y(n_2150)
);

CKINVDCx20_ASAP7_75t_R g2151 ( 
.A(n_1907),
.Y(n_2151)
);

AO22x2_ASAP7_75t_L g2152 ( 
.A1(n_1924),
.A2(n_735),
.B1(n_736),
.B2(n_734),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_SL g2153 ( 
.A(n_1981),
.B(n_69),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_R g2154 ( 
.A(n_1819),
.B(n_734),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1867),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1965),
.B(n_70),
.Y(n_2156)
);

BUFx12f_ASAP7_75t_L g2157 ( 
.A(n_1777),
.Y(n_2157)
);

INVx8_ASAP7_75t_L g2158 ( 
.A(n_1921),
.Y(n_2158)
);

BUFx2_ASAP7_75t_L g2159 ( 
.A(n_1847),
.Y(n_2159)
);

INVx3_ASAP7_75t_L g2160 ( 
.A(n_1765),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1972),
.B(n_70),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1878),
.B(n_71),
.Y(n_2162)
);

A2O1A1Ixp33_ASAP7_75t_L g2163 ( 
.A1(n_1943),
.A2(n_1941),
.B(n_1904),
.C(n_1938),
.Y(n_2163)
);

O2A1O1Ixp33_ASAP7_75t_L g2164 ( 
.A1(n_1806),
.A2(n_74),
.B(n_71),
.C(n_73),
.Y(n_2164)
);

OAI22xp5_ASAP7_75t_L g2165 ( 
.A1(n_1822),
.A2(n_80),
.B1(n_75),
.B2(n_79),
.Y(n_2165)
);

A2O1A1Ixp33_ASAP7_75t_L g2166 ( 
.A1(n_1871),
.A2(n_1784),
.B(n_1791),
.C(n_1758),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1972),
.B(n_79),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1792),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1902),
.Y(n_2169)
);

INVx3_ASAP7_75t_L g2170 ( 
.A(n_1770),
.Y(n_2170)
);

NOR2xp33_ASAP7_75t_L g2171 ( 
.A(n_1873),
.B(n_82),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2021),
.B(n_82),
.Y(n_2172)
);

NAND3xp33_ASAP7_75t_L g2173 ( 
.A(n_1942),
.B(n_83),
.C(n_85),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_1877),
.B(n_727),
.Y(n_2174)
);

AOI22xp33_ASAP7_75t_L g2175 ( 
.A1(n_1839),
.A2(n_86),
.B1(n_83),
.B2(n_85),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1972),
.B(n_87),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1794),
.Y(n_2177)
);

AOI22xp5_ASAP7_75t_L g2178 ( 
.A1(n_1903),
.A2(n_1975),
.B1(n_1823),
.B2(n_1972),
.Y(n_2178)
);

INVx5_ASAP7_75t_L g2179 ( 
.A(n_1921),
.Y(n_2179)
);

A2O1A1Ixp33_ASAP7_75t_SL g2180 ( 
.A1(n_2009),
.A2(n_733),
.B(n_735),
.C(n_732),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_L g2181 ( 
.A(n_1837),
.B(n_732),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_1816),
.B(n_88),
.Y(n_2182)
);

AOI21xp5_ASAP7_75t_L g2183 ( 
.A1(n_1932),
.A2(n_89),
.B(n_90),
.Y(n_2183)
);

BUFx2_ASAP7_75t_L g2184 ( 
.A(n_1847),
.Y(n_2184)
);

AOI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_1935),
.A2(n_89),
.B(n_91),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_L g2186 ( 
.A(n_1866),
.B(n_741),
.Y(n_2186)
);

AOI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_1935),
.A2(n_94),
.B(n_97),
.Y(n_2187)
);

OAI22x1_ASAP7_75t_L g2188 ( 
.A1(n_1885),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1874),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_L g2190 ( 
.A(n_1760),
.B(n_746),
.Y(n_2190)
);

OAI22x1_ASAP7_75t_L g2191 ( 
.A1(n_1885),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_2191)
);

INVx4_ASAP7_75t_L g2192 ( 
.A(n_1921),
.Y(n_2192)
);

INVx5_ASAP7_75t_L g2193 ( 
.A(n_1921),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1799),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1802),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1891),
.Y(n_2196)
);

INVx1_ASAP7_75t_SL g2197 ( 
.A(n_2024),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_SL g2198 ( 
.A(n_1829),
.B(n_103),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_SL g2199 ( 
.A(n_1787),
.B(n_1803),
.Y(n_2199)
);

A2O1A1Ixp33_ASAP7_75t_L g2200 ( 
.A1(n_1762),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_2200)
);

NOR2xp67_ASAP7_75t_L g2201 ( 
.A(n_1889),
.B(n_104),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1897),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1903),
.B(n_107),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1956),
.B(n_108),
.Y(n_2204)
);

AOI21xp5_ASAP7_75t_L g2205 ( 
.A1(n_1936),
.A2(n_108),
.B(n_109),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1900),
.Y(n_2206)
);

INVx3_ASAP7_75t_L g2207 ( 
.A(n_1770),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1876),
.Y(n_2208)
);

NAND2x1p5_ASAP7_75t_L g2209 ( 
.A(n_1859),
.B(n_112),
.Y(n_2209)
);

OAI22xp33_ASAP7_75t_L g2210 ( 
.A1(n_1930),
.A2(n_114),
.B1(n_110),
.B2(n_113),
.Y(n_2210)
);

AOI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_1781),
.A2(n_1962),
.B1(n_1861),
.B2(n_1952),
.Y(n_2211)
);

NAND2xp33_ASAP7_75t_SL g2212 ( 
.A(n_1770),
.B(n_745),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1823),
.Y(n_2213)
);

NAND2x1p5_ASAP7_75t_L g2214 ( 
.A(n_1859),
.B(n_116),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_1848),
.Y(n_2215)
);

CKINVDCx5p33_ASAP7_75t_R g2216 ( 
.A(n_1796),
.Y(n_2216)
);

INVx1_ASAP7_75t_SL g2217 ( 
.A(n_1884),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1914),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1963),
.B(n_115),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1915),
.Y(n_2220)
);

OAI22xp5_ASAP7_75t_SL g2221 ( 
.A1(n_1923),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_2221)
);

AOI21xp5_ASAP7_75t_L g2222 ( 
.A1(n_1974),
.A2(n_120),
.B(n_121),
.Y(n_2222)
);

OAI22xp5_ASAP7_75t_SL g2223 ( 
.A1(n_1937),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1862),
.Y(n_2224)
);

INVx8_ASAP7_75t_L g2225 ( 
.A(n_1859),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1862),
.Y(n_2226)
);

INVxp67_ASAP7_75t_L g2227 ( 
.A(n_2004),
.Y(n_2227)
);

BUFx6f_ASAP7_75t_L g2228 ( 
.A(n_1790),
.Y(n_2228)
);

INVx5_ASAP7_75t_L g2229 ( 
.A(n_1790),
.Y(n_2229)
);

AOI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_1928),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2008),
.Y(n_2231)
);

INVxp67_ASAP7_75t_L g2232 ( 
.A(n_2010),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_L g2233 ( 
.A(n_1767),
.B(n_733),
.Y(n_2233)
);

O2A1O1Ixp33_ASAP7_75t_L g2234 ( 
.A1(n_1830),
.A2(n_128),
.B(n_125),
.C(n_126),
.Y(n_2234)
);

BUFx2_ASAP7_75t_L g2235 ( 
.A(n_1937),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_1884),
.B(n_129),
.Y(n_2236)
);

O2A1O1Ixp33_ASAP7_75t_L g2237 ( 
.A1(n_1835),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_2237)
);

OAI22x1_ASAP7_75t_L g2238 ( 
.A1(n_1885),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_2238)
);

BUFx8_ASAP7_75t_L g2239 ( 
.A(n_1815),
.Y(n_2239)
);

A2O1A1Ixp33_ASAP7_75t_L g2240 ( 
.A1(n_1845),
.A2(n_136),
.B(n_134),
.C(n_135),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1880),
.Y(n_2241)
);

AOI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_1846),
.A2(n_135),
.B(n_136),
.Y(n_2242)
);

AOI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_1939),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1970),
.B(n_138),
.Y(n_2244)
);

OR2x6_ASAP7_75t_L g2245 ( 
.A(n_1810),
.B(n_140),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_1850),
.B(n_731),
.Y(n_2246)
);

AOI21xp5_ASAP7_75t_L g2247 ( 
.A1(n_1858),
.A2(n_141),
.B(n_142),
.Y(n_2247)
);

INVx1_ASAP7_75t_SL g2248 ( 
.A(n_1884),
.Y(n_2248)
);

CKINVDCx14_ASAP7_75t_R g2249 ( 
.A(n_1929),
.Y(n_2249)
);

OAI22x1_ASAP7_75t_L g2250 ( 
.A1(n_1929),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_2250)
);

O2A1O1Ixp33_ASAP7_75t_L g2251 ( 
.A1(n_1888),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_1790),
.B(n_147),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2013),
.Y(n_2253)
);

A2O1A1Ixp33_ASAP7_75t_L g2254 ( 
.A1(n_1953),
.A2(n_151),
.B(n_149),
.C(n_150),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2014),
.Y(n_2255)
);

AOI21xp5_ASAP7_75t_L g2256 ( 
.A1(n_1927),
.A2(n_155),
.B(n_156),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_L g2257 ( 
.A(n_1934),
.B(n_737),
.Y(n_2257)
);

INVx1_ASAP7_75t_SL g2258 ( 
.A(n_1869),
.Y(n_2258)
);

BUFx12f_ASAP7_75t_L g2259 ( 
.A(n_1929),
.Y(n_2259)
);

INVx4_ASAP7_75t_L g2260 ( 
.A(n_2011),
.Y(n_2260)
);

O2A1O1Ixp33_ASAP7_75t_L g2261 ( 
.A1(n_1985),
.A2(n_163),
.B(n_160),
.C(n_162),
.Y(n_2261)
);

NAND2xp33_ASAP7_75t_R g2262 ( 
.A(n_1978),
.B(n_162),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1945),
.Y(n_2263)
);

NOR3xp33_ASAP7_75t_SL g2264 ( 
.A(n_1759),
.B(n_163),
.C(n_164),
.Y(n_2264)
);

OR2x2_ASAP7_75t_L g2265 ( 
.A(n_1842),
.B(n_164),
.Y(n_2265)
);

BUFx6f_ASAP7_75t_L g2266 ( 
.A(n_2011),
.Y(n_2266)
);

BUFx2_ASAP7_75t_L g2267 ( 
.A(n_1840),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_1857),
.B(n_744),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_1955),
.B(n_165),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_SL g2270 ( 
.A(n_2011),
.B(n_166),
.Y(n_2270)
);

INVx4_ASAP7_75t_L g2271 ( 
.A(n_2000),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1946),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1980),
.Y(n_2273)
);

OAI21x1_ASAP7_75t_L g2274 ( 
.A1(n_2001),
.A2(n_167),
.B(n_168),
.Y(n_2274)
);

BUFx2_ASAP7_75t_L g2275 ( 
.A(n_1854),
.Y(n_2275)
);

NOR2xp33_ASAP7_75t_L g2276 ( 
.A(n_1875),
.B(n_725),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1994),
.B(n_168),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1886),
.B(n_169),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_1836),
.B(n_169),
.Y(n_2279)
);

OAI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_1988),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_2280)
);

OAI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_1899),
.A2(n_173),
.B1(n_170),
.B2(n_171),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_1916),
.Y(n_2282)
);

O2A1O1Ixp33_ASAP7_75t_L g2283 ( 
.A1(n_1983),
.A2(n_175),
.B(n_173),
.C(n_174),
.Y(n_2283)
);

BUFx3_ASAP7_75t_L g2284 ( 
.A(n_1949),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_1951),
.B(n_174),
.Y(n_2285)
);

NOR2xp33_ASAP7_75t_L g2286 ( 
.A(n_1933),
.B(n_740),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_1998),
.B(n_1980),
.Y(n_2287)
);

OAI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_1964),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_1949),
.B(n_179),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1801),
.Y(n_2290)
);

AOI21xp5_ASAP7_75t_L g2291 ( 
.A1(n_1821),
.A2(n_180),
.B(n_181),
.Y(n_2291)
);

OAI22xp5_ASAP7_75t_SL g2292 ( 
.A1(n_1949),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_2292)
);

A2O1A1Ixp33_ASAP7_75t_L g2293 ( 
.A1(n_2007),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_2293)
);

AOI21xp5_ASAP7_75t_L g2294 ( 
.A1(n_1999),
.A2(n_185),
.B(n_186),
.Y(n_2294)
);

INVx3_ASAP7_75t_L g2295 ( 
.A(n_1954),
.Y(n_2295)
);

A2O1A1Ixp33_ASAP7_75t_L g2296 ( 
.A1(n_2023),
.A2(n_188),
.B(n_185),
.C(n_187),
.Y(n_2296)
);

BUFx6f_ASAP7_75t_L g2297 ( 
.A(n_1954),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_1995),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_1856),
.B(n_190),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_1993),
.B(n_191),
.Y(n_2300)
);

INVx2_ASAP7_75t_SL g2301 ( 
.A(n_1752),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_2020),
.B(n_193),
.Y(n_2302)
);

BUFx3_ASAP7_75t_L g2303 ( 
.A(n_1958),
.Y(n_2303)
);

AOI21x1_ASAP7_75t_L g2304 ( 
.A1(n_1984),
.A2(n_1982),
.B(n_1977),
.Y(n_2304)
);

INVx2_ASAP7_75t_SL g2305 ( 
.A(n_2022),
.Y(n_2305)
);

BUFx6f_ASAP7_75t_L g2306 ( 
.A(n_2002),
.Y(n_2306)
);

INVx4_ASAP7_75t_L g2307 ( 
.A(n_1828),
.Y(n_2307)
);

OAI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_1996),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_1804),
.B(n_197),
.Y(n_2309)
);

AOI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_1979),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_2310)
);

A2O1A1Ixp33_ASAP7_75t_L g2311 ( 
.A1(n_1961),
.A2(n_201),
.B(n_199),
.C(n_200),
.Y(n_2311)
);

NOR3xp33_ASAP7_75t_L g2312 ( 
.A(n_1979),
.B(n_200),
.C(n_201),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_1961),
.B(n_202),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1750),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_1912),
.B(n_203),
.Y(n_2315)
);

BUFx6f_ASAP7_75t_L g2316 ( 
.A(n_1852),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_1757),
.B(n_205),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_SL g2318 ( 
.A(n_1757),
.B(n_205),
.Y(n_2318)
);

OAI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_1865),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_1813),
.Y(n_2320)
);

INVxp67_ASAP7_75t_L g2321 ( 
.A(n_1756),
.Y(n_2321)
);

AOI22x1_ASAP7_75t_SL g2322 ( 
.A1(n_1764),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_2322)
);

OAI22xp5_ASAP7_75t_L g2323 ( 
.A1(n_1865),
.A2(n_215),
.B1(n_212),
.B2(n_214),
.Y(n_2323)
);

OAI22xp5_ASAP7_75t_SL g2324 ( 
.A1(n_1825),
.A2(n_215),
.B1(n_212),
.B2(n_214),
.Y(n_2324)
);

OAI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_1865),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_2325)
);

A2O1A1Ixp33_ASAP7_75t_L g2326 ( 
.A1(n_1910),
.A2(n_220),
.B(n_217),
.C(n_219),
.Y(n_2326)
);

INVx3_ASAP7_75t_L g2327 ( 
.A(n_1765),
.Y(n_2327)
);

OAI21xp33_ASAP7_75t_L g2328 ( 
.A1(n_1797),
.A2(n_219),
.B(n_221),
.Y(n_2328)
);

AND2x2_ASAP7_75t_SL g2329 ( 
.A(n_1793),
.B(n_222),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_1808),
.B(n_222),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_1912),
.B(n_223),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1750),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1750),
.Y(n_2333)
);

BUFx2_ASAP7_75t_L g2334 ( 
.A(n_1756),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_1813),
.Y(n_2335)
);

AOI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_2018),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_2336)
);

AND2x4_ASAP7_75t_L g2337 ( 
.A(n_1909),
.B(n_229),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_1797),
.B(n_229),
.Y(n_2338)
);

NAND2xp33_ASAP7_75t_SL g2339 ( 
.A(n_1793),
.B(n_231),
.Y(n_2339)
);

NOR3xp33_ASAP7_75t_SL g2340 ( 
.A(n_1775),
.B(n_231),
.C(n_232),
.Y(n_2340)
);

OAI22xp5_ASAP7_75t_SL g2341 ( 
.A1(n_1825),
.A2(n_236),
.B1(n_233),
.B2(n_234),
.Y(n_2341)
);

OR2x6_ASAP7_75t_L g2342 ( 
.A(n_1774),
.B(n_233),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_R g2343 ( 
.A(n_1764),
.B(n_237),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_L g2344 ( 
.A(n_1808),
.B(n_240),
.Y(n_2344)
);

INVx4_ASAP7_75t_L g2345 ( 
.A(n_1757),
.Y(n_2345)
);

AND2x4_ASAP7_75t_L g2346 ( 
.A(n_1909),
.B(n_241),
.Y(n_2346)
);

A2O1A1Ixp33_ASAP7_75t_L g2347 ( 
.A1(n_1910),
.A2(n_245),
.B(n_242),
.C(n_243),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_1757),
.B(n_246),
.Y(n_2348)
);

OAI21x1_ASAP7_75t_L g2349 ( 
.A1(n_1917),
.A2(n_246),
.B(n_247),
.Y(n_2349)
);

A2O1A1Ixp33_ASAP7_75t_L g2350 ( 
.A1(n_1910),
.A2(n_251),
.B(n_248),
.C(n_249),
.Y(n_2350)
);

AND2x6_ASAP7_75t_L g2351 ( 
.A(n_1793),
.B(n_252),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_SL g2352 ( 
.A(n_1757),
.B(n_252),
.Y(n_2352)
);

OAI21xp5_ASAP7_75t_L g2353 ( 
.A1(n_1910),
.A2(n_253),
.B(n_255),
.Y(n_2353)
);

AND2x4_ASAP7_75t_L g2354 ( 
.A(n_1909),
.B(n_253),
.Y(n_2354)
);

NOR2xp33_ASAP7_75t_L g2355 ( 
.A(n_1808),
.B(n_255),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1750),
.Y(n_2356)
);

A2O1A1Ixp33_ASAP7_75t_L g2357 ( 
.A1(n_1910),
.A2(n_259),
.B(n_257),
.C(n_258),
.Y(n_2357)
);

O2A1O1Ixp33_ASAP7_75t_L g2358 ( 
.A1(n_1913),
.A2(n_260),
.B(n_257),
.C(n_259),
.Y(n_2358)
);

NOR2x1_ASAP7_75t_L g2359 ( 
.A(n_1959),
.B(n_262),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_1813),
.Y(n_2360)
);

INVxp67_ASAP7_75t_SL g2361 ( 
.A(n_1793),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_1757),
.B(n_264),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_1853),
.Y(n_2363)
);

OR2x2_ASAP7_75t_L g2364 ( 
.A(n_1811),
.B(n_264),
.Y(n_2364)
);

A2O1A1Ixp33_ASAP7_75t_L g2365 ( 
.A1(n_1910),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_2365)
);

NOR3xp33_ASAP7_75t_SL g2366 ( 
.A(n_1775),
.B(n_265),
.C(n_266),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_1797),
.B(n_267),
.Y(n_2367)
);

O2A1O1Ixp33_ASAP7_75t_L g2368 ( 
.A1(n_1913),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_2368)
);

AOI22xp5_ASAP7_75t_L g2369 ( 
.A1(n_2018),
.A2(n_272),
.B1(n_268),
.B2(n_269),
.Y(n_2369)
);

OA22x2_ASAP7_75t_L g2370 ( 
.A1(n_1825),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_1912),
.B(n_276),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_1750),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_1912),
.B(n_276),
.Y(n_2373)
);

BUFx3_ASAP7_75t_L g2374 ( 
.A(n_1757),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_R g2375 ( 
.A(n_1764),
.B(n_277),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_1813),
.Y(n_2376)
);

OAI22xp5_ASAP7_75t_L g2377 ( 
.A1(n_1865),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1797),
.B(n_283),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_1813),
.Y(n_2379)
);

OAI22x1_ASAP7_75t_L g2380 ( 
.A1(n_1766),
.A2(n_288),
.B1(n_283),
.B2(n_284),
.Y(n_2380)
);

AOI22xp5_ASAP7_75t_L g2381 ( 
.A1(n_2018),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.Y(n_2381)
);

INVx2_ASAP7_75t_SL g2382 ( 
.A(n_1757),
.Y(n_2382)
);

INVxp67_ASAP7_75t_L g2383 ( 
.A(n_1756),
.Y(n_2383)
);

CKINVDCx5p33_ASAP7_75t_R g2384 ( 
.A(n_1853),
.Y(n_2384)
);

AOI21x1_ASAP7_75t_L g2385 ( 
.A1(n_1911),
.A2(n_291),
.B(n_292),
.Y(n_2385)
);

NOR3xp33_ASAP7_75t_SL g2386 ( 
.A(n_1775),
.B(n_294),
.C(n_295),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_1813),
.Y(n_2387)
);

AO22x1_ASAP7_75t_L g2388 ( 
.A1(n_1832),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_2388)
);

INVxp67_ASAP7_75t_SL g2389 ( 
.A(n_1793),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_1808),
.B(n_300),
.Y(n_2390)
);

AND2x4_ASAP7_75t_L g2391 ( 
.A(n_1909),
.B(n_302),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_1797),
.B(n_303),
.Y(n_2392)
);

BUFx8_ASAP7_75t_L g2393 ( 
.A(n_1774),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_1808),
.B(n_307),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_L g2395 ( 
.A(n_1808),
.B(n_308),
.Y(n_2395)
);

INVx4_ASAP7_75t_L g2396 ( 
.A(n_1757),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_1797),
.B(n_308),
.Y(n_2397)
);

HB1xp67_ASAP7_75t_L g2398 ( 
.A(n_1756),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_1756),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_L g2400 ( 
.A(n_1808),
.B(n_313),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_1912),
.B(n_314),
.Y(n_2401)
);

OAI21xp5_ASAP7_75t_L g2402 ( 
.A1(n_1910),
.A2(n_314),
.B(n_315),
.Y(n_2402)
);

NOR2xp33_ASAP7_75t_L g2403 ( 
.A(n_1808),
.B(n_316),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_1808),
.B(n_316),
.Y(n_2404)
);

OAI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_1865),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_2405)
);

INVx1_ASAP7_75t_SL g2406 ( 
.A(n_1756),
.Y(n_2406)
);

AO21x1_ASAP7_75t_L g2407 ( 
.A1(n_1908),
.A2(n_318),
.B(n_319),
.Y(n_2407)
);

OAI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_1865),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.Y(n_2408)
);

BUFx6f_ASAP7_75t_L g2409 ( 
.A(n_1852),
.Y(n_2409)
);

OAI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_1865),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_1797),
.B(n_323),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_1750),
.Y(n_2412)
);

AOI21x1_ASAP7_75t_L g2413 ( 
.A1(n_1911),
.A2(n_327),
.B(n_328),
.Y(n_2413)
);

NOR3xp33_ASAP7_75t_L g2414 ( 
.A(n_1863),
.B(n_330),
.C(n_331),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_1750),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1750),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_1797),
.B(n_332),
.Y(n_2417)
);

NAND2x1p5_ASAP7_75t_L g2418 ( 
.A(n_1757),
.B(n_333),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_1797),
.B(n_333),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1750),
.Y(n_2420)
);

AO32x1_ASAP7_75t_L g2421 ( 
.A1(n_1917),
.A2(n_336),
.A3(n_334),
.B1(n_335),
.B2(n_337),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_L g2422 ( 
.A(n_1808),
.B(n_335),
.Y(n_2422)
);

NAND3xp33_ASAP7_75t_SL g2423 ( 
.A(n_1831),
.B(n_337),
.C(n_338),
.Y(n_2423)
);

HB1xp67_ASAP7_75t_L g2424 ( 
.A(n_1756),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_1813),
.Y(n_2425)
);

INVxp67_ASAP7_75t_L g2426 ( 
.A(n_1756),
.Y(n_2426)
);

INVx5_ASAP7_75t_L g2427 ( 
.A(n_2005),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_1797),
.B(n_339),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_L g2429 ( 
.A(n_1808),
.B(n_339),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_1808),
.B(n_340),
.Y(n_2430)
);

NOR2xp33_ASAP7_75t_L g2431 ( 
.A(n_1808),
.B(n_341),
.Y(n_2431)
);

XOR2xp5_ASAP7_75t_L g2432 ( 
.A(n_1825),
.B(n_343),
.Y(n_2432)
);

CKINVDCx11_ASAP7_75t_R g2433 ( 
.A(n_1774),
.Y(n_2433)
);

OAI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_1865),
.A2(n_346),
.B1(n_343),
.B2(n_344),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_1813),
.Y(n_2435)
);

AO31x2_ASAP7_75t_L g2436 ( 
.A1(n_1917),
.A2(n_347),
.A3(n_344),
.B(n_346),
.Y(n_2436)
);

AO32x2_ASAP7_75t_L g2437 ( 
.A1(n_1890),
.A2(n_350),
.A3(n_348),
.B1(n_349),
.B2(n_351),
.Y(n_2437)
);

NOR3xp33_ASAP7_75t_SL g2438 ( 
.A(n_1775),
.B(n_351),
.C(n_352),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_1797),
.B(n_353),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_1750),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_1813),
.Y(n_2441)
);

AOI21xp5_ASAP7_75t_L g2442 ( 
.A1(n_1944),
.A2(n_356),
.B(n_358),
.Y(n_2442)
);

AOI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_1944),
.A2(n_358),
.B(n_359),
.Y(n_2443)
);

OAI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_1865),
.A2(n_363),
.B1(n_360),
.B2(n_361),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_SL g2445 ( 
.A(n_1780),
.B(n_360),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_1813),
.Y(n_2446)
);

NOR2xp33_ASAP7_75t_L g2447 ( 
.A(n_1808),
.B(n_364),
.Y(n_2447)
);

OA21x2_ASAP7_75t_L g2448 ( 
.A1(n_2349),
.A2(n_2274),
.B(n_2353),
.Y(n_2448)
);

INVx3_ASAP7_75t_L g2449 ( 
.A(n_2260),
.Y(n_2449)
);

BUFx4_ASAP7_75t_SL g2450 ( 
.A(n_2082),
.Y(n_2450)
);

INVx5_ASAP7_75t_SL g2451 ( 
.A(n_2342),
.Y(n_2451)
);

BUFx2_ASAP7_75t_L g2452 ( 
.A(n_2239),
.Y(n_2452)
);

INVx3_ASAP7_75t_L g2453 ( 
.A(n_2260),
.Y(n_2453)
);

AOI22x1_ASAP7_75t_L g2454 ( 
.A1(n_2085),
.A2(n_370),
.B1(n_365),
.B2(n_369),
.Y(n_2454)
);

INVx3_ASAP7_75t_L g2455 ( 
.A(n_2229),
.Y(n_2455)
);

AND2x4_ASAP7_75t_L g2456 ( 
.A(n_2058),
.B(n_369),
.Y(n_2456)
);

BUFx12f_ASAP7_75t_L g2457 ( 
.A(n_2086),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2329),
.B(n_370),
.Y(n_2458)
);

BUFx2_ASAP7_75t_R g2459 ( 
.A(n_2363),
.Y(n_2459)
);

AO21x2_ASAP7_75t_L g2460 ( 
.A1(n_2402),
.A2(n_371),
.B(n_372),
.Y(n_2460)
);

INVx4_ASAP7_75t_L g2461 ( 
.A(n_2225),
.Y(n_2461)
);

BUFx4_ASAP7_75t_SL g2462 ( 
.A(n_2384),
.Y(n_2462)
);

OAI22xp5_ASAP7_75t_L g2463 ( 
.A1(n_2178),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2112),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2117),
.Y(n_2465)
);

HB1xp67_ASAP7_75t_L g2466 ( 
.A(n_2098),
.Y(n_2466)
);

OR2x2_ASAP7_75t_L g2467 ( 
.A(n_2406),
.B(n_375),
.Y(n_2467)
);

INVx3_ASAP7_75t_L g2468 ( 
.A(n_2229),
.Y(n_2468)
);

OA21x2_ASAP7_75t_L g2469 ( 
.A1(n_2407),
.A2(n_376),
.B(n_377),
.Y(n_2469)
);

OR2x2_ASAP7_75t_L g2470 ( 
.A(n_2051),
.B(n_376),
.Y(n_2470)
);

CKINVDCx20_ASAP7_75t_R g2471 ( 
.A(n_2125),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2231),
.B(n_377),
.Y(n_2472)
);

CKINVDCx20_ASAP7_75t_R g2473 ( 
.A(n_2056),
.Y(n_2473)
);

INVx1_ASAP7_75t_SL g2474 ( 
.A(n_2334),
.Y(n_2474)
);

INVx1_ASAP7_75t_SL g2475 ( 
.A(n_2399),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2039),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2320),
.Y(n_2477)
);

BUFx3_ASAP7_75t_L g2478 ( 
.A(n_2225),
.Y(n_2478)
);

OAI21xp5_ASAP7_75t_L g2479 ( 
.A1(n_2089),
.A2(n_379),
.B(n_380),
.Y(n_2479)
);

INVx3_ASAP7_75t_L g2480 ( 
.A(n_2229),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2335),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_SL g2482 ( 
.A(n_2359),
.B(n_2201),
.Y(n_2482)
);

BUFx2_ASAP7_75t_R g2483 ( 
.A(n_2215),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_L g2484 ( 
.A(n_2031),
.B(n_2211),
.Y(n_2484)
);

NAND2x1p5_ASAP7_75t_L g2485 ( 
.A(n_2074),
.B(n_381),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2071),
.Y(n_2486)
);

OAI21xp5_ASAP7_75t_L g2487 ( 
.A1(n_2163),
.A2(n_382),
.B(n_383),
.Y(n_2487)
);

NAND2x1p5_ASAP7_75t_L g2488 ( 
.A(n_2074),
.B(n_382),
.Y(n_2488)
);

INVx5_ASAP7_75t_L g2489 ( 
.A(n_2158),
.Y(n_2489)
);

AOI21xp5_ASAP7_75t_L g2490 ( 
.A1(n_2131),
.A2(n_383),
.B(n_384),
.Y(n_2490)
);

AO21x2_ASAP7_75t_L g2491 ( 
.A1(n_2385),
.A2(n_384),
.B(n_386),
.Y(n_2491)
);

INVx2_ASAP7_75t_SL g2492 ( 
.A(n_2056),
.Y(n_2492)
);

CKINVDCx16_ASAP7_75t_R g2493 ( 
.A(n_2065),
.Y(n_2493)
);

AO21x2_ASAP7_75t_L g2494 ( 
.A1(n_2413),
.A2(n_386),
.B(n_387),
.Y(n_2494)
);

INVx2_ASAP7_75t_SL g2495 ( 
.A(n_2393),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2360),
.Y(n_2496)
);

AOI22x1_ASAP7_75t_L g2497 ( 
.A1(n_2050),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_2497)
);

CKINVDCx5p33_ASAP7_75t_R g2498 ( 
.A(n_2033),
.Y(n_2498)
);

INVx5_ASAP7_75t_L g2499 ( 
.A(n_2158),
.Y(n_2499)
);

NOR2xp33_ASAP7_75t_L g2500 ( 
.A(n_2197),
.B(n_388),
.Y(n_2500)
);

AOI22xp5_ASAP7_75t_L g2501 ( 
.A1(n_2178),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.Y(n_2501)
);

NAND2x1p5_ASAP7_75t_L g2502 ( 
.A(n_2179),
.B(n_391),
.Y(n_2502)
);

BUFx12f_ASAP7_75t_L g2503 ( 
.A(n_2063),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2376),
.Y(n_2504)
);

OAI21x1_ASAP7_75t_SL g2505 ( 
.A1(n_2192),
.A2(n_394),
.B(n_395),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2379),
.Y(n_2506)
);

OAI21x1_ASAP7_75t_L g2507 ( 
.A1(n_2304),
.A2(n_396),
.B(n_399),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2387),
.Y(n_2508)
);

AOI22x1_ASAP7_75t_L g2509 ( 
.A1(n_2109),
.A2(n_402),
.B1(n_399),
.B2(n_401),
.Y(n_2509)
);

NAND2xp33_ASAP7_75t_L g2510 ( 
.A(n_2158),
.B(n_402),
.Y(n_2510)
);

NOR2x1_ASAP7_75t_L g2511 ( 
.A(n_2345),
.B(n_403),
.Y(n_2511)
);

INVx1_ASAP7_75t_SL g2512 ( 
.A(n_2258),
.Y(n_2512)
);

BUFx6f_ASAP7_75t_L g2513 ( 
.A(n_2053),
.Y(n_2513)
);

BUFx4f_ASAP7_75t_L g2514 ( 
.A(n_2342),
.Y(n_2514)
);

NAND2x1p5_ASAP7_75t_L g2515 ( 
.A(n_2179),
.B(n_404),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2425),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2253),
.B(n_405),
.Y(n_2517)
);

INVx4_ASAP7_75t_L g2518 ( 
.A(n_2225),
.Y(n_2518)
);

OAI21x1_ASAP7_75t_L g2519 ( 
.A1(n_2295),
.A2(n_406),
.B(n_408),
.Y(n_2519)
);

NAND2x1p5_ASAP7_75t_L g2520 ( 
.A(n_2179),
.B(n_406),
.Y(n_2520)
);

OAI21x1_ASAP7_75t_L g2521 ( 
.A1(n_2295),
.A2(n_408),
.B(n_409),
.Y(n_2521)
);

BUFx3_ASAP7_75t_L g2522 ( 
.A(n_2239),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2435),
.Y(n_2523)
);

AND2x4_ASAP7_75t_L g2524 ( 
.A(n_2058),
.B(n_409),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2441),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2446),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2053),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2034),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2314),
.Y(n_2529)
);

BUFx3_ASAP7_75t_L g2530 ( 
.A(n_2374),
.Y(n_2530)
);

OA21x2_ASAP7_75t_L g2531 ( 
.A1(n_2328),
.A2(n_410),
.B(n_411),
.Y(n_2531)
);

BUFx2_ASAP7_75t_R g2532 ( 
.A(n_2216),
.Y(n_2532)
);

AO21x2_ASAP7_75t_L g2533 ( 
.A1(n_2137),
.A2(n_2201),
.B(n_2166),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2332),
.Y(n_2534)
);

OR2x6_ASAP7_75t_L g2535 ( 
.A(n_2192),
.B(n_412),
.Y(n_2535)
);

BUFx12f_ASAP7_75t_L g2536 ( 
.A(n_2433),
.Y(n_2536)
);

INVx3_ASAP7_75t_L g2537 ( 
.A(n_2345),
.Y(n_2537)
);

CKINVDCx6p67_ASAP7_75t_R g2538 ( 
.A(n_2095),
.Y(n_2538)
);

INVx1_ASAP7_75t_SL g2539 ( 
.A(n_2061),
.Y(n_2539)
);

INVxp67_ASAP7_75t_L g2540 ( 
.A(n_2127),
.Y(n_2540)
);

AO21x2_ASAP7_75t_L g2541 ( 
.A1(n_2180),
.A2(n_413),
.B(n_415),
.Y(n_2541)
);

OAI21x1_ASAP7_75t_L g2542 ( 
.A1(n_2072),
.A2(n_416),
.B(n_418),
.Y(n_2542)
);

OAI21x1_ASAP7_75t_L g2543 ( 
.A1(n_2072),
.A2(n_416),
.B(n_418),
.Y(n_2543)
);

INVx2_ASAP7_75t_SL g2544 ( 
.A(n_2393),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2099),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2255),
.B(n_419),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2333),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2356),
.Y(n_2548)
);

BUFx4_ASAP7_75t_SL g2549 ( 
.A(n_2130),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2099),
.Y(n_2550)
);

CKINVDCx11_ASAP7_75t_R g2551 ( 
.A(n_2087),
.Y(n_2551)
);

CKINVDCx20_ASAP7_75t_R g2552 ( 
.A(n_2151),
.Y(n_2552)
);

AOI22x1_ASAP7_75t_L g2553 ( 
.A1(n_2242),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_2553)
);

BUFx3_ASAP7_75t_L g2554 ( 
.A(n_2120),
.Y(n_2554)
);

NAND2x1p5_ASAP7_75t_L g2555 ( 
.A(n_2193),
.B(n_2044),
.Y(n_2555)
);

INVx5_ASAP7_75t_L g2556 ( 
.A(n_2351),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2372),
.Y(n_2557)
);

BUFx4_ASAP7_75t_SL g2558 ( 
.A(n_2130),
.Y(n_2558)
);

BUFx3_ASAP7_75t_L g2559 ( 
.A(n_2228),
.Y(n_2559)
);

BUFx2_ASAP7_75t_L g2560 ( 
.A(n_2028),
.Y(n_2560)
);

CKINVDCx6p67_ASAP7_75t_R g2561 ( 
.A(n_2245),
.Y(n_2561)
);

BUFx2_ASAP7_75t_SL g2562 ( 
.A(n_2044),
.Y(n_2562)
);

INVx6_ASAP7_75t_L g2563 ( 
.A(n_2396),
.Y(n_2563)
);

BUFx8_ASAP7_75t_SL g2564 ( 
.A(n_2075),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_2227),
.B(n_422),
.Y(n_2565)
);

AO21x2_ASAP7_75t_L g2566 ( 
.A1(n_2313),
.A2(n_423),
.B(n_424),
.Y(n_2566)
);

BUFx2_ASAP7_75t_R g2567 ( 
.A(n_2092),
.Y(n_2567)
);

OAI21x1_ASAP7_75t_L g2568 ( 
.A1(n_2359),
.A2(n_423),
.B(n_425),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2135),
.Y(n_2569)
);

BUFx3_ASAP7_75t_L g2570 ( 
.A(n_2228),
.Y(n_2570)
);

AO21x2_ASAP7_75t_L g2571 ( 
.A1(n_2052),
.A2(n_425),
.B(n_426),
.Y(n_2571)
);

BUFx3_ASAP7_75t_L g2572 ( 
.A(n_2228),
.Y(n_2572)
);

AOI22x1_ASAP7_75t_L g2573 ( 
.A1(n_2247),
.A2(n_429),
.B1(n_427),
.B2(n_428),
.Y(n_2573)
);

BUFx2_ASAP7_75t_R g2574 ( 
.A(n_2199),
.Y(n_2574)
);

OAI21xp5_ASAP7_75t_L g2575 ( 
.A1(n_2080),
.A2(n_427),
.B(n_428),
.Y(n_2575)
);

INVx1_ASAP7_75t_SL g2576 ( 
.A(n_2217),
.Y(n_2576)
);

BUFx3_ASAP7_75t_L g2577 ( 
.A(n_2266),
.Y(n_2577)
);

BUFx2_ASAP7_75t_L g2578 ( 
.A(n_2398),
.Y(n_2578)
);

NOR2x1_ASAP7_75t_R g2579 ( 
.A(n_2044),
.B(n_429),
.Y(n_2579)
);

AOI22xp5_ASAP7_75t_L g2580 ( 
.A1(n_2047),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.Y(n_2580)
);

BUFx2_ASAP7_75t_SL g2581 ( 
.A(n_2073),
.Y(n_2581)
);

BUFx3_ASAP7_75t_L g2582 ( 
.A(n_2266),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2412),
.Y(n_2583)
);

NAND2x1p5_ASAP7_75t_L g2584 ( 
.A(n_2193),
.B(n_432),
.Y(n_2584)
);

INVx6_ASAP7_75t_L g2585 ( 
.A(n_2396),
.Y(n_2585)
);

HB1xp67_ASAP7_75t_L g2586 ( 
.A(n_2337),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2415),
.Y(n_2587)
);

AO21x2_ASAP7_75t_L g2588 ( 
.A1(n_2326),
.A2(n_434),
.B(n_437),
.Y(n_2588)
);

BUFx12f_ASAP7_75t_L g2589 ( 
.A(n_2259),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2169),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2138),
.B(n_437),
.Y(n_2591)
);

AO21x2_ASAP7_75t_L g2592 ( 
.A1(n_2347),
.A2(n_438),
.B(n_439),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2316),
.Y(n_2593)
);

BUFx2_ASAP7_75t_L g2594 ( 
.A(n_2424),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2416),
.Y(n_2595)
);

BUFx4_ASAP7_75t_SL g2596 ( 
.A(n_2245),
.Y(n_2596)
);

INVx1_ASAP7_75t_SL g2597 ( 
.A(n_2248),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2420),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2316),
.Y(n_2599)
);

INVx4_ASAP7_75t_L g2600 ( 
.A(n_2073),
.Y(n_2600)
);

BUFx2_ASAP7_75t_L g2601 ( 
.A(n_2321),
.Y(n_2601)
);

AOI22x1_ASAP7_75t_L g2602 ( 
.A1(n_2256),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2440),
.Y(n_2603)
);

OAI21x1_ASAP7_75t_L g2604 ( 
.A1(n_2183),
.A2(n_2187),
.B(n_2185),
.Y(n_2604)
);

OAI21x1_ASAP7_75t_L g2605 ( 
.A1(n_2205),
.A2(n_443),
.B(n_445),
.Y(n_2605)
);

BUFx3_ASAP7_75t_L g2606 ( 
.A(n_2111),
.Y(n_2606)
);

AOI22x1_ASAP7_75t_L g2607 ( 
.A1(n_2222),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.Y(n_2607)
);

INVx4_ASAP7_75t_L g2608 ( 
.A(n_2073),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2168),
.B(n_447),
.Y(n_2609)
);

BUFx3_ASAP7_75t_L g2610 ( 
.A(n_2036),
.Y(n_2610)
);

HB1xp67_ASAP7_75t_L g2611 ( 
.A(n_2337),
.Y(n_2611)
);

AND2x4_ASAP7_75t_L g2612 ( 
.A(n_2083),
.B(n_448),
.Y(n_2612)
);

OAI21x1_ASAP7_75t_L g2613 ( 
.A1(n_2055),
.A2(n_450),
.B(n_451),
.Y(n_2613)
);

NAND2x1p5_ASAP7_75t_L g2614 ( 
.A(n_2193),
.B(n_450),
.Y(n_2614)
);

INVx1_ASAP7_75t_SL g2615 ( 
.A(n_2159),
.Y(n_2615)
);

BUFx3_ASAP7_75t_L g2616 ( 
.A(n_2382),
.Y(n_2616)
);

INVx5_ASAP7_75t_SL g2617 ( 
.A(n_2075),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2064),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_2081),
.Y(n_2619)
);

AO21x2_ASAP7_75t_L g2620 ( 
.A1(n_2350),
.A2(n_453),
.B(n_454),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_L g2621 ( 
.A(n_2232),
.B(n_454),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2067),
.Y(n_2622)
);

AO21x2_ASAP7_75t_L g2623 ( 
.A1(n_2357),
.A2(n_455),
.B(n_456),
.Y(n_2623)
);

INVxp67_ASAP7_75t_SL g2624 ( 
.A(n_2346),
.Y(n_2624)
);

AO21x2_ASAP7_75t_L g2625 ( 
.A1(n_2365),
.A2(n_457),
.B(n_458),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2315),
.B(n_458),
.Y(n_2626)
);

NAND2x1p5_ASAP7_75t_L g2627 ( 
.A(n_2083),
.B(n_460),
.Y(n_2627)
);

HB1xp67_ASAP7_75t_L g2628 ( 
.A(n_2346),
.Y(n_2628)
);

CKINVDCx16_ASAP7_75t_R g2629 ( 
.A(n_2153),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2177),
.B(n_461),
.Y(n_2630)
);

INVx4_ASAP7_75t_L g2631 ( 
.A(n_2083),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_2331),
.B(n_461),
.Y(n_2632)
);

BUFx12f_ASAP7_75t_L g2633 ( 
.A(n_2157),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2068),
.Y(n_2634)
);

BUFx3_ASAP7_75t_L g2635 ( 
.A(n_2306),
.Y(n_2635)
);

OAI21xp5_ASAP7_75t_L g2636 ( 
.A1(n_2041),
.A2(n_462),
.B(n_463),
.Y(n_2636)
);

OAI21xp5_ASAP7_75t_L g2637 ( 
.A1(n_2042),
.A2(n_464),
.B(n_465),
.Y(n_2637)
);

AND2x4_ASAP7_75t_L g2638 ( 
.A(n_2427),
.B(n_464),
.Y(n_2638)
);

INVx1_ASAP7_75t_SL g2639 ( 
.A(n_2184),
.Y(n_2639)
);

AND2x4_ASAP7_75t_L g2640 ( 
.A(n_2427),
.B(n_467),
.Y(n_2640)
);

INVx6_ASAP7_75t_L g2641 ( 
.A(n_2306),
.Y(n_2641)
);

OAI21x1_ASAP7_75t_SL g2642 ( 
.A1(n_2307),
.A2(n_469),
.B(n_470),
.Y(n_2642)
);

BUFx8_ASAP7_75t_SL g2643 ( 
.A(n_2235),
.Y(n_2643)
);

BUFx3_ASAP7_75t_L g2644 ( 
.A(n_2306),
.Y(n_2644)
);

AO21x2_ASAP7_75t_L g2645 ( 
.A1(n_2043),
.A2(n_471),
.B(n_472),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2069),
.Y(n_2646)
);

AND2x4_ASAP7_75t_L g2647 ( 
.A(n_2427),
.B(n_471),
.Y(n_2647)
);

INVx6_ASAP7_75t_L g2648 ( 
.A(n_2271),
.Y(n_2648)
);

BUFx2_ASAP7_75t_L g2649 ( 
.A(n_2383),
.Y(n_2649)
);

INVx2_ASAP7_75t_SL g2650 ( 
.A(n_2148),
.Y(n_2650)
);

OAI21xp5_ASAP7_75t_L g2651 ( 
.A1(n_2030),
.A2(n_2367),
.B(n_2338),
.Y(n_2651)
);

INVx6_ASAP7_75t_SL g2652 ( 
.A(n_2148),
.Y(n_2652)
);

HB1xp67_ASAP7_75t_L g2653 ( 
.A(n_2354),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2090),
.Y(n_2654)
);

OAI21x1_ASAP7_75t_L g2655 ( 
.A1(n_2442),
.A2(n_474),
.B(n_475),
.Y(n_2655)
);

BUFx3_ASAP7_75t_L g2656 ( 
.A(n_2297),
.Y(n_2656)
);

BUFx4f_ASAP7_75t_L g2657 ( 
.A(n_2351),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2097),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2371),
.B(n_474),
.Y(n_2659)
);

BUFx12f_ASAP7_75t_L g2660 ( 
.A(n_2271),
.Y(n_2660)
);

BUFx12f_ASAP7_75t_L g2661 ( 
.A(n_2289),
.Y(n_2661)
);

BUFx2_ASAP7_75t_R g2662 ( 
.A(n_2054),
.Y(n_2662)
);

INVx1_ASAP7_75t_SL g2663 ( 
.A(n_2267),
.Y(n_2663)
);

NAND2x1p5_ASAP7_75t_L g2664 ( 
.A(n_2354),
.B(n_475),
.Y(n_2664)
);

OAI21x1_ASAP7_75t_L g2665 ( 
.A1(n_2443),
.A2(n_476),
.B(n_477),
.Y(n_2665)
);

AOI22x1_ASAP7_75t_L g2666 ( 
.A1(n_2294),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2122),
.Y(n_2667)
);

INVxp67_ASAP7_75t_L g2668 ( 
.A(n_2391),
.Y(n_2668)
);

OAI21x1_ASAP7_75t_SL g2669 ( 
.A1(n_2307),
.A2(n_481),
.B(n_482),
.Y(n_2669)
);

AO21x2_ASAP7_75t_L g2670 ( 
.A1(n_2277),
.A2(n_484),
.B(n_485),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2132),
.Y(n_2671)
);

INVxp67_ASAP7_75t_L g2672 ( 
.A(n_2391),
.Y(n_2672)
);

AOI22x1_ASAP7_75t_L g2673 ( 
.A1(n_2291),
.A2(n_487),
.B1(n_485),
.B2(n_486),
.Y(n_2673)
);

HB1xp67_ASAP7_75t_L g2674 ( 
.A(n_2093),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2409),
.Y(n_2675)
);

NOR2xp67_ASAP7_75t_L g2676 ( 
.A(n_2078),
.B(n_486),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2194),
.B(n_489),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2195),
.B(n_489),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2373),
.B(n_490),
.Y(n_2679)
);

OAI21xp5_ASAP7_75t_L g2680 ( 
.A1(n_2378),
.A2(n_491),
.B(n_492),
.Y(n_2680)
);

HB1xp67_ASAP7_75t_L g2681 ( 
.A(n_2093),
.Y(n_2681)
);

OAI21x1_ASAP7_75t_SL g2682 ( 
.A1(n_2336),
.A2(n_491),
.B(n_493),
.Y(n_2682)
);

INVx8_ASAP7_75t_L g2683 ( 
.A(n_2351),
.Y(n_2683)
);

AO21x1_ASAP7_75t_L g2684 ( 
.A1(n_2339),
.A2(n_493),
.B(n_494),
.Y(n_2684)
);

NAND2x1p5_ASAP7_75t_L g2685 ( 
.A(n_2409),
.B(n_494),
.Y(n_2685)
);

AO21x2_ASAP7_75t_L g2686 ( 
.A1(n_2293),
.A2(n_495),
.B(n_496),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2290),
.B(n_497),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2060),
.B(n_497),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2155),
.Y(n_2689)
);

BUFx8_ASAP7_75t_L g2690 ( 
.A(n_2289),
.Y(n_2690)
);

INVx5_ASAP7_75t_L g2691 ( 
.A(n_2351),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2218),
.Y(n_2692)
);

AO21x2_ASAP7_75t_L g2693 ( 
.A1(n_2161),
.A2(n_498),
.B(n_500),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2401),
.B(n_500),
.Y(n_2694)
);

CKINVDCx11_ASAP7_75t_R g2695 ( 
.A(n_2115),
.Y(n_2695)
);

BUFx2_ASAP7_75t_L g2696 ( 
.A(n_2426),
.Y(n_2696)
);

CKINVDCx14_ASAP7_75t_R g2697 ( 
.A(n_2110),
.Y(n_2697)
);

OAI21xp5_ASAP7_75t_L g2698 ( 
.A1(n_2392),
.A2(n_501),
.B(n_503),
.Y(n_2698)
);

INVx3_ASAP7_75t_L g2699 ( 
.A(n_2035),
.Y(n_2699)
);

BUFx2_ASAP7_75t_SL g2700 ( 
.A(n_2108),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_2343),
.Y(n_2701)
);

AO21x2_ASAP7_75t_L g2702 ( 
.A1(n_2167),
.A2(n_501),
.B(n_503),
.Y(n_2702)
);

OAI21x1_ASAP7_75t_L g2703 ( 
.A1(n_2126),
.A2(n_504),
.B(n_507),
.Y(n_2703)
);

AND2x6_ASAP7_75t_L g2704 ( 
.A(n_2108),
.B(n_504),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2220),
.B(n_508),
.Y(n_2705)
);

INVx1_ASAP7_75t_SL g2706 ( 
.A(n_2102),
.Y(n_2706)
);

BUFx2_ASAP7_75t_SL g2707 ( 
.A(n_2284),
.Y(n_2707)
);

OA21x2_ASAP7_75t_L g2708 ( 
.A1(n_2200),
.A2(n_508),
.B(n_509),
.Y(n_2708)
);

OAI21xp5_ASAP7_75t_L g2709 ( 
.A1(n_2397),
.A2(n_509),
.B(n_510),
.Y(n_2709)
);

AO21x2_ASAP7_75t_L g2710 ( 
.A1(n_2176),
.A2(n_510),
.B(n_511),
.Y(n_2710)
);

BUFx2_ASAP7_75t_L g2711 ( 
.A(n_2119),
.Y(n_2711)
);

NAND2x1p5_ASAP7_75t_L g2712 ( 
.A(n_2160),
.B(n_512),
.Y(n_2712)
);

OAI21xp5_ASAP7_75t_L g2713 ( 
.A1(n_2411),
.A2(n_512),
.B(n_515),
.Y(n_2713)
);

OAI21x1_ASAP7_75t_L g2714 ( 
.A1(n_2160),
.A2(n_515),
.B(n_516),
.Y(n_2714)
);

AOI22x1_ASAP7_75t_L g2715 ( 
.A1(n_2188),
.A2(n_519),
.B1(n_517),
.B2(n_518),
.Y(n_2715)
);

AND2x2_ASAP7_75t_SL g2716 ( 
.A(n_2142),
.B(n_743),
.Y(n_2716)
);

BUFx6f_ASAP7_75t_L g2717 ( 
.A(n_2303),
.Y(n_2717)
);

BUFx3_ASAP7_75t_L g2718 ( 
.A(n_2170),
.Y(n_2718)
);

OAI21xp5_ASAP7_75t_L g2719 ( 
.A1(n_2417),
.A2(n_518),
.B(n_520),
.Y(n_2719)
);

BUFx2_ASAP7_75t_L g2720 ( 
.A(n_2249),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_2375),
.Y(n_2721)
);

AO21x2_ASAP7_75t_L g2722 ( 
.A1(n_2240),
.A2(n_520),
.B(n_521),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2263),
.Y(n_2723)
);

NAND2x1p5_ASAP7_75t_L g2724 ( 
.A(n_2207),
.B(n_522),
.Y(n_2724)
);

INVx4_ASAP7_75t_L g2725 ( 
.A(n_2418),
.Y(n_2725)
);

AO21x2_ASAP7_75t_L g2726 ( 
.A1(n_2254),
.A2(n_523),
.B(n_524),
.Y(n_2726)
);

INVx3_ASAP7_75t_L g2727 ( 
.A(n_2327),
.Y(n_2727)
);

HB1xp67_ASAP7_75t_L g2728 ( 
.A(n_2273),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2272),
.Y(n_2729)
);

INVx6_ASAP7_75t_L g2730 ( 
.A(n_2302),
.Y(n_2730)
);

INVx3_ASAP7_75t_L g2731 ( 
.A(n_2327),
.Y(n_2731)
);

OAI21x1_ASAP7_75t_L g2732 ( 
.A1(n_2236),
.A2(n_526),
.B(n_528),
.Y(n_2732)
);

BUFx2_ASAP7_75t_R g2733 ( 
.A(n_2054),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2146),
.Y(n_2734)
);

BUFx12f_ASAP7_75t_L g2735 ( 
.A(n_2209),
.Y(n_2735)
);

AOI22x1_ASAP7_75t_L g2736 ( 
.A1(n_2191),
.A2(n_530),
.B1(n_526),
.B2(n_529),
.Y(n_2736)
);

INVxp67_ASAP7_75t_SL g2737 ( 
.A(n_2336),
.Y(n_2737)
);

CKINVDCx20_ASAP7_75t_R g2738 ( 
.A(n_2154),
.Y(n_2738)
);

HB1xp67_ASAP7_75t_L g2739 ( 
.A(n_2214),
.Y(n_2739)
);

OR2x2_ASAP7_75t_L g2740 ( 
.A(n_2079),
.B(n_530),
.Y(n_2740)
);

BUFx2_ASAP7_75t_L g2741 ( 
.A(n_2275),
.Y(n_2741)
);

INVxp67_ASAP7_75t_SL g2742 ( 
.A(n_2369),
.Y(n_2742)
);

AOI21xp5_ASAP7_75t_L g2743 ( 
.A1(n_2419),
.A2(n_2439),
.B(n_2428),
.Y(n_2743)
);

BUFx2_ASAP7_75t_L g2744 ( 
.A(n_2136),
.Y(n_2744)
);

BUFx12f_ASAP7_75t_L g2745 ( 
.A(n_2301),
.Y(n_2745)
);

BUFx3_ASAP7_75t_L g2746 ( 
.A(n_2189),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_SL g2747 ( 
.A1(n_2152),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.Y(n_2747)
);

OAI21xp5_ASAP7_75t_L g2748 ( 
.A1(n_2032),
.A2(n_531),
.B(n_534),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2147),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2150),
.Y(n_2750)
);

INVx3_ASAP7_75t_L g2751 ( 
.A(n_2196),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2282),
.B(n_535),
.Y(n_2752)
);

HB1xp67_ASAP7_75t_L g2753 ( 
.A(n_2202),
.Y(n_2753)
);

AO21x2_ASAP7_75t_L g2754 ( 
.A1(n_2296),
.A2(n_535),
.B(n_537),
.Y(n_2754)
);

HB1xp67_ASAP7_75t_L g2755 ( 
.A(n_2206),
.Y(n_2755)
);

INVxp67_ASAP7_75t_L g2756 ( 
.A(n_2257),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2208),
.Y(n_2757)
);

OAI21xp5_ASAP7_75t_L g2758 ( 
.A1(n_2156),
.A2(n_537),
.B(n_539),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_L g2759 ( 
.A(n_2287),
.B(n_539),
.Y(n_2759)
);

OAI21x1_ASAP7_75t_L g2760 ( 
.A1(n_2317),
.A2(n_540),
.B(n_541),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2057),
.B(n_2116),
.Y(n_2761)
);

BUFx3_ASAP7_75t_L g2762 ( 
.A(n_2241),
.Y(n_2762)
);

CKINVDCx20_ASAP7_75t_R g2763 ( 
.A(n_2062),
.Y(n_2763)
);

AOI22xp5_ASAP7_75t_L g2764 ( 
.A1(n_2077),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_2764)
);

AND2x6_ASAP7_75t_L g2765 ( 
.A(n_2302),
.B(n_543),
.Y(n_2765)
);

INVx4_ASAP7_75t_L g2766 ( 
.A(n_2152),
.Y(n_2766)
);

NAND2x1p5_ASAP7_75t_L g2767 ( 
.A(n_2029),
.B(n_543),
.Y(n_2767)
);

OAI21x1_ASAP7_75t_SL g2768 ( 
.A1(n_2369),
.A2(n_2381),
.B(n_2310),
.Y(n_2768)
);

NAND2xp33_ASAP7_75t_L g2769 ( 
.A(n_2264),
.B(n_544),
.Y(n_2769)
);

INVx3_ASAP7_75t_L g2770 ( 
.A(n_2298),
.Y(n_2770)
);

AO21x2_ASAP7_75t_L g2771 ( 
.A1(n_2088),
.A2(n_544),
.B(n_545),
.Y(n_2771)
);

INVx4_ASAP7_75t_L g2772 ( 
.A(n_2364),
.Y(n_2772)
);

CKINVDCx20_ASAP7_75t_R g2773 ( 
.A(n_2223),
.Y(n_2773)
);

BUFx2_ASAP7_75t_SL g2774 ( 
.A(n_2038),
.Y(n_2774)
);

AOI22x1_ASAP7_75t_L g2775 ( 
.A1(n_2238),
.A2(n_549),
.B1(n_546),
.B2(n_548),
.Y(n_2775)
);

OAI21x1_ASAP7_75t_L g2776 ( 
.A1(n_2318),
.A2(n_546),
.B(n_548),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2027),
.B(n_550),
.Y(n_2777)
);

OR2x2_ASAP7_75t_L g2778 ( 
.A(n_2027),
.B(n_550),
.Y(n_2778)
);

NAND2x1p5_ASAP7_75t_L g2779 ( 
.A(n_2348),
.B(n_551),
.Y(n_2779)
);

AND2x4_ASAP7_75t_L g2780 ( 
.A(n_2279),
.B(n_551),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2124),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2436),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2128),
.Y(n_2783)
);

INVx3_ASAP7_75t_L g2784 ( 
.A(n_2172),
.Y(n_2784)
);

NAND2x1p5_ASAP7_75t_L g2785 ( 
.A(n_2352),
.B(n_552),
.Y(n_2785)
);

AND2x4_ASAP7_75t_L g2786 ( 
.A(n_2305),
.B(n_552),
.Y(n_2786)
);

BUFx3_ASAP7_75t_L g2787 ( 
.A(n_2213),
.Y(n_2787)
);

BUFx6f_ASAP7_75t_L g2788 ( 
.A(n_2362),
.Y(n_2788)
);

HB1xp67_ASAP7_75t_L g2789 ( 
.A(n_2224),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2269),
.B(n_553),
.Y(n_2790)
);

BUFx2_ASAP7_75t_L g2791 ( 
.A(n_2212),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2246),
.B(n_2162),
.Y(n_2792)
);

AND2x4_ASAP7_75t_L g2793 ( 
.A(n_2226),
.B(n_553),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2381),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2437),
.Y(n_2795)
);

AO21x2_ASAP7_75t_L g2796 ( 
.A1(n_2204),
.A2(n_555),
.B(n_556),
.Y(n_2796)
);

BUFx3_ASAP7_75t_L g2797 ( 
.A(n_2106),
.Y(n_2797)
);

AO21x2_ASAP7_75t_L g2798 ( 
.A1(n_2219),
.A2(n_556),
.B(n_557),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2101),
.B(n_558),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2244),
.Y(n_2800)
);

INVx4_ASAP7_75t_L g2801 ( 
.A(n_2265),
.Y(n_2801)
);

INVx1_ASAP7_75t_SL g2802 ( 
.A(n_2134),
.Y(n_2802)
);

INVx2_ASAP7_75t_SL g2803 ( 
.A(n_2143),
.Y(n_2803)
);

OAI21xp5_ASAP7_75t_L g2804 ( 
.A1(n_2045),
.A2(n_559),
.B(n_560),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2186),
.B(n_560),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2310),
.Y(n_2806)
);

OAI21x1_ASAP7_75t_L g2807 ( 
.A1(n_2066),
.A2(n_561),
.B(n_562),
.Y(n_2807)
);

AOI22xp33_ASAP7_75t_L g2808 ( 
.A1(n_2414),
.A2(n_561),
.B1(n_562),
.B2(n_563),
.Y(n_2808)
);

INVx1_ASAP7_75t_SL g2809 ( 
.A(n_2103),
.Y(n_2809)
);

BUFx12f_ASAP7_75t_L g2810 ( 
.A(n_2445),
.Y(n_2810)
);

BUFx2_ASAP7_75t_L g2811 ( 
.A(n_2107),
.Y(n_2811)
);

CKINVDCx5p33_ASAP7_75t_R g2812 ( 
.A(n_2262),
.Y(n_2812)
);

HB1xp67_ASAP7_75t_L g2813 ( 
.A(n_2144),
.Y(n_2813)
);

BUFx8_ASAP7_75t_L g2814 ( 
.A(n_2437),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2300),
.B(n_564),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2278),
.Y(n_2816)
);

BUFx3_ASAP7_75t_L g2817 ( 
.A(n_2149),
.Y(n_2817)
);

AO21x2_ASAP7_75t_L g2818 ( 
.A1(n_2311),
.A2(n_565),
.B(n_566),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2437),
.Y(n_2819)
);

AND2x4_ASAP7_75t_L g2820 ( 
.A(n_2361),
.B(n_566),
.Y(n_2820)
);

NAND2x1p5_ASAP7_75t_L g2821 ( 
.A(n_2252),
.B(n_2270),
.Y(n_2821)
);

BUFx3_ASAP7_75t_L g2822 ( 
.A(n_2118),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2285),
.Y(n_2823)
);

AND2x2_ASAP7_75t_L g2824 ( 
.A(n_2040),
.B(n_567),
.Y(n_2824)
);

AO21x2_ASAP7_75t_L g2825 ( 
.A1(n_2070),
.A2(n_567),
.B(n_568),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2141),
.Y(n_2826)
);

AND2x4_ASAP7_75t_L g2827 ( 
.A(n_2389),
.B(n_568),
.Y(n_2827)
);

AND2x2_ASAP7_75t_L g2828 ( 
.A(n_2133),
.B(n_570),
.Y(n_2828)
);

AOI22x1_ASAP7_75t_L g2829 ( 
.A1(n_2250),
.A2(n_571),
.B1(n_572),
.B2(n_573),
.Y(n_2829)
);

NOR2xp33_ASAP7_75t_L g2830 ( 
.A(n_2037),
.B(n_572),
.Y(n_2830)
);

BUFx3_ASAP7_75t_L g2831 ( 
.A(n_2299),
.Y(n_2831)
);

INVx5_ASAP7_75t_L g2832 ( 
.A(n_2292),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2506),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2692),
.Y(n_2834)
);

BUFx2_ASAP7_75t_L g2835 ( 
.A(n_2652),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2723),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2506),
.Y(n_2837)
);

INVx1_ASAP7_75t_SL g2838 ( 
.A(n_2700),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2729),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2508),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2528),
.Y(n_2841)
);

AOI21x1_ASAP7_75t_L g2842 ( 
.A1(n_2482),
.A2(n_2113),
.B(n_2091),
.Y(n_2842)
);

INVx2_ASAP7_75t_SL g2843 ( 
.A(n_2478),
.Y(n_2843)
);

AOI22xp33_ASAP7_75t_L g2844 ( 
.A1(n_2766),
.A2(n_2105),
.B1(n_2123),
.B2(n_2100),
.Y(n_2844)
);

BUFx3_ASAP7_75t_L g2845 ( 
.A(n_2473),
.Y(n_2845)
);

BUFx3_ASAP7_75t_L g2846 ( 
.A(n_2473),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2529),
.Y(n_2847)
);

OAI22xp5_ASAP7_75t_L g2848 ( 
.A1(n_2624),
.A2(n_2141),
.B1(n_2104),
.B2(n_2175),
.Y(n_2848)
);

AOI22xp33_ASAP7_75t_L g2849 ( 
.A1(n_2766),
.A2(n_2484),
.B1(n_2768),
.B2(n_2801),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2508),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2534),
.Y(n_2851)
);

NOR2xp33_ASAP7_75t_SL g2852 ( 
.A(n_2657),
.B(n_2173),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2526),
.Y(n_2853)
);

CKINVDCx11_ASAP7_75t_R g2854 ( 
.A(n_2457),
.Y(n_2854)
);

CKINVDCx20_ASAP7_75t_R g2855 ( 
.A(n_2471),
.Y(n_2855)
);

CKINVDCx11_ASAP7_75t_R g2856 ( 
.A(n_2457),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2526),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2464),
.B(n_2370),
.Y(n_2858)
);

AOI22xp33_ASAP7_75t_SL g2859 ( 
.A1(n_2716),
.A2(n_2322),
.B1(n_2221),
.B2(n_2324),
.Y(n_2859)
);

AOI22xp33_ASAP7_75t_L g2860 ( 
.A1(n_2484),
.A2(n_2312),
.B1(n_2423),
.B2(n_2341),
.Y(n_2860)
);

BUFx12f_ASAP7_75t_L g2861 ( 
.A(n_2503),
.Y(n_2861)
);

INVx5_ASAP7_75t_L g2862 ( 
.A(n_2589),
.Y(n_2862)
);

INVx1_ASAP7_75t_SL g2863 ( 
.A(n_2466),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2465),
.B(n_2432),
.Y(n_2864)
);

BUFx3_ASAP7_75t_L g2865 ( 
.A(n_2589),
.Y(n_2865)
);

BUFx8_ASAP7_75t_SL g2866 ( 
.A(n_2503),
.Y(n_2866)
);

BUFx2_ASAP7_75t_L g2867 ( 
.A(n_2652),
.Y(n_2867)
);

NAND2x1p5_ASAP7_75t_L g2868 ( 
.A(n_2489),
.B(n_2182),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2486),
.Y(n_2869)
);

INVx1_ASAP7_75t_SL g2870 ( 
.A(n_2466),
.Y(n_2870)
);

AOI21x1_ASAP7_75t_L g2871 ( 
.A1(n_2482),
.A2(n_2280),
.B(n_2388),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2486),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2547),
.Y(n_2873)
);

OAI22xp33_ASAP7_75t_SL g2874 ( 
.A1(n_2458),
.A2(n_2281),
.B1(n_2308),
.B2(n_2319),
.Y(n_2874)
);

AND2x2_ASAP7_75t_L g2875 ( 
.A(n_2761),
.B(n_2048),
.Y(n_2875)
);

AOI22xp5_ASAP7_75t_L g2876 ( 
.A1(n_2737),
.A2(n_2210),
.B1(n_2140),
.B2(n_2380),
.Y(n_2876)
);

CKINVDCx6p67_ASAP7_75t_R g2877 ( 
.A(n_2633),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2548),
.Y(n_2878)
);

AOI22xp5_ASAP7_75t_L g2879 ( 
.A1(n_2737),
.A2(n_2288),
.B1(n_2094),
.B2(n_2323),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2557),
.Y(n_2880)
);

INVx3_ASAP7_75t_L g2881 ( 
.A(n_2489),
.Y(n_2881)
);

INVx1_ASAP7_75t_SL g2882 ( 
.A(n_2576),
.Y(n_2882)
);

BUFx6f_ASAP7_75t_L g2883 ( 
.A(n_2478),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2583),
.Y(n_2884)
);

OAI22xp5_ASAP7_75t_L g2885 ( 
.A1(n_2624),
.A2(n_2742),
.B1(n_2657),
.B2(n_2664),
.Y(n_2885)
);

AOI22xp33_ASAP7_75t_L g2886 ( 
.A1(n_2801),
.A2(n_2233),
.B1(n_2276),
.B2(n_2268),
.Y(n_2886)
);

NAND2x1p5_ASAP7_75t_L g2887 ( 
.A(n_2489),
.B(n_2499),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_2772),
.B(n_2181),
.Y(n_2888)
);

AOI22xp5_ASAP7_75t_L g2889 ( 
.A1(n_2742),
.A2(n_2325),
.B1(n_2405),
.B2(n_2377),
.Y(n_2889)
);

BUFx2_ASAP7_75t_L g2890 ( 
.A(n_2690),
.Y(n_2890)
);

AOI22xp33_ASAP7_75t_SL g2891 ( 
.A1(n_2772),
.A2(n_2410),
.B1(n_2434),
.B2(n_2408),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2587),
.Y(n_2892)
);

CKINVDCx11_ASAP7_75t_R g2893 ( 
.A(n_2536),
.Y(n_2893)
);

CKINVDCx20_ASAP7_75t_R g2894 ( 
.A(n_2471),
.Y(n_2894)
);

INVxp67_ASAP7_75t_L g2895 ( 
.A(n_2601),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2595),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2598),
.Y(n_2897)
);

AOI22xp5_ASAP7_75t_L g2898 ( 
.A1(n_2806),
.A2(n_2444),
.B1(n_2330),
.B2(n_2355),
.Y(n_2898)
);

INVxp67_ASAP7_75t_L g2899 ( 
.A(n_2649),
.Y(n_2899)
);

OR2x2_ASAP7_75t_L g2900 ( 
.A(n_2539),
.B(n_2203),
.Y(n_2900)
);

AO21x1_ASAP7_75t_SL g2901 ( 
.A1(n_2586),
.A2(n_2628),
.B(n_2611),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2603),
.Y(n_2902)
);

AOI22xp33_ASAP7_75t_L g2903 ( 
.A1(n_2794),
.A2(n_2286),
.B1(n_2190),
.B2(n_2447),
.Y(n_2903)
);

AO21x2_ASAP7_75t_L g2904 ( 
.A1(n_2782),
.A2(n_2368),
.B(n_2358),
.Y(n_2904)
);

INVx3_ASAP7_75t_L g2905 ( 
.A(n_2489),
.Y(n_2905)
);

INVxp67_ASAP7_75t_L g2906 ( 
.A(n_2696),
.Y(n_2906)
);

BUFx2_ASAP7_75t_L g2907 ( 
.A(n_2690),
.Y(n_2907)
);

INVx4_ASAP7_75t_L g2908 ( 
.A(n_2461),
.Y(n_2908)
);

BUFx3_ASAP7_75t_L g2909 ( 
.A(n_2554),
.Y(n_2909)
);

AOI22xp33_ASAP7_75t_L g2910 ( 
.A1(n_2832),
.A2(n_2390),
.B1(n_2394),
.B2(n_2344),
.Y(n_2910)
);

INVx3_ASAP7_75t_SL g2911 ( 
.A(n_2498),
.Y(n_2911)
);

BUFx12f_ASAP7_75t_L g2912 ( 
.A(n_2498),
.Y(n_2912)
);

NAND2x1p5_ASAP7_75t_L g2913 ( 
.A(n_2499),
.B(n_2198),
.Y(n_2913)
);

BUFx2_ASAP7_75t_L g2914 ( 
.A(n_2661),
.Y(n_2914)
);

HB1xp67_ASAP7_75t_L g2915 ( 
.A(n_2540),
.Y(n_2915)
);

HB1xp67_ASAP7_75t_L g2916 ( 
.A(n_2540),
.Y(n_2916)
);

CKINVDCx11_ASAP7_75t_R g2917 ( 
.A(n_2536),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2618),
.Y(n_2918)
);

CKINVDCx16_ASAP7_75t_R g2919 ( 
.A(n_2493),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2622),
.Y(n_2920)
);

AND2x2_ASAP7_75t_L g2921 ( 
.A(n_2777),
.B(n_2340),
.Y(n_2921)
);

INVx3_ASAP7_75t_L g2922 ( 
.A(n_2499),
.Y(n_2922)
);

AOI22xp33_ASAP7_75t_SL g2923 ( 
.A1(n_2716),
.A2(n_2400),
.B1(n_2403),
.B2(n_2395),
.Y(n_2923)
);

BUFx3_ASAP7_75t_L g2924 ( 
.A(n_2554),
.Y(n_2924)
);

AOI22xp33_ASAP7_75t_L g2925 ( 
.A1(n_2832),
.A2(n_2422),
.B1(n_2429),
.B2(n_2404),
.Y(n_2925)
);

INVxp67_ASAP7_75t_L g2926 ( 
.A(n_2560),
.Y(n_2926)
);

NAND3xp33_ASAP7_75t_SL g2927 ( 
.A(n_2747),
.B(n_2386),
.C(n_2366),
.Y(n_2927)
);

HB1xp67_ASAP7_75t_L g2928 ( 
.A(n_2578),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2556),
.B(n_2438),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2456),
.B(n_2430),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2634),
.Y(n_2931)
);

CKINVDCx11_ASAP7_75t_R g2932 ( 
.A(n_2538),
.Y(n_2932)
);

CKINVDCx6p67_ASAP7_75t_R g2933 ( 
.A(n_2633),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2646),
.Y(n_2934)
);

BUFx3_ASAP7_75t_L g2935 ( 
.A(n_2522),
.Y(n_2935)
);

CKINVDCx11_ASAP7_75t_R g2936 ( 
.A(n_2552),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2654),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2658),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2667),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2671),
.Y(n_2940)
);

INVx1_ASAP7_75t_SL g2941 ( 
.A(n_2597),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2456),
.B(n_2431),
.Y(n_2942)
);

AND2x4_ASAP7_75t_L g2943 ( 
.A(n_2556),
.B(n_2309),
.Y(n_2943)
);

BUFx4f_ASAP7_75t_L g2944 ( 
.A(n_2561),
.Y(n_2944)
);

AO21x1_ASAP7_75t_L g2945 ( 
.A1(n_2458),
.A2(n_2510),
.B(n_2575),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2524),
.B(n_2171),
.Y(n_2946)
);

AOI22xp33_ASAP7_75t_L g2947 ( 
.A1(n_2832),
.A2(n_2174),
.B1(n_2145),
.B2(n_2129),
.Y(n_2947)
);

AOI22xp33_ASAP7_75t_SL g2948 ( 
.A1(n_2617),
.A2(n_2165),
.B1(n_2059),
.B2(n_2046),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2826),
.B(n_2139),
.Y(n_2949)
);

AOI22xp33_ASAP7_75t_L g2950 ( 
.A1(n_2832),
.A2(n_2243),
.B1(n_2230),
.B2(n_2076),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2689),
.Y(n_2951)
);

BUFx6f_ASAP7_75t_L g2952 ( 
.A(n_2513),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2476),
.Y(n_2953)
);

INVx1_ASAP7_75t_SL g2954 ( 
.A(n_2753),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2524),
.B(n_2049),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2477),
.Y(n_2956)
);

BUFx2_ASAP7_75t_L g2957 ( 
.A(n_2661),
.Y(n_2957)
);

AOI22xp33_ASAP7_75t_SL g2958 ( 
.A1(n_2617),
.A2(n_2421),
.B1(n_2164),
.B2(n_2261),
.Y(n_2958)
);

BUFx5_ASAP7_75t_L g2959 ( 
.A(n_2656),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2481),
.Y(n_2960)
);

AOI22xp33_ASAP7_75t_L g2961 ( 
.A1(n_2765),
.A2(n_2084),
.B1(n_2283),
.B2(n_2251),
.Y(n_2961)
);

AOI22xp33_ASAP7_75t_L g2962 ( 
.A1(n_2765),
.A2(n_2237),
.B1(n_2234),
.B2(n_2121),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2496),
.Y(n_2963)
);

AOI22xp5_ASAP7_75t_L g2964 ( 
.A1(n_2765),
.A2(n_2114),
.B1(n_2096),
.B2(n_2421),
.Y(n_2964)
);

CKINVDCx20_ASAP7_75t_R g2965 ( 
.A(n_2552),
.Y(n_2965)
);

INVx2_ASAP7_75t_SL g2966 ( 
.A(n_2461),
.Y(n_2966)
);

OAI22xp5_ASAP7_75t_L g2967 ( 
.A1(n_2664),
.A2(n_573),
.B1(n_574),
.B2(n_575),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2504),
.Y(n_2968)
);

AOI22xp33_ASAP7_75t_SL g2969 ( 
.A1(n_2617),
.A2(n_576),
.B1(n_577),
.B2(n_578),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2516),
.Y(n_2970)
);

INVx2_ASAP7_75t_SL g2971 ( 
.A(n_2518),
.Y(n_2971)
);

HB1xp67_ASAP7_75t_L g2972 ( 
.A(n_2594),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2591),
.B(n_576),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2523),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2525),
.Y(n_2975)
);

BUFx3_ASAP7_75t_L g2976 ( 
.A(n_2522),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2743),
.B(n_577),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2609),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2609),
.Y(n_2979)
);

OA21x2_ASAP7_75t_L g2980 ( 
.A1(n_2795),
.A2(n_2819),
.B(n_2507),
.Y(n_2980)
);

INVx1_ASAP7_75t_SL g2981 ( 
.A(n_2753),
.Y(n_2981)
);

HB1xp67_ASAP7_75t_L g2982 ( 
.A(n_2474),
.Y(n_2982)
);

AOI22xp33_ASAP7_75t_L g2983 ( 
.A1(n_2765),
.A2(n_581),
.B1(n_582),
.B2(n_583),
.Y(n_2983)
);

OAI22xp5_ASAP7_75t_L g2984 ( 
.A1(n_2535),
.A2(n_583),
.B1(n_585),
.B2(n_586),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2630),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2630),
.Y(n_2986)
);

NOR2xp33_ASAP7_75t_L g2987 ( 
.A(n_2773),
.B(n_586),
.Y(n_2987)
);

AOI22xp33_ASAP7_75t_L g2988 ( 
.A1(n_2765),
.A2(n_587),
.B1(n_588),
.B2(n_589),
.Y(n_2988)
);

AOI21xp5_ASAP7_75t_L g2989 ( 
.A1(n_2510),
.A2(n_588),
.B(n_590),
.Y(n_2989)
);

BUFx3_ASAP7_75t_L g2990 ( 
.A(n_2720),
.Y(n_2990)
);

AOI22xp33_ASAP7_75t_L g2991 ( 
.A1(n_2514),
.A2(n_2704),
.B1(n_2730),
.B2(n_2564),
.Y(n_2991)
);

CKINVDCx20_ASAP7_75t_R g2992 ( 
.A(n_2551),
.Y(n_2992)
);

HB1xp67_ASAP7_75t_L g2993 ( 
.A(n_2475),
.Y(n_2993)
);

BUFx2_ASAP7_75t_SL g2994 ( 
.A(n_2518),
.Y(n_2994)
);

CKINVDCx11_ASAP7_75t_R g2995 ( 
.A(n_2551),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2755),
.Y(n_2996)
);

OAI22xp5_ASAP7_75t_SL g2997 ( 
.A1(n_2773),
.A2(n_591),
.B1(n_592),
.B2(n_593),
.Y(n_2997)
);

OAI22xp33_ASAP7_75t_L g2998 ( 
.A1(n_2514),
.A2(n_591),
.B1(n_592),
.B2(n_595),
.Y(n_2998)
);

OAI22xp33_ASAP7_75t_L g2999 ( 
.A1(n_2629),
.A2(n_595),
.B1(n_596),
.B2(n_597),
.Y(n_2999)
);

BUFx2_ASAP7_75t_L g3000 ( 
.A(n_2735),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2755),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2746),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2746),
.Y(n_3003)
);

INVx1_ASAP7_75t_SL g3004 ( 
.A(n_2730),
.Y(n_3004)
);

AND2x2_ASAP7_75t_L g3005 ( 
.A(n_2626),
.B(n_596),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2677),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2677),
.Y(n_3007)
);

INVx3_ASAP7_75t_L g3008 ( 
.A(n_2499),
.Y(n_3008)
);

OAI22xp5_ASAP7_75t_L g3009 ( 
.A1(n_2535),
.A2(n_597),
.B1(n_598),
.B2(n_599),
.Y(n_3009)
);

AOI21x1_ASAP7_75t_L g3010 ( 
.A1(n_2448),
.A2(n_598),
.B(n_599),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2678),
.Y(n_3011)
);

INVx2_ASAP7_75t_SL g3012 ( 
.A(n_2450),
.Y(n_3012)
);

NAND2x1_ASAP7_75t_L g3013 ( 
.A(n_2535),
.B(n_601),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2678),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2762),
.Y(n_3015)
);

AOI22xp33_ASAP7_75t_SL g3016 ( 
.A1(n_2704),
.A2(n_601),
.B1(n_602),
.B2(n_603),
.Y(n_3016)
);

INVx3_ASAP7_75t_L g3017 ( 
.A(n_2555),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2705),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2751),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2705),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2472),
.Y(n_3021)
);

AOI22xp33_ASAP7_75t_L g3022 ( 
.A1(n_2704),
.A2(n_2730),
.B1(n_2564),
.B2(n_2817),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2751),
.Y(n_3023)
);

OAI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_2586),
.A2(n_602),
.B1(n_603),
.B2(n_605),
.Y(n_3024)
);

AOI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_2704),
.A2(n_605),
.B1(n_606),
.B2(n_607),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2472),
.Y(n_3026)
);

INVx3_ASAP7_75t_L g3027 ( 
.A(n_2555),
.Y(n_3027)
);

AOI22xp33_ASAP7_75t_SL g3028 ( 
.A1(n_2704),
.A2(n_606),
.B1(n_607),
.B2(n_608),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_2632),
.B(n_609),
.Y(n_3029)
);

AOI22xp33_ASAP7_75t_L g3030 ( 
.A1(n_2817),
.A2(n_610),
.B1(n_611),
.B2(n_612),
.Y(n_3030)
);

CKINVDCx20_ASAP7_75t_R g3031 ( 
.A(n_2452),
.Y(n_3031)
);

BUFx2_ASAP7_75t_R g3032 ( 
.A(n_2619),
.Y(n_3032)
);

BUFx3_ASAP7_75t_L g3033 ( 
.A(n_2660),
.Y(n_3033)
);

OA21x2_ASAP7_75t_L g3034 ( 
.A1(n_2795),
.A2(n_611),
.B(n_612),
.Y(n_3034)
);

BUFx3_ASAP7_75t_L g3035 ( 
.A(n_2660),
.Y(n_3035)
);

AND2x2_ASAP7_75t_L g3036 ( 
.A(n_2659),
.B(n_613),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2734),
.B(n_614),
.Y(n_3037)
);

INVxp67_ASAP7_75t_SL g3038 ( 
.A(n_2611),
.Y(n_3038)
);

INVx4_ASAP7_75t_L g3039 ( 
.A(n_2683),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2757),
.Y(n_3040)
);

AOI22xp33_ASAP7_75t_L g3041 ( 
.A1(n_2822),
.A2(n_614),
.B1(n_615),
.B2(n_616),
.Y(n_3041)
);

AOI22xp5_ASAP7_75t_L g3042 ( 
.A1(n_2697),
.A2(n_615),
.B1(n_616),
.B2(n_617),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2517),
.Y(n_3043)
);

BUFx2_ASAP7_75t_R g3044 ( 
.A(n_2701),
.Y(n_3044)
);

OAI22xp5_ASAP7_75t_L g3045 ( 
.A1(n_2628),
.A2(n_617),
.B1(n_620),
.B2(n_621),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2679),
.B(n_620),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2749),
.B(n_621),
.Y(n_3047)
);

BUFx3_ASAP7_75t_L g3048 ( 
.A(n_2606),
.Y(n_3048)
);

CKINVDCx20_ASAP7_75t_R g3049 ( 
.A(n_2643),
.Y(n_3049)
);

AOI22xp33_ASAP7_75t_L g3050 ( 
.A1(n_2822),
.A2(n_623),
.B1(n_624),
.B2(n_625),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2517),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2694),
.B(n_623),
.Y(n_3052)
);

AND2x4_ASAP7_75t_L g3053 ( 
.A(n_2556),
.B(n_624),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2546),
.Y(n_3054)
);

AOI22xp33_ASAP7_75t_L g3055 ( 
.A1(n_2830),
.A2(n_625),
.B1(n_626),
.B2(n_627),
.Y(n_3055)
);

HB1xp67_ASAP7_75t_L g3056 ( 
.A(n_2512),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2757),
.Y(n_3057)
);

INVx4_ASAP7_75t_SL g3058 ( 
.A(n_2735),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_2470),
.B(n_2565),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2546),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2687),
.Y(n_3061)
);

OAI21x1_ASAP7_75t_SL g3062 ( 
.A1(n_2682),
.A2(n_627),
.B(n_628),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2687),
.Y(n_3063)
);

INVx3_ASAP7_75t_L g3064 ( 
.A(n_2683),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2740),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2793),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2750),
.B(n_628),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2793),
.Y(n_3068)
);

OAI22xp5_ASAP7_75t_L g3069 ( 
.A1(n_2653),
.A2(n_629),
.B1(n_630),
.B2(n_631),
.Y(n_3069)
);

OAI21xp5_ASAP7_75t_L g3070 ( 
.A1(n_2490),
.A2(n_629),
.B(n_630),
.Y(n_3070)
);

INVx1_ASAP7_75t_SL g3071 ( 
.A(n_2563),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2757),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2752),
.Y(n_3073)
);

AOI22xp5_ASAP7_75t_L g3074 ( 
.A1(n_2697),
.A2(n_632),
.B1(n_634),
.B2(n_635),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2752),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2728),
.Y(n_3076)
);

AOI22xp33_ASAP7_75t_SL g3077 ( 
.A1(n_2653),
.A2(n_634),
.B1(n_635),
.B2(n_636),
.Y(n_3077)
);

OAI22xp33_ASAP7_75t_L g3078 ( 
.A1(n_2812),
.A2(n_637),
.B1(n_638),
.B2(n_639),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2728),
.Y(n_3079)
);

BUFx2_ASAP7_75t_L g3080 ( 
.A(n_2643),
.Y(n_3080)
);

CKINVDCx20_ASAP7_75t_R g3081 ( 
.A(n_2451),
.Y(n_3081)
);

OAI22xp5_ASAP7_75t_L g3082 ( 
.A1(n_2674),
.A2(n_638),
.B1(n_640),
.B2(n_641),
.Y(n_3082)
);

OA21x2_ASAP7_75t_L g3083 ( 
.A1(n_2819),
.A2(n_642),
.B(n_643),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2789),
.Y(n_3084)
);

BUFx2_ASAP7_75t_R g3085 ( 
.A(n_2721),
.Y(n_3085)
);

OAI22xp5_ASAP7_75t_L g3086 ( 
.A1(n_2674),
.A2(n_644),
.B1(n_646),
.B2(n_647),
.Y(n_3086)
);

BUFx8_ASAP7_75t_L g3087 ( 
.A(n_2492),
.Y(n_3087)
);

AOI21x1_ASAP7_75t_L g3088 ( 
.A1(n_2448),
.A2(n_644),
.B(n_646),
.Y(n_3088)
);

OAI21x1_ASAP7_75t_L g3089 ( 
.A1(n_2604),
.A2(n_648),
.B(n_649),
.Y(n_3089)
);

BUFx12f_ASAP7_75t_L g3090 ( 
.A(n_2495),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2789),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2688),
.Y(n_3092)
);

AO21x2_ASAP7_75t_L g3093 ( 
.A1(n_2479),
.A2(n_743),
.B(n_650),
.Y(n_3093)
);

AOI22xp33_ASAP7_75t_L g3094 ( 
.A1(n_2830),
.A2(n_649),
.B1(n_651),
.B2(n_653),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2688),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2786),
.Y(n_3096)
);

AND2x4_ASAP7_75t_L g3097 ( 
.A(n_2556),
.B(n_653),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2786),
.Y(n_3098)
);

BUFx3_ASAP7_75t_L g3099 ( 
.A(n_2544),
.Y(n_3099)
);

AOI22xp33_ASAP7_75t_L g3100 ( 
.A1(n_2681),
.A2(n_2797),
.B1(n_2769),
.B2(n_2451),
.Y(n_3100)
);

INVx1_ASAP7_75t_SL g3101 ( 
.A(n_2563),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_2519),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2521),
.Y(n_3103)
);

OAI22xp5_ASAP7_75t_L g3104 ( 
.A1(n_2681),
.A2(n_654),
.B1(n_655),
.B2(n_656),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2703),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2714),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2712),
.Y(n_3107)
);

OR2x2_ASAP7_75t_L g3108 ( 
.A(n_2706),
.B(n_655),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2712),
.Y(n_3109)
);

INVx1_ASAP7_75t_SL g3110 ( 
.A(n_2563),
.Y(n_3110)
);

CKINVDCx20_ASAP7_75t_R g3111 ( 
.A(n_2451),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2724),
.Y(n_3112)
);

BUFx2_ASAP7_75t_L g3113 ( 
.A(n_2455),
.Y(n_3113)
);

NAND2x1p5_ASAP7_75t_L g3114 ( 
.A(n_2691),
.B(n_656),
.Y(n_3114)
);

OAI21xp5_ASAP7_75t_SL g3115 ( 
.A1(n_2747),
.A2(n_657),
.B(n_658),
.Y(n_3115)
);

CKINVDCx20_ASAP7_75t_R g3116 ( 
.A(n_2738),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2778),
.Y(n_3117)
);

HB1xp67_ASAP7_75t_L g3118 ( 
.A(n_2549),
.Y(n_3118)
);

CKINVDCx11_ASAP7_75t_R g3119 ( 
.A(n_2695),
.Y(n_3119)
);

OA21x2_ASAP7_75t_L g3120 ( 
.A1(n_2613),
.A2(n_657),
.B(n_659),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2807),
.Y(n_3121)
);

BUFx2_ASAP7_75t_L g3122 ( 
.A(n_2455),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2565),
.Y(n_3123)
);

AND2x2_ASAP7_75t_L g3124 ( 
.A(n_2621),
.B(n_659),
.Y(n_3124)
);

INVx3_ASAP7_75t_L g3125 ( 
.A(n_2683),
.Y(n_3125)
);

AOI21x1_ASAP7_75t_L g3126 ( 
.A1(n_2448),
.A2(n_660),
.B(n_661),
.Y(n_3126)
);

AND2x2_ASAP7_75t_L g3127 ( 
.A(n_2621),
.B(n_661),
.Y(n_3127)
);

INVx3_ASAP7_75t_L g3128 ( 
.A(n_2600),
.Y(n_3128)
);

BUFx2_ASAP7_75t_L g3129 ( 
.A(n_2468),
.Y(n_3129)
);

BUFx2_ASAP7_75t_L g3130 ( 
.A(n_2468),
.Y(n_3130)
);

INVx3_ASAP7_75t_L g3131 ( 
.A(n_2600),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2542),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2790),
.B(n_662),
.Y(n_3133)
);

AOI22xp33_ASAP7_75t_SL g3134 ( 
.A1(n_2814),
.A2(n_662),
.B1(n_663),
.B2(n_664),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2543),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_L g3136 ( 
.A1(n_2797),
.A2(n_663),
.B1(n_665),
.B2(n_666),
.Y(n_3136)
);

AOI22xp33_ASAP7_75t_L g3137 ( 
.A1(n_2769),
.A2(n_665),
.B1(n_668),
.B2(n_669),
.Y(n_3137)
);

INVx3_ASAP7_75t_L g3138 ( 
.A(n_2608),
.Y(n_3138)
);

OAI22xp33_ASAP7_75t_L g3139 ( 
.A1(n_2810),
.A2(n_670),
.B1(n_671),
.B2(n_672),
.Y(n_3139)
);

INVx6_ASAP7_75t_L g3140 ( 
.A(n_2648),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2781),
.B(n_670),
.Y(n_3141)
);

AOI21x1_ASAP7_75t_L g3142 ( 
.A1(n_2531),
.A2(n_671),
.B(n_672),
.Y(n_3142)
);

AOI22xp33_ASAP7_75t_SL g3143 ( 
.A1(n_2814),
.A2(n_673),
.B1(n_675),
.B2(n_676),
.Y(n_3143)
);

AOI21x1_ASAP7_75t_L g3144 ( 
.A1(n_2531),
.A2(n_676),
.B(n_677),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2767),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_2500),
.B(n_678),
.Y(n_3146)
);

INVx2_ASAP7_75t_SL g3147 ( 
.A(n_2450),
.Y(n_3147)
);

BUFx3_ASAP7_75t_L g3148 ( 
.A(n_2530),
.Y(n_3148)
);

NAND2x1p5_ASAP7_75t_L g3149 ( 
.A(n_2691),
.B(n_678),
.Y(n_3149)
);

AOI22xp33_ASAP7_75t_SL g3150 ( 
.A1(n_2810),
.A2(n_679),
.B1(n_680),
.B2(n_681),
.Y(n_3150)
);

BUFx2_ASAP7_75t_L g3151 ( 
.A(n_2480),
.Y(n_3151)
);

INVxp67_ASAP7_75t_L g3152 ( 
.A(n_2662),
.Y(n_3152)
);

AOI21x1_ASAP7_75t_L g3153 ( 
.A1(n_2531),
.A2(n_679),
.B(n_681),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2511),
.Y(n_3154)
);

INVx2_ASAP7_75t_SL g3155 ( 
.A(n_2462),
.Y(n_3155)
);

AOI22xp5_ASAP7_75t_L g3156 ( 
.A1(n_2738),
.A2(n_682),
.B1(n_683),
.B2(n_684),
.Y(n_3156)
);

CKINVDCx20_ASAP7_75t_R g3157 ( 
.A(n_2695),
.Y(n_3157)
);

AOI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_2533),
.A2(n_682),
.B(n_685),
.Y(n_3158)
);

BUFx2_ASAP7_75t_R g3159 ( 
.A(n_2549),
.Y(n_3159)
);

AO21x2_ASAP7_75t_L g3160 ( 
.A1(n_2487),
.A2(n_742),
.B(n_686),
.Y(n_3160)
);

BUFx2_ASAP7_75t_L g3161 ( 
.A(n_2480),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2500),
.Y(n_3162)
);

OAI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2490),
.A2(n_685),
.B(n_686),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2796),
.Y(n_3164)
);

OAI22xp33_ASAP7_75t_L g3165 ( 
.A1(n_2668),
.A2(n_687),
.B1(n_688),
.B2(n_689),
.Y(n_3165)
);

AOI21x1_ASAP7_75t_L g3166 ( 
.A1(n_2791),
.A2(n_687),
.B(n_688),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2796),
.Y(n_3167)
);

AND2x2_ASAP7_75t_L g3168 ( 
.A(n_2650),
.B(n_690),
.Y(n_3168)
);

AND2x2_ASAP7_75t_L g3169 ( 
.A(n_2780),
.B(n_2828),
.Y(n_3169)
);

AND2x4_ASAP7_75t_L g3170 ( 
.A(n_2691),
.B(n_690),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2798),
.Y(n_3171)
);

BUFx2_ASAP7_75t_L g3172 ( 
.A(n_2744),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2798),
.Y(n_3173)
);

CKINVDCx11_ASAP7_75t_R g3174 ( 
.A(n_2745),
.Y(n_3174)
);

NOR2xp67_ASAP7_75t_R g3175 ( 
.A(n_2691),
.B(n_691),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2739),
.Y(n_3176)
);

BUFx4f_ASAP7_75t_SL g3177 ( 
.A(n_2763),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_2875),
.B(n_2610),
.Y(n_3178)
);

OAI22xp5_ASAP7_75t_L g3179 ( 
.A1(n_2859),
.A2(n_2672),
.B1(n_2668),
.B2(n_2574),
.Y(n_3179)
);

OAI22xp5_ASAP7_75t_L g3180 ( 
.A1(n_3025),
.A2(n_2672),
.B1(n_2574),
.B2(n_2501),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2834),
.Y(n_3181)
);

HB1xp67_ASAP7_75t_L g3182 ( 
.A(n_2954),
.Y(n_3182)
);

CKINVDCx5p33_ASAP7_75t_R g3183 ( 
.A(n_2866),
.Y(n_3183)
);

AOI22xp33_ASAP7_75t_L g3184 ( 
.A1(n_2927),
.A2(n_2799),
.B1(n_2736),
.B2(n_2775),
.Y(n_3184)
);

AND2x4_ASAP7_75t_L g3185 ( 
.A(n_3039),
.B(n_2612),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_3005),
.B(n_3029),
.Y(n_3186)
);

BUFx3_ASAP7_75t_L g3187 ( 
.A(n_2862),
.Y(n_3187)
);

AND2x2_ASAP7_75t_L g3188 ( 
.A(n_3036),
.B(n_2610),
.Y(n_3188)
);

AND2x2_ASAP7_75t_L g3189 ( 
.A(n_3046),
.B(n_2616),
.Y(n_3189)
);

OAI22xp5_ASAP7_75t_L g3190 ( 
.A1(n_3025),
.A2(n_2485),
.B1(n_2488),
.B2(n_2580),
.Y(n_3190)
);

OR2x2_ASAP7_75t_L g3191 ( 
.A(n_2863),
.B(n_2467),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2833),
.Y(n_3192)
);

NOR2x1_ASAP7_75t_SL g3193 ( 
.A(n_2901),
.B(n_2994),
.Y(n_3193)
);

AOI22xp33_ASAP7_75t_L g3194 ( 
.A1(n_2927),
.A2(n_2829),
.B1(n_2715),
.B2(n_2463),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3117),
.B(n_2813),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2836),
.Y(n_3196)
);

BUFx3_ASAP7_75t_L g3197 ( 
.A(n_2862),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2858),
.B(n_2813),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_3059),
.B(n_2783),
.Y(n_3199)
);

NOR2xp33_ASAP7_75t_R g3200 ( 
.A(n_2932),
.B(n_2558),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_2837),
.Y(n_3201)
);

NOR3xp33_ASAP7_75t_SL g3202 ( 
.A(n_2919),
.B(n_2733),
.C(n_2662),
.Y(n_3202)
);

OR2x6_ASAP7_75t_L g3203 ( 
.A(n_3000),
.B(n_2707),
.Y(n_3203)
);

NOR3xp33_ASAP7_75t_SL g3204 ( 
.A(n_2997),
.B(n_2733),
.C(n_2558),
.Y(n_3204)
);

NOR2xp33_ASAP7_75t_R g3205 ( 
.A(n_2854),
.B(n_2596),
.Y(n_3205)
);

NOR3xp33_ASAP7_75t_SL g3206 ( 
.A(n_2997),
.B(n_2596),
.C(n_2792),
.Y(n_3206)
);

INVx2_ASAP7_75t_L g3207 ( 
.A(n_2840),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_3123),
.B(n_2809),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2839),
.Y(n_3209)
);

NOR2x1p5_ASAP7_75t_L g3210 ( 
.A(n_2877),
.B(n_2933),
.Y(n_3210)
);

OR2x2_ASAP7_75t_L g3211 ( 
.A(n_2863),
.B(n_2663),
.Y(n_3211)
);

NOR3xp33_ASAP7_75t_SL g3212 ( 
.A(n_3115),
.B(n_2792),
.C(n_2759),
.Y(n_3212)
);

CKINVDCx20_ASAP7_75t_R g3213 ( 
.A(n_2856),
.Y(n_3213)
);

CKINVDCx16_ASAP7_75t_R g3214 ( 
.A(n_2861),
.Y(n_3214)
);

NOR2xp33_ASAP7_75t_R g3215 ( 
.A(n_2862),
.B(n_3049),
.Y(n_3215)
);

AND2x2_ASAP7_75t_L g3216 ( 
.A(n_3052),
.B(n_2616),
.Y(n_3216)
);

CKINVDCx5p33_ASAP7_75t_R g3217 ( 
.A(n_2912),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2841),
.B(n_2615),
.Y(n_3218)
);

INVx3_ASAP7_75t_L g3219 ( 
.A(n_2908),
.Y(n_3219)
);

NAND3xp33_ASAP7_75t_SL g3220 ( 
.A(n_3150),
.B(n_2802),
.C(n_2488),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2847),
.Y(n_3221)
);

AND2x4_ASAP7_75t_L g3222 ( 
.A(n_3039),
.B(n_2954),
.Y(n_3222)
);

CKINVDCx5p33_ASAP7_75t_R g3223 ( 
.A(n_3087),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2851),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_2850),
.Y(n_3225)
);

CKINVDCx5p33_ASAP7_75t_R g3226 ( 
.A(n_3087),
.Y(n_3226)
);

OAI22xp33_ASAP7_75t_L g3227 ( 
.A1(n_3042),
.A2(n_2725),
.B1(n_2485),
.B2(n_2739),
.Y(n_3227)
);

NOR2xp33_ASAP7_75t_R g3228 ( 
.A(n_2855),
.B(n_2462),
.Y(n_3228)
);

AOI22xp33_ASAP7_75t_L g3229 ( 
.A1(n_2921),
.A2(n_2831),
.B1(n_2756),
.B2(n_2811),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2873),
.B(n_2639),
.Y(n_3230)
);

AOI22xp33_ASAP7_75t_L g3231 ( 
.A1(n_2849),
.A2(n_2831),
.B1(n_2756),
.B2(n_2784),
.Y(n_3231)
);

CKINVDCx16_ASAP7_75t_R g3232 ( 
.A(n_2894),
.Y(n_3232)
);

CKINVDCx5p33_ASAP7_75t_R g3233 ( 
.A(n_2936),
.Y(n_3233)
);

OAI22xp5_ASAP7_75t_L g3234 ( 
.A1(n_2991),
.A2(n_2627),
.B1(n_2502),
.B2(n_2520),
.Y(n_3234)
);

NAND2xp33_ASAP7_75t_SL g3235 ( 
.A(n_2885),
.B(n_2725),
.Y(n_3235)
);

BUFx2_ASAP7_75t_SL g3236 ( 
.A(n_3033),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2878),
.B(n_2784),
.Y(n_3237)
);

AOI22xp33_ASAP7_75t_SL g3238 ( 
.A1(n_2885),
.A2(n_2638),
.B1(n_2640),
.B2(n_2612),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2853),
.Y(n_3239)
);

CKINVDCx5p33_ASAP7_75t_R g3240 ( 
.A(n_2995),
.Y(n_3240)
);

AOI22xp5_ASAP7_75t_L g3241 ( 
.A1(n_2876),
.A2(n_2763),
.B1(n_2759),
.B2(n_2824),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_2857),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_2973),
.B(n_2530),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_3133),
.B(n_2741),
.Y(n_3244)
);

AND2x4_ASAP7_75t_L g3245 ( 
.A(n_2981),
.B(n_2638),
.Y(n_3245)
);

AO31x2_ASAP7_75t_L g3246 ( 
.A1(n_3102),
.A2(n_2684),
.A3(n_2545),
.B(n_2550),
.Y(n_3246)
);

AND2x2_ASAP7_75t_L g3247 ( 
.A(n_2864),
.B(n_2780),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2880),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_2884),
.B(n_2787),
.Y(n_3249)
);

NAND2xp33_ASAP7_75t_R g3250 ( 
.A(n_2890),
.B(n_2640),
.Y(n_3250)
);

AND2x2_ASAP7_75t_L g3251 ( 
.A(n_2981),
.B(n_2635),
.Y(n_3251)
);

INVxp67_ASAP7_75t_L g3252 ( 
.A(n_2928),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_2869),
.Y(n_3253)
);

AND2x2_ASAP7_75t_L g3254 ( 
.A(n_3169),
.B(n_2635),
.Y(n_3254)
);

OR2x6_ASAP7_75t_L g3255 ( 
.A(n_3012),
.B(n_2562),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_2870),
.B(n_2644),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2892),
.Y(n_3257)
);

CKINVDCx5p33_ASAP7_75t_R g3258 ( 
.A(n_2893),
.Y(n_3258)
);

INVx6_ASAP7_75t_L g3259 ( 
.A(n_3058),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_2896),
.Y(n_3260)
);

INVx2_ASAP7_75t_SL g3261 ( 
.A(n_3058),
.Y(n_3261)
);

AND2x4_ASAP7_75t_L g3262 ( 
.A(n_2881),
.B(n_2905),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_2870),
.B(n_2644),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_2897),
.B(n_2787),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_2955),
.B(n_2711),
.Y(n_3265)
);

NOR3xp33_ASAP7_75t_SL g3266 ( 
.A(n_3115),
.B(n_2967),
.C(n_2999),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2902),
.Y(n_3267)
);

HB1xp67_ASAP7_75t_L g3268 ( 
.A(n_2972),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_2872),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_2996),
.B(n_3001),
.Y(n_3270)
);

CKINVDCx5p33_ASAP7_75t_R g3271 ( 
.A(n_2917),
.Y(n_3271)
);

INVx2_ASAP7_75t_SL g3272 ( 
.A(n_3058),
.Y(n_3272)
);

OAI22xp33_ASAP7_75t_SL g3273 ( 
.A1(n_3013),
.A2(n_2627),
.B1(n_2502),
.B2(n_2520),
.Y(n_3273)
);

NAND2xp33_ASAP7_75t_R g3274 ( 
.A(n_2907),
.B(n_3080),
.Y(n_3274)
);

NAND2xp33_ASAP7_75t_R g3275 ( 
.A(n_3159),
.B(n_2914),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_3148),
.B(n_2676),
.Y(n_3276)
);

HB1xp67_ASAP7_75t_L g3277 ( 
.A(n_2915),
.Y(n_3277)
);

BUFx2_ASAP7_75t_L g3278 ( 
.A(n_2883),
.Y(n_3278)
);

OR2x2_ASAP7_75t_L g3279 ( 
.A(n_2882),
.B(n_2537),
.Y(n_3279)
);

BUFx8_ASAP7_75t_L g3280 ( 
.A(n_3147),
.Y(n_3280)
);

AND2x4_ASAP7_75t_L g3281 ( 
.A(n_2881),
.B(n_2647),
.Y(n_3281)
);

NAND4xp25_ASAP7_75t_L g3282 ( 
.A(n_3042),
.B(n_2764),
.C(n_2808),
.D(n_2804),
.Y(n_3282)
);

OAI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_2989),
.A2(n_2748),
.B(n_2808),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_2918),
.B(n_2800),
.Y(n_3284)
);

NAND2xp33_ASAP7_75t_R g3285 ( 
.A(n_3159),
.B(n_2647),
.Y(n_3285)
);

INVx3_ASAP7_75t_L g3286 ( 
.A(n_3035),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2920),
.Y(n_3287)
);

NAND3xp33_ASAP7_75t_L g3288 ( 
.A(n_2947),
.B(n_2573),
.C(n_2553),
.Y(n_3288)
);

OR2x6_ASAP7_75t_L g3289 ( 
.A(n_3155),
.B(n_2581),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2931),
.B(n_2816),
.Y(n_3290)
);

AND2x2_ASAP7_75t_L g3291 ( 
.A(n_2843),
.B(n_2537),
.Y(n_3291)
);

HB1xp67_ASAP7_75t_L g3292 ( 
.A(n_2916),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_2934),
.Y(n_3293)
);

AO31x2_ASAP7_75t_L g3294 ( 
.A1(n_3103),
.A2(n_2545),
.A3(n_2550),
.B(n_2527),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_3146),
.B(n_2449),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2937),
.B(n_2823),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2938),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2939),
.Y(n_3298)
);

NAND2xp33_ASAP7_75t_R g3299 ( 
.A(n_2957),
.B(n_2449),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_2940),
.Y(n_3300)
);

AOI22xp33_ASAP7_75t_L g3301 ( 
.A1(n_2860),
.A2(n_2651),
.B1(n_2497),
.B2(n_2637),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_2951),
.B(n_2803),
.Y(n_3302)
);

NAND2xp33_ASAP7_75t_R g3303 ( 
.A(n_2905),
.B(n_2453),
.Y(n_3303)
);

NOR2xp33_ASAP7_75t_R g3304 ( 
.A(n_2965),
.B(n_2648),
.Y(n_3304)
);

AND2x4_ASAP7_75t_L g3305 ( 
.A(n_2922),
.B(n_2453),
.Y(n_3305)
);

AOI22xp33_ASAP7_75t_L g3306 ( 
.A1(n_2923),
.A2(n_2636),
.B1(n_2666),
.B2(n_2607),
.Y(n_3306)
);

NOR2xp33_ASAP7_75t_R g3307 ( 
.A(n_3031),
.B(n_2648),
.Y(n_3307)
);

HB1xp67_ASAP7_75t_L g3308 ( 
.A(n_2982),
.Y(n_3308)
);

AOI22xp33_ASAP7_75t_L g3309 ( 
.A1(n_2923),
.A2(n_2602),
.B1(n_2673),
.B2(n_2758),
.Y(n_3309)
);

NAND2xp33_ASAP7_75t_R g3310 ( 
.A(n_2922),
.B(n_2469),
.Y(n_3310)
);

AOI22xp33_ASAP7_75t_L g3311 ( 
.A1(n_2945),
.A2(n_2698),
.B1(n_2709),
.B2(n_2680),
.Y(n_3311)
);

CKINVDCx5p33_ASAP7_75t_R g3312 ( 
.A(n_2865),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2953),
.Y(n_3313)
);

CKINVDCx16_ASAP7_75t_R g3314 ( 
.A(n_2992),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2956),
.Y(n_3315)
);

NOR2xp33_ASAP7_75t_R g3316 ( 
.A(n_2944),
.B(n_2745),
.Y(n_3316)
);

NAND3xp33_ASAP7_75t_L g3317 ( 
.A(n_2844),
.B(n_2719),
.C(n_2713),
.Y(n_3317)
);

BUFx12f_ASAP7_75t_L g3318 ( 
.A(n_3174),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_2960),
.Y(n_3319)
);

OR2x6_ASAP7_75t_L g3320 ( 
.A(n_3118),
.B(n_2774),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3162),
.B(n_2805),
.Y(n_3321)
);

CKINVDCx16_ASAP7_75t_R g3322 ( 
.A(n_3157),
.Y(n_3322)
);

AOI22xp33_ASAP7_75t_L g3323 ( 
.A1(n_2891),
.A2(n_2876),
.B1(n_2848),
.B2(n_2984),
.Y(n_3323)
);

NAND3xp33_ASAP7_75t_SL g3324 ( 
.A(n_3150),
.B(n_2584),
.C(n_2515),
.Y(n_3324)
);

NOR2xp33_ASAP7_75t_L g3325 ( 
.A(n_2888),
.B(n_2459),
.Y(n_3325)
);

CKINVDCx5p33_ASAP7_75t_R g3326 ( 
.A(n_2911),
.Y(n_3326)
);

CKINVDCx5p33_ASAP7_75t_R g3327 ( 
.A(n_3119),
.Y(n_3327)
);

BUFx3_ASAP7_75t_L g3328 ( 
.A(n_2935),
.Y(n_3328)
);

NAND2xp33_ASAP7_75t_R g3329 ( 
.A(n_3008),
.B(n_2469),
.Y(n_3329)
);

NOR2xp33_ASAP7_75t_R g3330 ( 
.A(n_2944),
.B(n_3081),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_2963),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_R g3332 ( 
.A(n_3111),
.B(n_2585),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2968),
.B(n_2805),
.Y(n_3333)
);

NOR3xp33_ASAP7_75t_SL g3334 ( 
.A(n_2967),
.B(n_2815),
.C(n_2459),
.Y(n_3334)
);

OR2x6_ASAP7_75t_L g3335 ( 
.A(n_2887),
.B(n_2515),
.Y(n_3335)
);

O2A1O1Ixp33_ASAP7_75t_SL g3336 ( 
.A1(n_2984),
.A2(n_2579),
.B(n_2815),
.C(n_2699),
.Y(n_3336)
);

NOR3xp33_ASAP7_75t_SL g3337 ( 
.A(n_2998),
.B(n_2532),
.C(n_2483),
.Y(n_3337)
);

AND2x2_ASAP7_75t_L g3338 ( 
.A(n_3048),
.B(n_2770),
.Y(n_3338)
);

NAND2xp33_ASAP7_75t_SL g3339 ( 
.A(n_3022),
.B(n_3009),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_R g3340 ( 
.A(n_3116),
.B(n_2585),
.Y(n_3340)
);

AOI22xp33_ASAP7_75t_L g3341 ( 
.A1(n_2891),
.A2(n_2642),
.B1(n_2669),
.B2(n_2505),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_2970),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_2974),
.B(n_3065),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_2975),
.Y(n_3344)
);

NOR2xp33_ASAP7_75t_R g3345 ( 
.A(n_3090),
.B(n_2585),
.Y(n_3345)
);

BUFx3_ASAP7_75t_L g3346 ( 
.A(n_2976),
.Y(n_3346)
);

NOR2x1_ASAP7_75t_L g3347 ( 
.A(n_3009),
.B(n_2693),
.Y(n_3347)
);

CKINVDCx5p33_ASAP7_75t_R g3348 ( 
.A(n_2845),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3092),
.B(n_2670),
.Y(n_3349)
);

NAND2xp33_ASAP7_75t_SL g3350 ( 
.A(n_3053),
.B(n_3097),
.Y(n_3350)
);

AND2x2_ASAP7_75t_L g3351 ( 
.A(n_2883),
.B(n_3176),
.Y(n_3351)
);

AND2x2_ASAP7_75t_L g3352 ( 
.A(n_3124),
.B(n_693),
.Y(n_3352)
);

OR2x2_ASAP7_75t_L g3353 ( 
.A(n_2882),
.B(n_2693),
.Y(n_3353)
);

AND2x2_ASAP7_75t_L g3354 ( 
.A(n_3127),
.B(n_694),
.Y(n_3354)
);

NOR2xp33_ASAP7_75t_R g3355 ( 
.A(n_2966),
.B(n_2641),
.Y(n_3355)
);

NOR2xp33_ASAP7_75t_R g3356 ( 
.A(n_2971),
.B(n_2641),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3076),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3095),
.B(n_2670),
.Y(n_3358)
);

HB1xp67_ASAP7_75t_L g3359 ( 
.A(n_2993),
.Y(n_3359)
);

NOR3xp33_ASAP7_75t_SL g3360 ( 
.A(n_3139),
.B(n_2532),
.C(n_2483),
.Y(n_3360)
);

CKINVDCx5p33_ASAP7_75t_R g3361 ( 
.A(n_2846),
.Y(n_3361)
);

CKINVDCx20_ASAP7_75t_R g3362 ( 
.A(n_3177),
.Y(n_3362)
);

CKINVDCx16_ASAP7_75t_R g3363 ( 
.A(n_2909),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3079),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3084),
.Y(n_3365)
);

NOR2x1_ASAP7_75t_R g3366 ( 
.A(n_2924),
.B(n_2567),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_2930),
.B(n_694),
.Y(n_3367)
);

BUFx6f_ASAP7_75t_L g3368 ( 
.A(n_2887),
.Y(n_3368)
);

INVx3_ASAP7_75t_L g3369 ( 
.A(n_3008),
.Y(n_3369)
);

NAND2xp33_ASAP7_75t_R g3370 ( 
.A(n_3064),
.B(n_2469),
.Y(n_3370)
);

OR2x6_ASAP7_75t_L g3371 ( 
.A(n_3152),
.B(n_2584),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3091),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3037),
.Y(n_3373)
);

AND2x4_ASAP7_75t_L g3374 ( 
.A(n_3064),
.B(n_2559),
.Y(n_3374)
);

NOR2xp33_ASAP7_75t_R g3375 ( 
.A(n_3017),
.B(n_2641),
.Y(n_3375)
);

NOR2xp33_ASAP7_75t_R g3376 ( 
.A(n_3017),
.B(n_2717),
.Y(n_3376)
);

CKINVDCx20_ASAP7_75t_R g3377 ( 
.A(n_3099),
.Y(n_3377)
);

OR2x2_ASAP7_75t_L g3378 ( 
.A(n_2941),
.B(n_2702),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_3047),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_2978),
.B(n_2702),
.Y(n_3380)
);

CKINVDCx5p33_ASAP7_75t_R g3381 ( 
.A(n_3032),
.Y(n_3381)
);

CKINVDCx11_ASAP7_75t_R g3382 ( 
.A(n_2990),
.Y(n_3382)
);

CKINVDCx20_ASAP7_75t_R g3383 ( 
.A(n_3172),
.Y(n_3383)
);

NOR2xp33_ASAP7_75t_R g3384 ( 
.A(n_3027),
.B(n_2717),
.Y(n_3384)
);

CKINVDCx16_ASAP7_75t_R g3385 ( 
.A(n_3074),
.Y(n_3385)
);

AND2x2_ASAP7_75t_L g3386 ( 
.A(n_2942),
.B(n_2946),
.Y(n_3386)
);

AND2x2_ASAP7_75t_L g3387 ( 
.A(n_2941),
.B(n_695),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_2979),
.B(n_2710),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3047),
.Y(n_3389)
);

NAND2xp33_ASAP7_75t_R g3390 ( 
.A(n_3125),
.B(n_2708),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_2985),
.B(n_2710),
.Y(n_3391)
);

NOR3xp33_ASAP7_75t_SL g3392 ( 
.A(n_2987),
.B(n_2567),
.C(n_2614),
.Y(n_3392)
);

NOR2xp33_ASAP7_75t_R g3393 ( 
.A(n_3125),
.B(n_2717),
.Y(n_3393)
);

OR2x2_ASAP7_75t_L g3394 ( 
.A(n_3056),
.B(n_2820),
.Y(n_3394)
);

BUFx3_ASAP7_75t_L g3395 ( 
.A(n_3140),
.Y(n_3395)
);

AOI22xp33_ASAP7_75t_L g3396 ( 
.A1(n_2848),
.A2(n_2686),
.B1(n_2726),
.B2(n_2722),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3067),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3067),
.Y(n_3398)
);

NOR2xp33_ASAP7_75t_R g3399 ( 
.A(n_3128),
.B(n_2559),
.Y(n_3399)
);

NOR3xp33_ASAP7_75t_SL g3400 ( 
.A(n_3078),
.B(n_2614),
.C(n_2686),
.Y(n_3400)
);

OR2x2_ASAP7_75t_L g3401 ( 
.A(n_2926),
.B(n_2820),
.Y(n_3401)
);

AO31x2_ASAP7_75t_L g3402 ( 
.A1(n_3105),
.A2(n_2675),
.A3(n_2590),
.B(n_2569),
.Y(n_3402)
);

AND2x2_ASAP7_75t_L g3403 ( 
.A(n_3168),
.B(n_696),
.Y(n_3403)
);

INVx2_ASAP7_75t_SL g3404 ( 
.A(n_3140),
.Y(n_3404)
);

NOR2xp33_ASAP7_75t_R g3405 ( 
.A(n_3128),
.B(n_2570),
.Y(n_3405)
);

CKINVDCx16_ASAP7_75t_R g3406 ( 
.A(n_3074),
.Y(n_3406)
);

INVx4_ASAP7_75t_L g3407 ( 
.A(n_3131),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_2986),
.B(n_2722),
.Y(n_3408)
);

INVx2_ASAP7_75t_SL g3409 ( 
.A(n_2838),
.Y(n_3409)
);

HB1xp67_ASAP7_75t_L g3410 ( 
.A(n_3113),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_3122),
.B(n_696),
.Y(n_3411)
);

BUFx3_ASAP7_75t_L g3412 ( 
.A(n_3129),
.Y(n_3412)
);

AND2x4_ASAP7_75t_L g3413 ( 
.A(n_3131),
.B(n_2570),
.Y(n_3413)
);

NOR2xp33_ASAP7_75t_L g3414 ( 
.A(n_2895),
.B(n_2727),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_2977),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3006),
.B(n_2726),
.Y(n_3416)
);

AND2x2_ASAP7_75t_L g3417 ( 
.A(n_3130),
.B(n_698),
.Y(n_3417)
);

AND2x2_ASAP7_75t_L g3418 ( 
.A(n_3151),
.B(n_698),
.Y(n_3418)
);

AOI22xp33_ASAP7_75t_L g3419 ( 
.A1(n_2948),
.A2(n_2625),
.B1(n_2623),
.B2(n_2620),
.Y(n_3419)
);

CKINVDCx5p33_ASAP7_75t_R g3420 ( 
.A(n_3032),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3141),
.Y(n_3421)
);

OR2x2_ASAP7_75t_L g3422 ( 
.A(n_2899),
.B(n_2827),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3096),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_3161),
.B(n_699),
.Y(n_3424)
);

NOR2x1_ASAP7_75t_SL g3425 ( 
.A(n_3107),
.B(n_2631),
.Y(n_3425)
);

AO31x2_ASAP7_75t_L g3426 ( 
.A1(n_3106),
.A2(n_2590),
.A3(n_2593),
.B(n_2599),
.Y(n_3426)
);

OAI22xp5_ASAP7_75t_L g3427 ( 
.A1(n_3016),
.A2(n_2779),
.B1(n_2785),
.B2(n_2685),
.Y(n_3427)
);

CKINVDCx5p33_ASAP7_75t_R g3428 ( 
.A(n_3044),
.Y(n_3428)
);

INVx2_ASAP7_75t_SL g3429 ( 
.A(n_2838),
.Y(n_3429)
);

CKINVDCx5p33_ASAP7_75t_R g3430 ( 
.A(n_3044),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3034),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_2900),
.B(n_700),
.Y(n_3432)
);

NAND2xp33_ASAP7_75t_SL g3433 ( 
.A(n_3053),
.B(n_3097),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3034),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3098),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_3156),
.B(n_700),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_3083),
.Y(n_3437)
);

OR2x6_ASAP7_75t_L g3438 ( 
.A(n_3170),
.B(n_2685),
.Y(n_3438)
);

HB1xp67_ASAP7_75t_L g3439 ( 
.A(n_3002),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_3083),
.Y(n_3440)
);

OR2x6_ASAP7_75t_L g3441 ( 
.A(n_3170),
.B(n_2779),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3156),
.B(n_701),
.Y(n_3442)
);

BUFx2_ASAP7_75t_L g3443 ( 
.A(n_3138),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3066),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3068),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_R g3446 ( 
.A(n_3138),
.B(n_2572),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_3007),
.B(n_2645),
.Y(n_3447)
);

BUFx10_ASAP7_75t_L g3448 ( 
.A(n_3109),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3154),
.Y(n_3449)
);

OR2x6_ASAP7_75t_L g3450 ( 
.A(n_2989),
.B(n_2785),
.Y(n_3450)
);

BUFx4f_ASAP7_75t_SL g3451 ( 
.A(n_2835),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3038),
.Y(n_3452)
);

HB1xp67_ASAP7_75t_L g3453 ( 
.A(n_3003),
.Y(n_3453)
);

NOR2xp33_ASAP7_75t_R g3454 ( 
.A(n_3166),
.B(n_2867),
.Y(n_3454)
);

AND2x4_ASAP7_75t_L g3455 ( 
.A(n_3112),
.B(n_2572),
.Y(n_3455)
);

OR2x6_ASAP7_75t_L g3456 ( 
.A(n_3114),
.B(n_2827),
.Y(n_3456)
);

AND2x2_ASAP7_75t_L g3457 ( 
.A(n_3108),
.B(n_701),
.Y(n_3457)
);

AND2x2_ASAP7_75t_SL g3458 ( 
.A(n_2929),
.B(n_2708),
.Y(n_3458)
);

AOI22xp33_ASAP7_75t_L g3459 ( 
.A1(n_2948),
.A2(n_2592),
.B1(n_2625),
.B2(n_2623),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3073),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_SL g3461 ( 
.A(n_3134),
.B(n_2788),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3075),
.Y(n_3462)
);

AND2x4_ASAP7_75t_L g3463 ( 
.A(n_2929),
.B(n_2577),
.Y(n_3463)
);

AOI22xp33_ASAP7_75t_L g3464 ( 
.A1(n_2949),
.A2(n_2588),
.B1(n_2592),
.B2(n_2620),
.Y(n_3464)
);

AND2x2_ASAP7_75t_L g3465 ( 
.A(n_2969),
.B(n_702),
.Y(n_3465)
);

CKINVDCx20_ASAP7_75t_R g3466 ( 
.A(n_2906),
.Y(n_3466)
);

OAI22xp5_ASAP7_75t_L g3467 ( 
.A1(n_3016),
.A2(n_2821),
.B1(n_2708),
.B2(n_2509),
.Y(n_3467)
);

OAI222xp33_ASAP7_75t_L g3468 ( 
.A1(n_3134),
.A2(n_2454),
.B1(n_2821),
.B2(n_2727),
.C1(n_2731),
.C2(n_2718),
.Y(n_3468)
);

NAND2xp33_ASAP7_75t_R g3469 ( 
.A(n_3120),
.B(n_702),
.Y(n_3469)
);

INVxp67_ASAP7_75t_L g3470 ( 
.A(n_3015),
.Y(n_3470)
);

AND2x4_ASAP7_75t_L g3471 ( 
.A(n_3071),
.B(n_2577),
.Y(n_3471)
);

AND2x2_ASAP7_75t_L g3472 ( 
.A(n_2969),
.B(n_703),
.Y(n_3472)
);

INVx1_ASAP7_75t_SL g3473 ( 
.A(n_3071),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_3192),
.Y(n_3474)
);

AND2x2_ASAP7_75t_L g3475 ( 
.A(n_3386),
.B(n_3101),
.Y(n_3475)
);

AOI22xp33_ASAP7_75t_L g3476 ( 
.A1(n_3339),
.A2(n_3143),
.B1(n_3028),
.B2(n_2874),
.Y(n_3476)
);

OR2x2_ASAP7_75t_L g3477 ( 
.A(n_3182),
.B(n_3101),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3201),
.Y(n_3478)
);

INVx2_ASAP7_75t_L g3479 ( 
.A(n_3207),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3225),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3239),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3242),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3181),
.Y(n_3483)
);

AND2x2_ASAP7_75t_L g3484 ( 
.A(n_3265),
.B(n_3110),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3196),
.Y(n_3485)
);

AND2x2_ASAP7_75t_L g3486 ( 
.A(n_3186),
.B(n_3110),
.Y(n_3486)
);

AND2x2_ASAP7_75t_L g3487 ( 
.A(n_3178),
.B(n_3019),
.Y(n_3487)
);

HB1xp67_ASAP7_75t_L g3488 ( 
.A(n_3410),
.Y(n_3488)
);

BUFx2_ASAP7_75t_L g3489 ( 
.A(n_3399),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3253),
.Y(n_3490)
);

HB1xp67_ASAP7_75t_L g3491 ( 
.A(n_3277),
.Y(n_3491)
);

AND2x2_ASAP7_75t_L g3492 ( 
.A(n_3270),
.B(n_3351),
.Y(n_3492)
);

INVxp67_ASAP7_75t_SL g3493 ( 
.A(n_3193),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_SL g3494 ( 
.A(n_3385),
.B(n_3143),
.Y(n_3494)
);

BUFx2_ASAP7_75t_L g3495 ( 
.A(n_3405),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3470),
.B(n_3023),
.Y(n_3496)
);

AND2x2_ASAP7_75t_L g3497 ( 
.A(n_3439),
.B(n_3028),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_3269),
.Y(n_3498)
);

OAI321xp33_ASAP7_75t_L g3499 ( 
.A1(n_3323),
.A2(n_3082),
.A3(n_3069),
.B1(n_3086),
.B2(n_3024),
.C(n_3045),
.Y(n_3499)
);

OAI33xp33_ASAP7_75t_L g3500 ( 
.A1(n_3179),
.A2(n_3086),
.A3(n_3104),
.B1(n_3082),
.B2(n_3069),
.B3(n_3045),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3209),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3453),
.B(n_3004),
.Y(n_3502)
);

AOI22xp5_ASAP7_75t_L g3503 ( 
.A1(n_3406),
.A2(n_2898),
.B1(n_3104),
.B2(n_2879),
.Y(n_3503)
);

AND2x2_ASAP7_75t_L g3504 ( 
.A(n_3243),
.B(n_3244),
.Y(n_3504)
);

AND2x2_ASAP7_75t_L g3505 ( 
.A(n_3188),
.B(n_3004),
.Y(n_3505)
);

AND2x4_ASAP7_75t_L g3506 ( 
.A(n_3222),
.B(n_3164),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3221),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3224),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3248),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3257),
.Y(n_3510)
);

AOI221xp5_ASAP7_75t_L g3511 ( 
.A1(n_3227),
.A2(n_2886),
.B1(n_3165),
.B2(n_2903),
.C(n_3014),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3415),
.B(n_3011),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3260),
.Y(n_3513)
);

OR2x2_ASAP7_75t_L g3514 ( 
.A(n_3268),
.B(n_3018),
.Y(n_3514)
);

BUFx2_ASAP7_75t_L g3515 ( 
.A(n_3446),
.Y(n_3515)
);

INVxp67_ASAP7_75t_SL g3516 ( 
.A(n_3292),
.Y(n_3516)
);

AND2x2_ASAP7_75t_L g3517 ( 
.A(n_3189),
.B(n_3216),
.Y(n_3517)
);

CKINVDCx5p33_ASAP7_75t_R g3518 ( 
.A(n_3200),
.Y(n_3518)
);

AOI22xp33_ASAP7_75t_SL g3519 ( 
.A1(n_3458),
.A2(n_3062),
.B1(n_3145),
.B2(n_3070),
.Y(n_3519)
);

OR2x2_ASAP7_75t_L g3520 ( 
.A(n_3211),
.B(n_3452),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3267),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3247),
.B(n_3020),
.Y(n_3522)
);

AND2x4_ASAP7_75t_L g3523 ( 
.A(n_3222),
.B(n_3167),
.Y(n_3523)
);

OR2x6_ASAP7_75t_L g3524 ( 
.A(n_3456),
.B(n_3114),
.Y(n_3524)
);

OR2x2_ASAP7_75t_L g3525 ( 
.A(n_3308),
.B(n_3021),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3287),
.Y(n_3526)
);

INVxp67_ASAP7_75t_L g3527 ( 
.A(n_3443),
.Y(n_3527)
);

AND2x2_ASAP7_75t_L g3528 ( 
.A(n_3256),
.B(n_3026),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3293),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3297),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3298),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3357),
.B(n_3364),
.Y(n_3532)
);

INVx3_ASAP7_75t_L g3533 ( 
.A(n_3407),
.Y(n_3533)
);

INVx3_ASAP7_75t_L g3534 ( 
.A(n_3407),
.Y(n_3534)
);

OR2x2_ASAP7_75t_L g3535 ( 
.A(n_3359),
.B(n_3043),
.Y(n_3535)
);

AND2x2_ASAP7_75t_L g3536 ( 
.A(n_3263),
.B(n_3051),
.Y(n_3536)
);

OR2x2_ASAP7_75t_L g3537 ( 
.A(n_3365),
.B(n_3054),
.Y(n_3537)
);

AND2x4_ASAP7_75t_L g3538 ( 
.A(n_3245),
.B(n_3171),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3372),
.B(n_3060),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3254),
.B(n_3061),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3300),
.Y(n_3541)
);

INVx4_ASAP7_75t_L g3542 ( 
.A(n_3259),
.Y(n_3542)
);

OR2x2_ASAP7_75t_L g3543 ( 
.A(n_3191),
.B(n_3063),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_3251),
.B(n_3173),
.Y(n_3544)
);

OR2x2_ASAP7_75t_L g3545 ( 
.A(n_3252),
.B(n_2949),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3313),
.Y(n_3546)
);

AND2x2_ASAP7_75t_L g3547 ( 
.A(n_3295),
.B(n_3040),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3315),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_3367),
.B(n_3057),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3319),
.Y(n_3550)
);

AND2x2_ASAP7_75t_L g3551 ( 
.A(n_3409),
.B(n_3429),
.Y(n_3551)
);

OAI22xp33_ASAP7_75t_L g3552 ( 
.A1(n_3250),
.A2(n_3149),
.B1(n_2852),
.B2(n_3070),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3331),
.Y(n_3553)
);

AND2x4_ASAP7_75t_L g3554 ( 
.A(n_3245),
.B(n_2943),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3342),
.Y(n_3555)
);

OR2x2_ASAP7_75t_L g3556 ( 
.A(n_3199),
.B(n_2980),
.Y(n_3556)
);

AND2x2_ASAP7_75t_L g3557 ( 
.A(n_3473),
.B(n_3072),
.Y(n_3557)
);

INVx2_ASAP7_75t_SL g3558 ( 
.A(n_3259),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3344),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3343),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3237),
.Y(n_3561)
);

NOR2xp67_ASAP7_75t_L g3562 ( 
.A(n_3324),
.B(n_3158),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3412),
.B(n_3077),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3444),
.Y(n_3564)
);

OR2x6_ASAP7_75t_L g3565 ( 
.A(n_3456),
.B(n_3149),
.Y(n_3565)
);

HB1xp67_ASAP7_75t_L g3566 ( 
.A(n_3279),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3445),
.Y(n_3567)
);

AND2x2_ASAP7_75t_L g3568 ( 
.A(n_3449),
.B(n_3077),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3447),
.B(n_2889),
.Y(n_3569)
);

AND2x4_ASAP7_75t_L g3570 ( 
.A(n_3262),
.B(n_3335),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3373),
.B(n_2889),
.Y(n_3571)
);

AND2x2_ASAP7_75t_L g3572 ( 
.A(n_3432),
.B(n_2566),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3423),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3338),
.B(n_2566),
.Y(n_3574)
);

INVxp67_ASAP7_75t_L g3575 ( 
.A(n_3353),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3435),
.Y(n_3576)
);

OAI211xp5_ASAP7_75t_L g3577 ( 
.A1(n_3204),
.A2(n_3100),
.B(n_2988),
.C(n_2983),
.Y(n_3577)
);

AND2x2_ASAP7_75t_L g3578 ( 
.A(n_3387),
.B(n_2959),
.Y(n_3578)
);

BUFx2_ASAP7_75t_L g3579 ( 
.A(n_3355),
.Y(n_3579)
);

NOR2xp33_ASAP7_75t_L g3580 ( 
.A(n_3232),
.B(n_3085),
.Y(n_3580)
);

INVx3_ASAP7_75t_L g3581 ( 
.A(n_3448),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3218),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3230),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3302),
.Y(n_3584)
);

HB1xp67_ASAP7_75t_L g3585 ( 
.A(n_3303),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3195),
.Y(n_3586)
);

AND2x4_ASAP7_75t_L g3587 ( 
.A(n_3335),
.B(n_3121),
.Y(n_3587)
);

OAI22xp5_ASAP7_75t_L g3588 ( 
.A1(n_3238),
.A2(n_2879),
.B1(n_3163),
.B2(n_2964),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3460),
.Y(n_3589)
);

AOI22xp33_ASAP7_75t_L g3590 ( 
.A1(n_3180),
.A2(n_2874),
.B1(n_2961),
.B2(n_3163),
.Y(n_3590)
);

HB1xp67_ASAP7_75t_L g3591 ( 
.A(n_3394),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3462),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3290),
.Y(n_3593)
);

AND2x4_ASAP7_75t_SL g3594 ( 
.A(n_3203),
.B(n_2731),
.Y(n_3594)
);

AND2x2_ASAP7_75t_L g3595 ( 
.A(n_3198),
.B(n_2959),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_3249),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3296),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3264),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3379),
.B(n_3093),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3284),
.Y(n_3600)
);

OR2x2_ASAP7_75t_L g3601 ( 
.A(n_3208),
.B(n_2645),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3401),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3422),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3448),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3389),
.Y(n_3605)
);

AND2x2_ASAP7_75t_L g3606 ( 
.A(n_3291),
.B(n_2818),
.Y(n_3606)
);

INVxp67_ASAP7_75t_SL g3607 ( 
.A(n_3378),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3397),
.B(n_3093),
.Y(n_3608)
);

OAI22xp5_ASAP7_75t_L g3609 ( 
.A1(n_3212),
.A2(n_2964),
.B1(n_2898),
.B2(n_3137),
.Y(n_3609)
);

NOR2x1_ASAP7_75t_L g3610 ( 
.A(n_3220),
.B(n_3160),
.Y(n_3610)
);

AOI22xp5_ASAP7_75t_L g3611 ( 
.A1(n_3436),
.A2(n_3055),
.B1(n_3094),
.B2(n_2950),
.Y(n_3611)
);

AND2x2_ASAP7_75t_L g3612 ( 
.A(n_3278),
.B(n_3352),
.Y(n_3612)
);

OAI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3317),
.A2(n_3158),
.B(n_2958),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_3431),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3398),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3421),
.Y(n_3616)
);

AND2x2_ASAP7_75t_L g3617 ( 
.A(n_3354),
.B(n_2818),
.Y(n_3617)
);

BUFx2_ASAP7_75t_L g3618 ( 
.A(n_3356),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3363),
.B(n_2771),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_3434),
.Y(n_3620)
);

INVx2_ASAP7_75t_L g3621 ( 
.A(n_3437),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3333),
.Y(n_3622)
);

AOI22xp33_ASAP7_75t_L g3623 ( 
.A1(n_3282),
.A2(n_2910),
.B1(n_2925),
.B2(n_2962),
.Y(n_3623)
);

INVx1_ASAP7_75t_SL g3624 ( 
.A(n_3350),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3380),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3440),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_3294),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3349),
.B(n_3358),
.Y(n_3628)
);

AND2x2_ASAP7_75t_L g3629 ( 
.A(n_3411),
.B(n_2771),
.Y(n_3629)
);

AND2x4_ASAP7_75t_L g3630 ( 
.A(n_3371),
.B(n_3132),
.Y(n_3630)
);

HB1xp67_ASAP7_75t_L g3631 ( 
.A(n_3299),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3388),
.Y(n_3632)
);

AND2x2_ASAP7_75t_L g3633 ( 
.A(n_3417),
.B(n_2491),
.Y(n_3633)
);

INVx2_ASAP7_75t_L g3634 ( 
.A(n_3294),
.Y(n_3634)
);

BUFx2_ASAP7_75t_L g3635 ( 
.A(n_3203),
.Y(n_3635)
);

OR2x2_ASAP7_75t_L g3636 ( 
.A(n_3391),
.B(n_2571),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_3418),
.B(n_2491),
.Y(n_3637)
);

OAI222xp33_ASAP7_75t_L g3638 ( 
.A1(n_3347),
.A2(n_2871),
.B1(n_3144),
.B2(n_3153),
.C1(n_3142),
.C2(n_3126),
.Y(n_3638)
);

INVx2_ASAP7_75t_L g3639 ( 
.A(n_3294),
.Y(n_3639)
);

AND2x2_ASAP7_75t_L g3640 ( 
.A(n_3424),
.B(n_2494),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_3403),
.B(n_2904),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3402),
.Y(n_3642)
);

OR2x2_ASAP7_75t_L g3643 ( 
.A(n_3328),
.B(n_2571),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3408),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3416),
.Y(n_3645)
);

AND2x2_ASAP7_75t_L g3646 ( 
.A(n_3414),
.B(n_2904),
.Y(n_3646)
);

AND2x2_ASAP7_75t_L g3647 ( 
.A(n_3457),
.B(n_3135),
.Y(n_3647)
);

AND2x4_ASAP7_75t_L g3648 ( 
.A(n_3371),
.B(n_2952),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3346),
.B(n_2825),
.Y(n_3649)
);

INVx4_ASAP7_75t_L g3650 ( 
.A(n_3368),
.Y(n_3650)
);

HB1xp67_ASAP7_75t_L g3651 ( 
.A(n_3219),
.Y(n_3651)
);

INVx2_ASAP7_75t_L g3652 ( 
.A(n_3402),
.Y(n_3652)
);

AND2x2_ASAP7_75t_L g3653 ( 
.A(n_3276),
.B(n_2825),
.Y(n_3653)
);

BUFx2_ASAP7_75t_L g3654 ( 
.A(n_3376),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3321),
.Y(n_3655)
);

HB1xp67_ASAP7_75t_L g3656 ( 
.A(n_3471),
.Y(n_3656)
);

OAI21xp5_ASAP7_75t_SL g3657 ( 
.A1(n_3468),
.A2(n_3136),
.B(n_3050),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3396),
.B(n_2588),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_3305),
.B(n_2582),
.Y(n_3659)
);

NOR2xp33_ASAP7_75t_SL g3660 ( 
.A(n_3493),
.B(n_3366),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3492),
.Y(n_3661)
);

AND2x2_ASAP7_75t_L g3662 ( 
.A(n_3517),
.B(n_3471),
.Y(n_3662)
);

AND2x4_ASAP7_75t_L g3663 ( 
.A(n_3538),
.B(n_3255),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3474),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3486),
.B(n_3229),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3625),
.B(n_3419),
.Y(n_3666)
);

BUFx2_ASAP7_75t_L g3667 ( 
.A(n_3489),
.Y(n_3667)
);

INVx2_ASAP7_75t_L g3668 ( 
.A(n_3478),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3532),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_3532),
.Y(n_3670)
);

AND2x2_ASAP7_75t_L g3671 ( 
.A(n_3504),
.B(n_3281),
.Y(n_3671)
);

HB1xp67_ASAP7_75t_L g3672 ( 
.A(n_3491),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3632),
.B(n_3459),
.Y(n_3673)
);

AND2x2_ASAP7_75t_L g3674 ( 
.A(n_3475),
.B(n_3281),
.Y(n_3674)
);

AND2x2_ASAP7_75t_L g3675 ( 
.A(n_3484),
.B(n_3455),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3483),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3485),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3501),
.Y(n_3678)
);

AND2x4_ASAP7_75t_L g3679 ( 
.A(n_3538),
.B(n_3255),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3507),
.Y(n_3680)
);

INVx2_ASAP7_75t_L g3681 ( 
.A(n_3479),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3644),
.B(n_3464),
.Y(n_3682)
);

OR2x2_ASAP7_75t_L g3683 ( 
.A(n_3566),
.B(n_3433),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3551),
.B(n_3455),
.Y(n_3684)
);

NAND3xp33_ASAP7_75t_L g3685 ( 
.A(n_3610),
.B(n_3266),
.C(n_3206),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3508),
.Y(n_3686)
);

AND2x2_ASAP7_75t_L g3687 ( 
.A(n_3505),
.B(n_3463),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3645),
.B(n_3311),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3509),
.Y(n_3689)
);

AND2x4_ASAP7_75t_L g3690 ( 
.A(n_3506),
.B(n_3289),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3480),
.Y(n_3691)
);

INVxp67_ASAP7_75t_SL g3692 ( 
.A(n_3533),
.Y(n_3692)
);

INVxp67_ASAP7_75t_SL g3693 ( 
.A(n_3533),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_SL g3694 ( 
.A(n_3495),
.B(n_3235),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3510),
.Y(n_3695)
);

NAND2x1p5_ASAP7_75t_L g3696 ( 
.A(n_3579),
.B(n_3210),
.Y(n_3696)
);

OR2x2_ASAP7_75t_L g3697 ( 
.A(n_3520),
.B(n_3516),
.Y(n_3697)
);

AND2x2_ASAP7_75t_L g3698 ( 
.A(n_3612),
.B(n_3463),
.Y(n_3698)
);

OR2x2_ASAP7_75t_L g3699 ( 
.A(n_3556),
.B(n_3236),
.Y(n_3699)
);

AND2x2_ASAP7_75t_L g3700 ( 
.A(n_3591),
.B(n_3413),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_3528),
.B(n_3413),
.Y(n_3701)
);

NOR3xp33_ASAP7_75t_L g3702 ( 
.A(n_3494),
.B(n_3288),
.C(n_3273),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3481),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3513),
.Y(n_3704)
);

INVxp67_ASAP7_75t_SL g3705 ( 
.A(n_3534),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3536),
.B(n_3305),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_SL g3707 ( 
.A(n_3515),
.B(n_3454),
.Y(n_3707)
);

AND2x2_ASAP7_75t_L g3708 ( 
.A(n_3602),
.B(n_3231),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3521),
.Y(n_3709)
);

AND2x2_ASAP7_75t_L g3710 ( 
.A(n_3603),
.B(n_3404),
.Y(n_3710)
);

OAI21xp5_ASAP7_75t_SL g3711 ( 
.A1(n_3624),
.A2(n_3272),
.B(n_3261),
.Y(n_3711)
);

OR2x2_ASAP7_75t_L g3712 ( 
.A(n_3488),
.B(n_3426),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3526),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3547),
.B(n_3450),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3628),
.B(n_3301),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3529),
.Y(n_3716)
);

NAND3xp33_ASAP7_75t_L g3717 ( 
.A(n_3610),
.B(n_3334),
.C(n_3184),
.Y(n_3717)
);

OR2x2_ASAP7_75t_L g3718 ( 
.A(n_3514),
.B(n_3426),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3502),
.B(n_3450),
.Y(n_3719)
);

AND2x4_ASAP7_75t_L g3720 ( 
.A(n_3506),
.B(n_3523),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3628),
.B(n_3569),
.Y(n_3721)
);

HB1xp67_ASAP7_75t_L g3722 ( 
.A(n_3651),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3530),
.Y(n_3723)
);

HB1xp67_ASAP7_75t_L g3724 ( 
.A(n_3527),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3531),
.Y(n_3725)
);

INVx2_ASAP7_75t_L g3726 ( 
.A(n_3482),
.Y(n_3726)
);

HB1xp67_ASAP7_75t_L g3727 ( 
.A(n_3527),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3569),
.B(n_3246),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3571),
.B(n_3246),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3571),
.B(n_3246),
.Y(n_3730)
);

AND2x4_ASAP7_75t_L g3731 ( 
.A(n_3523),
.B(n_3289),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3522),
.B(n_3369),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3541),
.Y(n_3733)
);

HB1xp67_ASAP7_75t_L g3734 ( 
.A(n_3477),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3595),
.B(n_3395),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3546),
.Y(n_3736)
);

HB1xp67_ASAP7_75t_L g3737 ( 
.A(n_3534),
.Y(n_3737)
);

NAND2x1_ASAP7_75t_SL g3738 ( 
.A(n_3631),
.B(n_3286),
.Y(n_3738)
);

AND2x4_ASAP7_75t_SL g3739 ( 
.A(n_3570),
.B(n_3377),
.Y(n_3739)
);

NOR2xp33_ASAP7_75t_L g3740 ( 
.A(n_3618),
.B(n_3314),
.Y(n_3740)
);

HB1xp67_ASAP7_75t_L g3741 ( 
.A(n_3656),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_3544),
.B(n_3187),
.Y(n_3742)
);

AND2x2_ASAP7_75t_L g3743 ( 
.A(n_3487),
.B(n_3197),
.Y(n_3743)
);

NOR2xp67_ASAP7_75t_L g3744 ( 
.A(n_3585),
.B(n_3427),
.Y(n_3744)
);

OR2x2_ASAP7_75t_L g3745 ( 
.A(n_3525),
.B(n_3426),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3548),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3605),
.B(n_3283),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3550),
.Y(n_3748)
);

OR2x2_ASAP7_75t_L g3749 ( 
.A(n_3535),
.B(n_3322),
.Y(n_3749)
);

INVx4_ASAP7_75t_L g3750 ( 
.A(n_3581),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3553),
.Y(n_3751)
);

NAND2x1_ASAP7_75t_L g3752 ( 
.A(n_3581),
.B(n_3320),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3490),
.Y(n_3753)
);

OR2x2_ASAP7_75t_L g3754 ( 
.A(n_3543),
.B(n_3320),
.Y(n_3754)
);

AND2x4_ASAP7_75t_L g3755 ( 
.A(n_3587),
.B(n_3368),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3555),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3498),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3664),
.Y(n_3758)
);

AND2x2_ASAP7_75t_L g3759 ( 
.A(n_3661),
.B(n_3721),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3676),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3668),
.Y(n_3761)
);

BUFx2_ASAP7_75t_L g3762 ( 
.A(n_3738),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_3721),
.B(n_3646),
.Y(n_3763)
);

OR2x2_ASAP7_75t_L g3764 ( 
.A(n_3697),
.B(n_3575),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3669),
.B(n_3606),
.Y(n_3765)
);

INVx2_ASAP7_75t_SL g3766 ( 
.A(n_3750),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3677),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3678),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3681),
.Y(n_3769)
);

AND2x2_ASAP7_75t_L g3770 ( 
.A(n_3670),
.B(n_3641),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3680),
.Y(n_3771)
);

INVx2_ASAP7_75t_SL g3772 ( 
.A(n_3750),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3691),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3715),
.B(n_3586),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3715),
.B(n_3622),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_3734),
.B(n_3653),
.Y(n_3776)
);

AND2x2_ASAP7_75t_L g3777 ( 
.A(n_3720),
.B(n_3719),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3720),
.B(n_3575),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3662),
.B(n_3574),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3686),
.Y(n_3780)
);

HB1xp67_ASAP7_75t_L g3781 ( 
.A(n_3722),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3724),
.B(n_3607),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3727),
.B(n_3647),
.Y(n_3783)
);

AND2x2_ASAP7_75t_L g3784 ( 
.A(n_3703),
.B(n_3617),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3726),
.B(n_3636),
.Y(n_3785)
);

AND2x2_ASAP7_75t_L g3786 ( 
.A(n_3753),
.B(n_3633),
.Y(n_3786)
);

AND2x2_ASAP7_75t_L g3787 ( 
.A(n_3757),
.B(n_3637),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3689),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3688),
.B(n_3655),
.Y(n_3789)
);

AND2x2_ASAP7_75t_L g3790 ( 
.A(n_3695),
.B(n_3640),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3704),
.B(n_3627),
.Y(n_3791)
);

AND2x2_ASAP7_75t_L g3792 ( 
.A(n_3709),
.B(n_3634),
.Y(n_3792)
);

AND2x2_ASAP7_75t_L g3793 ( 
.A(n_3713),
.B(n_3639),
.Y(n_3793)
);

OR2x2_ASAP7_75t_L g3794 ( 
.A(n_3672),
.B(n_3718),
.Y(n_3794)
);

INVx2_ASAP7_75t_L g3795 ( 
.A(n_3716),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_SL g3796 ( 
.A(n_3660),
.B(n_3624),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_3756),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3723),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3725),
.Y(n_3799)
);

BUFx2_ASAP7_75t_L g3800 ( 
.A(n_3667),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3733),
.B(n_3642),
.Y(n_3801)
);

INVxp67_ASAP7_75t_SL g3802 ( 
.A(n_3737),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3688),
.B(n_3582),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3736),
.Y(n_3804)
);

AND2x2_ASAP7_75t_L g3805 ( 
.A(n_3746),
.B(n_3652),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3748),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3747),
.B(n_3583),
.Y(n_3807)
);

INVx1_ASAP7_75t_SL g3808 ( 
.A(n_3739),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3751),
.B(n_3614),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3747),
.B(n_3598),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3741),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3745),
.Y(n_3812)
);

AND2x2_ASAP7_75t_L g3813 ( 
.A(n_3666),
.B(n_3620),
.Y(n_3813)
);

AND2x2_ASAP7_75t_L g3814 ( 
.A(n_3666),
.B(n_3621),
.Y(n_3814)
);

AND2x2_ASAP7_75t_L g3815 ( 
.A(n_3673),
.B(n_3626),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3712),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3673),
.B(n_3560),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3708),
.B(n_3561),
.Y(n_3818)
);

INVx2_ASAP7_75t_L g3819 ( 
.A(n_3682),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3699),
.Y(n_3820)
);

AND2x4_ASAP7_75t_L g3821 ( 
.A(n_3744),
.B(n_3587),
.Y(n_3821)
);

AND2x2_ASAP7_75t_L g3822 ( 
.A(n_3682),
.B(n_3557),
.Y(n_3822)
);

AND2x2_ASAP7_75t_L g3823 ( 
.A(n_3714),
.B(n_3572),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3665),
.B(n_3593),
.Y(n_3824)
);

NAND2x1_ASAP7_75t_L g3825 ( 
.A(n_3690),
.B(n_3635),
.Y(n_3825)
);

OR2x2_ASAP7_75t_L g3826 ( 
.A(n_3728),
.B(n_3545),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3728),
.Y(n_3827)
);

OR2x2_ASAP7_75t_L g3828 ( 
.A(n_3700),
.B(n_3596),
.Y(n_3828)
);

AND2x4_ASAP7_75t_L g3829 ( 
.A(n_3744),
.B(n_3630),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3710),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3742),
.B(n_3597),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3692),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3812),
.Y(n_3833)
);

OAI22xp33_ASAP7_75t_L g3834 ( 
.A1(n_3825),
.A2(n_3660),
.B1(n_3711),
.B2(n_3685),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3827),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3778),
.B(n_3763),
.Y(n_3836)
);

NAND2x2_ASAP7_75t_L g3837 ( 
.A(n_3766),
.B(n_3752),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3800),
.Y(n_3838)
);

INVx2_ASAP7_75t_L g3839 ( 
.A(n_3794),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3827),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3778),
.B(n_3684),
.Y(n_3841)
);

OR2x6_ASAP7_75t_L g3842 ( 
.A(n_3796),
.B(n_3696),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3794),
.Y(n_3843)
);

AND2x4_ASAP7_75t_L g3844 ( 
.A(n_3766),
.B(n_3693),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3759),
.Y(n_3845)
);

INVx2_ASAP7_75t_SL g3846 ( 
.A(n_3808),
.Y(n_3846)
);

AND2x2_ASAP7_75t_L g3847 ( 
.A(n_3763),
.B(n_3698),
.Y(n_3847)
);

NAND2xp33_ASAP7_75t_SL g3848 ( 
.A(n_3796),
.B(n_3205),
.Y(n_3848)
);

AND2x2_ASAP7_75t_L g3849 ( 
.A(n_3776),
.B(n_3675),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_3819),
.B(n_3600),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3781),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3776),
.B(n_3777),
.Y(n_3852)
);

A2O1A1Ixp33_ASAP7_75t_L g3853 ( 
.A1(n_3772),
.A2(n_3711),
.B(n_3685),
.C(n_3702),
.Y(n_3853)
);

OA222x2_ASAP7_75t_L g3854 ( 
.A1(n_3764),
.A2(n_3683),
.B1(n_3565),
.B2(n_3524),
.C1(n_3754),
.C2(n_3749),
.Y(n_3854)
);

INVx2_ASAP7_75t_SL g3855 ( 
.A(n_3772),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3759),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3819),
.B(n_3729),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3795),
.Y(n_3858)
);

AOI22xp5_ASAP7_75t_L g3859 ( 
.A1(n_3820),
.A2(n_3717),
.B1(n_3588),
.B2(n_3503),
.Y(n_3859)
);

OAI322xp33_ASAP7_75t_L g3860 ( 
.A1(n_3826),
.A2(n_3707),
.A3(n_3503),
.B1(n_3717),
.B2(n_3588),
.C1(n_3740),
.C2(n_3694),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3777),
.B(n_3674),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3822),
.B(n_3729),
.Y(n_3862)
);

INVxp67_ASAP7_75t_L g3863 ( 
.A(n_3802),
.Y(n_3863)
);

OAI22xp33_ASAP7_75t_SL g3864 ( 
.A1(n_3762),
.A2(n_3705),
.B1(n_3731),
.B2(n_3690),
.Y(n_3864)
);

INVx2_ASAP7_75t_L g3865 ( 
.A(n_3758),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3822),
.B(n_3671),
.Y(n_3866)
);

AOI22xp5_ASAP7_75t_L g3867 ( 
.A1(n_3783),
.A2(n_3476),
.B1(n_3590),
.B2(n_3562),
.Y(n_3867)
);

INVx2_ASAP7_75t_L g3868 ( 
.A(n_3758),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_3761),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3816),
.Y(n_3870)
);

O2A1O1Ixp33_ASAP7_75t_L g3871 ( 
.A1(n_3774),
.A2(n_3775),
.B(n_3336),
.C(n_3609),
.Y(n_3871)
);

OR2x2_ASAP7_75t_L g3872 ( 
.A(n_3826),
.B(n_3730),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3761),
.Y(n_3873)
);

NAND4xp75_ASAP7_75t_L g3874 ( 
.A(n_3782),
.B(n_3202),
.C(n_3562),
.D(n_3580),
.Y(n_3874)
);

CKINVDCx16_ASAP7_75t_R g3875 ( 
.A(n_3783),
.Y(n_3875)
);

OAI322xp33_ASAP7_75t_L g3876 ( 
.A1(n_3817),
.A2(n_3609),
.A3(n_3274),
.B1(n_3584),
.B2(n_3552),
.C1(n_3643),
.C2(n_3601),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3770),
.B(n_3730),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3795),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3770),
.B(n_3813),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3797),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3797),
.Y(n_3881)
);

INVx3_ASAP7_75t_L g3882 ( 
.A(n_3821),
.Y(n_3882)
);

OAI22xp5_ASAP7_75t_L g3883 ( 
.A1(n_3831),
.A2(n_3731),
.B1(n_3679),
.B2(n_3663),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3813),
.B(n_3814),
.Y(n_3884)
);

OR2x2_ASAP7_75t_L g3885 ( 
.A(n_3814),
.B(n_3701),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3815),
.B(n_3615),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_3815),
.B(n_3616),
.Y(n_3887)
);

XNOR2x1_ASAP7_75t_L g3888 ( 
.A(n_3830),
.B(n_3240),
.Y(n_3888)
);

NOR2x1_ASAP7_75t_L g3889 ( 
.A(n_3821),
.B(n_3542),
.Y(n_3889)
);

INVx2_ASAP7_75t_SL g3890 ( 
.A(n_3828),
.Y(n_3890)
);

AND2x2_ASAP7_75t_L g3891 ( 
.A(n_3823),
.B(n_3687),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3760),
.Y(n_3892)
);

NAND2x1p5_ASAP7_75t_L g3893 ( 
.A(n_3832),
.B(n_3542),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3769),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3769),
.Y(n_3895)
);

INVx2_ASAP7_75t_L g3896 ( 
.A(n_3773),
.Y(n_3896)
);

OR2x2_ASAP7_75t_L g3897 ( 
.A(n_3765),
.B(n_3706),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3773),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3782),
.Y(n_3899)
);

NOR3xp33_ASAP7_75t_L g3900 ( 
.A(n_3834),
.B(n_3214),
.C(n_3500),
.Y(n_3900)
);

NOR4xp25_ASAP7_75t_SL g3901 ( 
.A(n_3848),
.B(n_3275),
.C(n_3285),
.D(n_3518),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3850),
.Y(n_3902)
);

AOI31xp33_ASAP7_75t_L g3903 ( 
.A1(n_3853),
.A2(n_3223),
.A3(n_3226),
.B(n_3663),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3870),
.Y(n_3904)
);

INVx2_ASAP7_75t_L g3905 ( 
.A(n_3844),
.Y(n_3905)
);

AOI21xp5_ASAP7_75t_L g3906 ( 
.A1(n_3864),
.A2(n_3821),
.B(n_3829),
.Y(n_3906)
);

A2O1A1Ixp33_ASAP7_75t_L g3907 ( 
.A1(n_3871),
.A2(n_3679),
.B(n_3829),
.C(n_3392),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3870),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3884),
.Y(n_3909)
);

INVx2_ASAP7_75t_SL g3910 ( 
.A(n_3844),
.Y(n_3910)
);

AOI22xp33_ASAP7_75t_L g3911 ( 
.A1(n_3860),
.A2(n_3500),
.B1(n_3623),
.B2(n_3563),
.Y(n_3911)
);

NOR2xp33_ASAP7_75t_L g3912 ( 
.A(n_3846),
.B(n_3327),
.Y(n_3912)
);

AND2x2_ASAP7_75t_L g3913 ( 
.A(n_3875),
.B(n_3779),
.Y(n_3913)
);

OAI221xp5_ASAP7_75t_SL g3914 ( 
.A1(n_3859),
.A2(n_3241),
.B1(n_3657),
.B2(n_3511),
.C(n_3577),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3845),
.Y(n_3915)
);

OAI21xp5_ASAP7_75t_L g3916 ( 
.A1(n_3842),
.A2(n_3519),
.B(n_3613),
.Y(n_3916)
);

OAI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3842),
.A2(n_3519),
.B(n_3613),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3856),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3890),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_3867),
.B(n_3790),
.Y(n_3920)
);

AOI21xp33_ASAP7_75t_L g3921 ( 
.A1(n_3883),
.A2(n_3619),
.B(n_3604),
.Y(n_3921)
);

AOI31xp33_ASAP7_75t_L g3922 ( 
.A1(n_3889),
.A2(n_3570),
.A3(n_3381),
.B(n_3428),
.Y(n_3922)
);

OAI21xp33_ASAP7_75t_L g3923 ( 
.A1(n_3838),
.A2(n_3789),
.B(n_3803),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3865),
.Y(n_3924)
);

INVx2_ASAP7_75t_L g3925 ( 
.A(n_3868),
.Y(n_3925)
);

OAI21xp5_ASAP7_75t_L g3926 ( 
.A1(n_3863),
.A2(n_3811),
.B(n_3657),
.Y(n_3926)
);

OR2x2_ASAP7_75t_L g3927 ( 
.A(n_3872),
.B(n_3824),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3833),
.Y(n_3928)
);

XOR2xp5_ASAP7_75t_L g3929 ( 
.A(n_3888),
.B(n_3213),
.Y(n_3929)
);

AOI31xp33_ASAP7_75t_L g3930 ( 
.A1(n_3893),
.A2(n_3420),
.A3(n_3430),
.B(n_3183),
.Y(n_3930)
);

O2A1O1Ixp33_ASAP7_75t_SL g3931 ( 
.A1(n_3854),
.A2(n_3383),
.B(n_3558),
.C(n_3466),
.Y(n_3931)
);

INVx2_ASAP7_75t_L g3932 ( 
.A(n_3869),
.Y(n_3932)
);

INVxp67_ASAP7_75t_L g3933 ( 
.A(n_3851),
.Y(n_3933)
);

OAI21xp33_ASAP7_75t_L g3934 ( 
.A1(n_3862),
.A2(n_3807),
.B(n_3810),
.Y(n_3934)
);

INVx1_ASAP7_75t_SL g3935 ( 
.A(n_3855),
.Y(n_3935)
);

AOI21xp33_ASAP7_75t_L g3936 ( 
.A1(n_3892),
.A2(n_3325),
.B(n_3577),
.Y(n_3936)
);

OAI21xp5_ASAP7_75t_L g3937 ( 
.A1(n_3874),
.A2(n_3499),
.B(n_3461),
.Y(n_3937)
);

OR2x2_ASAP7_75t_L g3938 ( 
.A(n_3877),
.B(n_3818),
.Y(n_3938)
);

HB1xp67_ASAP7_75t_L g3939 ( 
.A(n_3839),
.Y(n_3939)
);

OAI22xp33_ASAP7_75t_SL g3940 ( 
.A1(n_3837),
.A2(n_3524),
.B1(n_3565),
.B2(n_3829),
.Y(n_3940)
);

OAI22xp33_ASAP7_75t_L g3941 ( 
.A1(n_3882),
.A2(n_3885),
.B1(n_3897),
.B2(n_3879),
.Y(n_3941)
);

INVx2_ASAP7_75t_L g3942 ( 
.A(n_3873),
.Y(n_3942)
);

AOI22xp5_ASAP7_75t_L g3943 ( 
.A1(n_3900),
.A2(n_3511),
.B1(n_3568),
.B2(n_3442),
.Y(n_3943)
);

NOR2xp33_ASAP7_75t_L g3944 ( 
.A(n_3903),
.B(n_3318),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3902),
.Y(n_3945)
);

AOI211xp5_ASAP7_75t_L g3946 ( 
.A1(n_3931),
.A2(n_3876),
.B(n_3215),
.C(n_3228),
.Y(n_3946)
);

INVx1_ASAP7_75t_SL g3947 ( 
.A(n_3935),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3909),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3904),
.Y(n_3949)
);

AND2x2_ASAP7_75t_L g3950 ( 
.A(n_3910),
.B(n_3882),
.Y(n_3950)
);

NOR2xp33_ASAP7_75t_L g3951 ( 
.A(n_3903),
.B(n_3233),
.Y(n_3951)
);

OR2x2_ASAP7_75t_L g3952 ( 
.A(n_3938),
.B(n_3857),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3924),
.Y(n_3953)
);

O2A1O1Ixp33_ASAP7_75t_L g3954 ( 
.A1(n_3914),
.A2(n_3190),
.B(n_3360),
.C(n_3337),
.Y(n_3954)
);

NAND3xp33_ASAP7_75t_SL g3955 ( 
.A(n_3901),
.B(n_3307),
.C(n_3304),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3908),
.Y(n_3956)
);

AOI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3911),
.A2(n_3843),
.B1(n_3833),
.B2(n_3790),
.Y(n_3957)
);

OAI221xp5_ASAP7_75t_L g3958 ( 
.A1(n_3907),
.A2(n_3341),
.B1(n_3887),
.B2(n_3886),
.C(n_3899),
.Y(n_3958)
);

NAND2x1_ASAP7_75t_L g3959 ( 
.A(n_3922),
.B(n_3852),
.Y(n_3959)
);

OR2x2_ASAP7_75t_L g3960 ( 
.A(n_3927),
.B(n_3915),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_3925),
.Y(n_3961)
);

OAI22xp33_ASAP7_75t_L g3962 ( 
.A1(n_3922),
.A2(n_3524),
.B1(n_3565),
.B2(n_3654),
.Y(n_3962)
);

AND2x2_ASAP7_75t_L g3963 ( 
.A(n_3935),
.B(n_3836),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3934),
.B(n_3847),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_3920),
.B(n_3926),
.Y(n_3965)
);

INVx3_ASAP7_75t_L g3966 ( 
.A(n_3905),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3932),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_L g3968 ( 
.A(n_3923),
.B(n_3866),
.Y(n_3968)
);

NOR2xp67_ASAP7_75t_SL g3969 ( 
.A(n_3906),
.B(n_3258),
.Y(n_3969)
);

AOI22xp5_ASAP7_75t_L g3970 ( 
.A1(n_3937),
.A2(n_3465),
.B1(n_3472),
.B2(n_3497),
.Y(n_3970)
);

OAI22xp5_ASAP7_75t_L g3971 ( 
.A1(n_3941),
.A2(n_3849),
.B1(n_3891),
.B2(n_3841),
.Y(n_3971)
);

OAI21xp5_ASAP7_75t_L g3972 ( 
.A1(n_3916),
.A2(n_3917),
.B(n_3930),
.Y(n_3972)
);

OAI211xp5_ASAP7_75t_L g3973 ( 
.A1(n_3901),
.A2(n_3316),
.B(n_3330),
.C(n_3382),
.Y(n_3973)
);

OAI22xp5_ASAP7_75t_L g3974 ( 
.A1(n_3913),
.A2(n_3861),
.B1(n_3779),
.B2(n_3743),
.Y(n_3974)
);

OAI21xp5_ASAP7_75t_L g3975 ( 
.A1(n_3930),
.A2(n_3940),
.B(n_3936),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_L g3976 ( 
.A(n_3918),
.B(n_3823),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3919),
.B(n_3765),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3928),
.B(n_3767),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3933),
.B(n_3768),
.Y(n_3979)
);

OAI221xp5_ASAP7_75t_L g3980 ( 
.A1(n_3921),
.A2(n_3194),
.B1(n_3780),
.B2(n_3788),
.C(n_3771),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3939),
.Y(n_3981)
);

AND2x2_ASAP7_75t_L g3982 ( 
.A(n_3942),
.B(n_3784),
.Y(n_3982)
);

OAI22xp33_ASAP7_75t_L g3983 ( 
.A1(n_3912),
.A2(n_3390),
.B1(n_3895),
.B2(n_3894),
.Y(n_3983)
);

CKINVDCx16_ASAP7_75t_R g3984 ( 
.A(n_3929),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3902),
.Y(n_3985)
);

O2A1O1Ixp5_ASAP7_75t_L g3986 ( 
.A1(n_3907),
.A2(n_3799),
.B(n_3804),
.C(n_3798),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3902),
.Y(n_3987)
);

AOI21xp33_ASAP7_75t_L g3988 ( 
.A1(n_3903),
.A2(n_3361),
.B(n_3348),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3911),
.B(n_3806),
.Y(n_3989)
);

AND2x2_ASAP7_75t_L g3990 ( 
.A(n_3947),
.B(n_3784),
.Y(n_3990)
);

INVx2_ASAP7_75t_L g3991 ( 
.A(n_3963),
.Y(n_3991)
);

NOR2xp33_ASAP7_75t_L g3992 ( 
.A(n_3984),
.B(n_3271),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3960),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3943),
.B(n_3835),
.Y(n_3994)
);

AOI221xp5_ASAP7_75t_SL g3995 ( 
.A1(n_3972),
.A2(n_3962),
.B1(n_3975),
.B2(n_3954),
.C(n_3965),
.Y(n_3995)
);

OR3x1_ASAP7_75t_L g3996 ( 
.A(n_3955),
.B(n_3499),
.C(n_3280),
.Y(n_3996)
);

AND2x2_ASAP7_75t_L g3997 ( 
.A(n_3959),
.B(n_3786),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3950),
.B(n_3786),
.Y(n_3998)
);

NOR2xp33_ASAP7_75t_L g3999 ( 
.A(n_3944),
.B(n_3312),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3978),
.Y(n_4000)
);

NAND3xp33_ASAP7_75t_SL g4001 ( 
.A(n_3986),
.B(n_3946),
.C(n_3943),
.Y(n_4001)
);

INVx3_ASAP7_75t_L g4002 ( 
.A(n_3966),
.Y(n_4002)
);

AOI221xp5_ASAP7_75t_L g4003 ( 
.A1(n_3969),
.A2(n_3840),
.B1(n_3835),
.B2(n_3878),
.C(n_3858),
.Y(n_4003)
);

NOR2xp33_ASAP7_75t_L g4004 ( 
.A(n_3951),
.B(n_3326),
.Y(n_4004)
);

NAND3xp33_ASAP7_75t_L g4005 ( 
.A(n_3957),
.B(n_3280),
.C(n_3030),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3979),
.Y(n_4006)
);

NOR3xp33_ASAP7_75t_L g4007 ( 
.A(n_3973),
.B(n_3234),
.C(n_3217),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3981),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_SL g4009 ( 
.A(n_3971),
.B(n_3840),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3989),
.B(n_3948),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_3945),
.B(n_3791),
.Y(n_4011)
);

INVx2_ASAP7_75t_L g4012 ( 
.A(n_3966),
.Y(n_4012)
);

AOI21xp5_ASAP7_75t_L g4013 ( 
.A1(n_3988),
.A2(n_3362),
.B(n_3441),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3985),
.B(n_3791),
.Y(n_4014)
);

OA22x2_ASAP7_75t_L g4015 ( 
.A1(n_3970),
.A2(n_3441),
.B1(n_3735),
.B2(n_3611),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3987),
.B(n_3792),
.Y(n_4016)
);

OAI21xp5_ASAP7_75t_L g4017 ( 
.A1(n_3970),
.A2(n_3958),
.B(n_3983),
.Y(n_4017)
);

NAND3xp33_ASAP7_75t_L g4018 ( 
.A(n_3949),
.B(n_3956),
.C(n_3980),
.Y(n_4018)
);

NAND3xp33_ASAP7_75t_L g4019 ( 
.A(n_3964),
.B(n_3968),
.C(n_3961),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3977),
.B(n_3787),
.Y(n_4020)
);

AOI21xp5_ASAP7_75t_L g4021 ( 
.A1(n_4001),
.A2(n_3974),
.B(n_3967),
.Y(n_4021)
);

AOI21xp5_ASAP7_75t_L g4022 ( 
.A1(n_3992),
.A2(n_3953),
.B(n_3976),
.Y(n_4022)
);

AOI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_4004),
.A2(n_3952),
.B(n_3982),
.Y(n_4023)
);

NOR3xp33_ASAP7_75t_L g4024 ( 
.A(n_3995),
.B(n_2568),
.C(n_3467),
.Y(n_4024)
);

AOI22xp33_ASAP7_75t_L g4025 ( 
.A1(n_4015),
.A2(n_3630),
.B1(n_3755),
.B2(n_3554),
.Y(n_4025)
);

AND2x2_ASAP7_75t_L g4026 ( 
.A(n_3997),
.B(n_3787),
.Y(n_4026)
);

AOI22xp33_ASAP7_75t_SL g4027 ( 
.A1(n_4017),
.A2(n_3451),
.B1(n_3340),
.B2(n_3594),
.Y(n_4027)
);

AOI21xp5_ASAP7_75t_SL g4028 ( 
.A1(n_4003),
.A2(n_3345),
.B(n_3085),
.Y(n_4028)
);

AOI211xp5_ASAP7_75t_L g4029 ( 
.A1(n_4007),
.A2(n_3332),
.B(n_3648),
.C(n_3185),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_SL g4030 ( 
.A(n_4002),
.B(n_3894),
.Y(n_4030)
);

NOR3xp33_ASAP7_75t_L g4031 ( 
.A(n_4005),
.B(n_3088),
.C(n_3010),
.Y(n_4031)
);

NOR2xp67_ASAP7_75t_L g4032 ( 
.A(n_4019),
.B(n_703),
.Y(n_4032)
);

AOI211x1_ASAP7_75t_L g4033 ( 
.A1(n_4018),
.A2(n_3878),
.B(n_3881),
.C(n_3880),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_4006),
.B(n_3898),
.Y(n_4034)
);

AOI22xp33_ASAP7_75t_SL g4035 ( 
.A1(n_4005),
.A2(n_3185),
.B1(n_3648),
.B2(n_3393),
.Y(n_4035)
);

NOR3xp33_ASAP7_75t_L g4036 ( 
.A(n_4018),
.B(n_3089),
.C(n_2842),
.Y(n_4036)
);

AOI21xp5_ASAP7_75t_L g4037 ( 
.A1(n_3999),
.A2(n_3608),
.B(n_3599),
.Y(n_4037)
);

NAND3xp33_ASAP7_75t_L g4038 ( 
.A(n_4019),
.B(n_3400),
.C(n_3309),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3990),
.Y(n_4039)
);

NOR2xp67_ASAP7_75t_SL g4040 ( 
.A(n_4013),
.B(n_4002),
.Y(n_4040)
);

AND3x1_ASAP7_75t_L g4041 ( 
.A(n_4010),
.B(n_3611),
.C(n_2852),
.Y(n_4041)
);

INVxp67_ASAP7_75t_L g4042 ( 
.A(n_4008),
.Y(n_4042)
);

AND2x2_ASAP7_75t_L g4043 ( 
.A(n_3991),
.B(n_3785),
.Y(n_4043)
);

NOR3xp33_ASAP7_75t_L g4044 ( 
.A(n_4009),
.B(n_2665),
.C(n_2655),
.Y(n_4044)
);

OR3x1_ASAP7_75t_L g4045 ( 
.A(n_4039),
.B(n_3993),
.C(n_3996),
.Y(n_4045)
);

OAI221xp5_ASAP7_75t_L g4046 ( 
.A1(n_4027),
.A2(n_4035),
.B1(n_4024),
.B2(n_4040),
.C(n_4021),
.Y(n_4046)
);

NOR3xp33_ASAP7_75t_SL g4047 ( 
.A(n_4038),
.B(n_3994),
.C(n_4000),
.Y(n_4047)
);

AOI22xp33_ASAP7_75t_L g4048 ( 
.A1(n_4035),
.A2(n_4012),
.B1(n_4014),
.B2(n_4011),
.Y(n_4048)
);

AOI22xp5_ASAP7_75t_L g4049 ( 
.A1(n_4041),
.A2(n_3998),
.B1(n_4016),
.B2(n_4020),
.Y(n_4049)
);

NOR3xp33_ASAP7_75t_L g4050 ( 
.A(n_4032),
.B(n_2732),
.C(n_2760),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_4022),
.B(n_3895),
.Y(n_4051)
);

OAI31xp33_ASAP7_75t_L g4052 ( 
.A1(n_4042),
.A2(n_3649),
.A3(n_3638),
.B(n_2913),
.Y(n_4052)
);

AOI211xp5_ASAP7_75t_L g4053 ( 
.A1(n_4028),
.A2(n_3375),
.B(n_3638),
.C(n_3629),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_4034),
.Y(n_4054)
);

NAND3xp33_ASAP7_75t_L g4055 ( 
.A(n_4033),
.B(n_3041),
.C(n_3306),
.Y(n_4055)
);

BUFx2_ASAP7_75t_L g4056 ( 
.A(n_4043),
.Y(n_4056)
);

NOR2xp33_ASAP7_75t_L g4057 ( 
.A(n_4023),
.B(n_3898),
.Y(n_4057)
);

AOI211xp5_ASAP7_75t_L g4058 ( 
.A1(n_4036),
.A2(n_3496),
.B(n_3658),
.C(n_3512),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_SL g4059 ( 
.A(n_4029),
.B(n_3896),
.Y(n_4059)
);

O2A1O1Ixp33_ASAP7_75t_L g4060 ( 
.A1(n_4031),
.A2(n_2913),
.B(n_2868),
.C(n_3438),
.Y(n_4060)
);

NOR3xp33_ASAP7_75t_L g4061 ( 
.A(n_4044),
.B(n_4030),
.C(n_4037),
.Y(n_4061)
);

NAND2xp33_ASAP7_75t_R g4062 ( 
.A(n_4026),
.B(n_3384),
.Y(n_4062)
);

AOI221xp5_ASAP7_75t_L g4063 ( 
.A1(n_4025),
.A2(n_3539),
.B1(n_3512),
.B2(n_3559),
.C(n_3567),
.Y(n_4063)
);

OAI221xp5_ASAP7_75t_L g4064 ( 
.A1(n_4027),
.A2(n_3658),
.B1(n_3469),
.B2(n_3370),
.C(n_3310),
.Y(n_4064)
);

AO22x2_ASAP7_75t_L g4065 ( 
.A1(n_4054),
.A2(n_3650),
.B1(n_3537),
.B2(n_3732),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_4056),
.Y(n_4066)
);

AOI22xp5_ASAP7_75t_L g4067 ( 
.A1(n_4046),
.A2(n_3659),
.B1(n_3329),
.B2(n_3755),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_4051),
.Y(n_4068)
);

NOR2xp33_ASAP7_75t_L g4069 ( 
.A(n_4057),
.B(n_3539),
.Y(n_4069)
);

NOR2x1_ASAP7_75t_SL g4070 ( 
.A(n_4059),
.B(n_3438),
.Y(n_4070)
);

AND3x1_ASAP7_75t_L g4071 ( 
.A(n_4047),
.B(n_3540),
.C(n_3578),
.Y(n_4071)
);

NOR2x1_ASAP7_75t_L g4072 ( 
.A(n_4045),
.B(n_2460),
.Y(n_4072)
);

AOI22xp5_ASAP7_75t_L g4073 ( 
.A1(n_4053),
.A2(n_3554),
.B1(n_3549),
.B2(n_3785),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_4055),
.B(n_3809),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_4061),
.B(n_3809),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_4050),
.Y(n_4076)
);

AND2x4_ASAP7_75t_L g4077 ( 
.A(n_4049),
.B(n_3792),
.Y(n_4077)
);

AO22x2_ASAP7_75t_L g4078 ( 
.A1(n_4048),
.A2(n_3650),
.B1(n_3374),
.B2(n_3573),
.Y(n_4078)
);

NAND4xp75_ASAP7_75t_L g4079 ( 
.A(n_4072),
.B(n_4052),
.C(n_4063),
.D(n_4058),
.Y(n_4079)
);

AOI211xp5_ASAP7_75t_L g4080 ( 
.A1(n_4066),
.A2(n_4064),
.B(n_4060),
.C(n_4062),
.Y(n_4080)
);

OR2x2_ASAP7_75t_L g4081 ( 
.A(n_4075),
.B(n_3793),
.Y(n_4081)
);

AND2x2_ASAP7_75t_L g4082 ( 
.A(n_4070),
.B(n_3793),
.Y(n_4082)
);

AND3x2_ASAP7_75t_L g4083 ( 
.A(n_4076),
.B(n_3374),
.C(n_3175),
.Y(n_4083)
);

NOR3xp33_ASAP7_75t_L g4084 ( 
.A(n_4068),
.B(n_2776),
.C(n_2605),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_4071),
.B(n_3801),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_4074),
.Y(n_4086)
);

AOI221xp5_ASAP7_75t_L g4087 ( 
.A1(n_4067),
.A2(n_3564),
.B1(n_3589),
.B2(n_3576),
.C(n_3592),
.Y(n_4087)
);

NAND2xp5_ASAP7_75t_L g4088 ( 
.A(n_4069),
.B(n_3801),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_4077),
.B(n_3805),
.Y(n_4089)
);

XOR2x2_ASAP7_75t_L g4090 ( 
.A(n_4073),
.B(n_3425),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4081),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_4086),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_4083),
.Y(n_4093)
);

HB1xp67_ASAP7_75t_L g4094 ( 
.A(n_4080),
.Y(n_4094)
);

INVx1_ASAP7_75t_SL g4095 ( 
.A(n_4090),
.Y(n_4095)
);

HB1xp67_ASAP7_75t_L g4096 ( 
.A(n_4079),
.Y(n_4096)
);

BUFx2_ASAP7_75t_L g4097 ( 
.A(n_4082),
.Y(n_4097)
);

CKINVDCx5p33_ASAP7_75t_R g4098 ( 
.A(n_4085),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_4097),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_4096),
.B(n_4078),
.Y(n_4100)
);

AOI211xp5_ASAP7_75t_SL g4101 ( 
.A1(n_4094),
.A2(n_4087),
.B(n_4089),
.C(n_4088),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_4099),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_4100),
.B(n_4098),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_4101),
.Y(n_4104)
);

INVx2_ASAP7_75t_L g4105 ( 
.A(n_4102),
.Y(n_4105)
);

OAI22xp5_ASAP7_75t_SL g4106 ( 
.A1(n_4105),
.A2(n_4094),
.B1(n_4104),
.B2(n_4103),
.Y(n_4106)
);

BUFx2_ASAP7_75t_L g4107 ( 
.A(n_4106),
.Y(n_4107)
);

OAI21xp5_ASAP7_75t_L g4108 ( 
.A1(n_4107),
.A2(n_4092),
.B(n_4095),
.Y(n_4108)
);

AO22x2_ASAP7_75t_L g4109 ( 
.A1(n_4108),
.A2(n_4091),
.B1(n_4093),
.B2(n_4084),
.Y(n_4109)
);

AOI22xp5_ASAP7_75t_L g4110 ( 
.A1(n_4109),
.A2(n_4065),
.B1(n_2541),
.B2(n_2754),
.Y(n_4110)
);


endmodule