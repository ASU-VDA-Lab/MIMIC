module fake_jpeg_372_n_297 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_297);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_41),
.Y(n_43)
);

INVx5_ASAP7_75t_SL g74 ( 
.A(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_47),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_45),
.B(n_54),
.Y(n_99)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_50),
.Y(n_104)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_25),
.B(n_27),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_29),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_31),
.B1(n_39),
.B2(n_30),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_2),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_4),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_70),
.A2(n_71),
.B1(n_85),
.B2(n_88),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_44),
.B1(n_64),
.B2(n_45),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_63),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_37),
.B1(n_19),
.B2(n_22),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_73),
.A2(n_93),
.B1(n_96),
.B2(n_103),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_30),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_78),
.B(n_79),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_33),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_80),
.B(n_109),
.Y(n_114)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_39),
.B1(n_31),
.B2(n_22),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_19),
.B1(n_22),
.B2(n_32),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_101),
.Y(n_121)
);

INVx5_ASAP7_75t_SL g91 ( 
.A(n_62),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_92),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_54),
.A2(n_32),
.B1(n_26),
.B2(n_25),
.Y(n_93)
);

BUFx2_ASAP7_75t_SL g94 ( 
.A(n_56),
.Y(n_94)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_57),
.A2(n_37),
.B1(n_22),
.B2(n_19),
.Y(n_96)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_46),
.B(n_26),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_49),
.A2(n_37),
.B1(n_42),
.B2(n_36),
.Y(n_103)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_6),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_6),
.B(n_7),
.Y(n_110)
);

NOR4xp25_ASAP7_75t_SL g173 ( 
.A(n_110),
.B(n_14),
.C(n_15),
.D(n_16),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_41),
.B(n_42),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_112),
.B(n_118),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_103),
.A2(n_67),
.B1(n_63),
.B2(n_36),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g164 ( 
.A1(n_115),
.A2(n_123),
.B1(n_23),
.B2(n_21),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_67),
.B1(n_63),
.B2(n_62),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_73),
.B1(n_87),
.B2(n_82),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_77),
.B(n_67),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_106),
.C(n_98),
.Y(n_152)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_122),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_92),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_8),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_8),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_10),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_10),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_134),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_75),
.B(n_10),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_135),
.Y(n_153)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_11),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_11),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_12),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_91),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_12),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_161),
.B1(n_162),
.B2(n_169),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_82),
.B1(n_76),
.B2(n_102),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_160),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_111),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_98),
.C(n_106),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_168),
.C(n_141),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_121),
.B(n_83),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_155),
.B(n_167),
.Y(n_191)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_159),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_136),
.A2(n_76),
.B1(n_87),
.B2(n_107),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_110),
.A2(n_100),
.B1(n_81),
.B2(n_89),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_115),
.A2(n_81),
.B1(n_107),
.B2(n_41),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_164),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_166),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_114),
.B(n_137),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_118),
.B(n_41),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_123),
.B1(n_131),
.B2(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_129),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_14),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_172),
.B(n_15),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_138),
.C(n_125),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_135),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_177),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_163),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_199),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_183),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_139),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_139),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_197),
.C(n_168),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_160),
.A2(n_125),
.B1(n_124),
.B2(n_119),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_161),
.B1(n_162),
.B2(n_145),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_111),
.B(n_113),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_185),
.A2(n_188),
.B(n_148),
.Y(n_215)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_133),
.C(n_113),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_167),
.B(n_16),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_165),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_156),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_151),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_170),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_176),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_198),
.B(n_158),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_204),
.B(n_207),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_211),
.C(n_223),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_191),
.B(n_156),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_168),
.C(n_171),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_183),
.B(n_165),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_213),
.Y(n_227)
);

OAI32xp33_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_157),
.A3(n_166),
.B1(n_172),
.B2(n_169),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_190),
.B(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_153),
.C(n_157),
.Y(n_223)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_153),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_199),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_215),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_218),
.A2(n_190),
.B1(n_203),
.B2(n_186),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_230),
.B1(n_231),
.B2(n_238),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_186),
.B1(n_179),
.B2(n_182),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_219),
.A2(n_182),
.B1(n_184),
.B2(n_202),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_204),
.B(n_178),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_237),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_205),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_224),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_219),
.A2(n_157),
.B1(n_200),
.B2(n_187),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_210),
.A2(n_200),
.B1(n_192),
.B2(n_201),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_241),
.B1(n_231),
.B2(n_228),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_213),
.A2(n_173),
.B1(n_151),
.B2(n_175),
.Y(n_241)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_146),
.C(n_176),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_229),
.C(n_222),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_244),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_234),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_212),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_257),
.B1(n_233),
.B2(n_237),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_206),
.C(n_223),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_255),
.C(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_232),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_227),
.B(n_211),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_235),
.B(n_207),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_256),
.B(n_221),
.Y(n_267)
);

AOI22x1_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_208),
.B1(n_214),
.B2(n_216),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_247),
.A2(n_233),
.B1(n_230),
.B2(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_245),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_263),
.Y(n_275)
);

OAI321xp33_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_235),
.A3(n_217),
.B1(n_221),
.B2(n_226),
.C(n_205),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_250),
.B(n_146),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_267),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_238),
.B(n_240),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_251),
.B(n_247),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_273),
.Y(n_283)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_252),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_255),
.C(n_249),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_276),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_246),
.C(n_214),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_272),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_280),
.Y(n_287)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

OAI221xp5_ASAP7_75t_L g281 ( 
.A1(n_275),
.A2(n_264),
.B1(n_261),
.B2(n_266),
.C(n_258),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_281),
.B(n_239),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_270),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_273),
.C(n_276),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_286),
.B(n_288),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_274),
.B(n_277),
.Y(n_288)
);

NOR2x1_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_278),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_291),
.B(n_193),
.Y(n_293)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_287),
.A3(n_248),
.B1(n_216),
.B2(n_242),
.C1(n_151),
.C2(n_209),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_293),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_289),
.B(n_242),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_175),
.C(n_159),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_159),
.Y(n_297)
);


endmodule