module fake_ariane_1876_n_880 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_880);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_880;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_818;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_821;
wire n_218;
wire n_839;
wire n_770;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_277;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_658;
wire n_616;
wire n_630;
wire n_705;
wire n_570;
wire n_362;
wire n_260;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_664;
wire n_629;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_66),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_161),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_130),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_46),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_86),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_51),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_61),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_175),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_156),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_65),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_60),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_143),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_127),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_34),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_94),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_183),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_2),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_124),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_109),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_6),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_149),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_113),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_97),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_37),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_74),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_56),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_6),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_163),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_3),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_103),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_99),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_92),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_137),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_87),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_5),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_10),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_54),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_69),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_95),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_146),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_167),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_20),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_125),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_16),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_142),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_4),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_191),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_24),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_136),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_100),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_122),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_176),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_152),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_123),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_155),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_26),
.Y(n_254)
);

INVx4_ASAP7_75t_R g255 ( 
.A(n_116),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_73),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_154),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_187),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_133),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_108),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_169),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_131),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_159),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_153),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_39),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_83),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_222),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_211),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_216),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_211),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_216),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_216),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_211),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_196),
.B(n_198),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_212),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_0),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_223),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_212),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_232),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_221),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_221),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_238),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_203),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_225),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_204),
.B(n_0),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_245),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_254),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_206),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_208),
.B(n_1),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_229),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_231),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_200),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_236),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_240),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_194),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_195),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_251),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_197),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_199),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_202),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_253),
.B(n_258),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_207),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_209),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_205),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_205),
.B(n_1),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_210),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_250),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_213),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_264),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_264),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_214),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_217),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_201),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_237),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_267),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_271),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_257),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_268),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_270),
.B(n_218),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_275),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_307),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_289),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_219),
.Y(n_330)
);

OAI21x1_ASAP7_75t_L g331 ( 
.A1(n_288),
.A2(n_255),
.B(n_193),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_301),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_193),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_291),
.B(n_193),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_220),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_303),
.B(n_224),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_310),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_270),
.A2(n_266),
.B1(n_265),
.B2(n_263),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_312),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_313),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_193),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_314),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_293),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_300),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_308),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_292),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_278),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_305),
.B(n_226),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_277),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_280),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_311),
.B(n_227),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_279),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_272),
.B(n_228),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_273),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_282),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_283),
.Y(n_359)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_287),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_306),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_309),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_309),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_316),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_316),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_281),
.Y(n_367)
);

AND2x6_ASAP7_75t_L g368 ( 
.A(n_272),
.B(n_27),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_284),
.Y(n_369)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_368),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_362),
.B(n_274),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g372 ( 
.A(n_346),
.B(n_290),
.C(n_274),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_337),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_348),
.B(n_230),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_301),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_233),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_344),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

INVx6_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_362),
.B(n_302),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_337),
.Y(n_382)
);

AND2x2_ASAP7_75t_SL g383 ( 
.A(n_362),
.B(n_302),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_323),
.B(n_315),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_324),
.B(n_315),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_234),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_349),
.A2(n_249),
.B1(n_262),
.B2(n_261),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_361),
.A2(n_247),
.B1(n_260),
.B2(n_259),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_345),
.Y(n_389)
);

NAND2xp33_ASAP7_75t_L g390 ( 
.A(n_362),
.B(n_235),
.Y(n_390)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_362),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_368),
.B(n_363),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_341),
.B(n_286),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_341),
.B(n_2),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_337),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_343),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_328),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_360),
.Y(n_399)
);

INVx4_ASAP7_75t_SL g400 ( 
.A(n_368),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_332),
.B(n_3),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_363),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_328),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_327),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_349),
.A2(n_256),
.B1(n_252),
.B2(n_248),
.Y(n_405)
);

OAI22xp33_ASAP7_75t_L g406 ( 
.A1(n_350),
.A2(n_347),
.B1(n_361),
.B2(n_363),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_327),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_353),
.B(n_239),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_327),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_319),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_339),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_363),
.Y(n_413)
);

NOR2x1p5_ASAP7_75t_L g414 ( 
.A(n_366),
.B(n_242),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_340),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_340),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_321),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_321),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_353),
.B(n_244),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_320),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_342),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_322),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_368),
.A2(n_246),
.B1(n_5),
.B2(n_7),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_333),
.B(n_28),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_364),
.Y(n_426)
);

BUFx4f_ASAP7_75t_L g427 ( 
.A(n_364),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_322),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_333),
.B(n_29),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_320),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_325),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_334),
.B(n_341),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_352),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_364),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_364),
.B(n_4),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_364),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_353),
.B(n_30),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_368),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_360),
.Y(n_440)
);

OAI221xp5_ASAP7_75t_L g441 ( 
.A1(n_387),
.A2(n_350),
.B1(n_318),
.B2(n_352),
.C(n_359),
.Y(n_441)
);

AO22x2_ASAP7_75t_L g442 ( 
.A1(n_394),
.A2(n_325),
.B1(n_358),
.B2(n_359),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_386),
.B(n_382),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_406),
.A2(n_365),
.B1(n_366),
.B2(n_367),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_434),
.Y(n_445)
);

AO22x2_ASAP7_75t_L g446 ( 
.A1(n_394),
.A2(n_358),
.B1(n_357),
.B2(n_365),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_395),
.B(n_414),
.Y(n_447)
);

INVx8_ASAP7_75t_L g448 ( 
.A(n_395),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_386),
.B(n_366),
.Y(n_449)
);

AO22x2_ASAP7_75t_L g450 ( 
.A1(n_381),
.A2(n_369),
.B1(n_367),
.B2(n_319),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_398),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_402),
.B(n_369),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_376),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_373),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_406),
.B(n_360),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_376),
.A2(n_329),
.B1(n_355),
.B2(n_368),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_385),
.B(n_360),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_393),
.A2(n_368),
.B1(n_356),
.B2(n_326),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_382),
.B(n_330),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_432),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_375),
.B(n_335),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_L g462 ( 
.A(n_372),
.B(n_338),
.Y(n_462)
);

AO22x2_ASAP7_75t_L g463 ( 
.A1(n_381),
.A2(n_329),
.B1(n_351),
.B2(n_336),
.Y(n_463)
);

BUFx8_ASAP7_75t_L g464 ( 
.A(n_384),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_383),
.B(n_354),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_413),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_398),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_378),
.Y(n_468)
);

OAI221xp5_ASAP7_75t_L g469 ( 
.A1(n_387),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_469)
);

OAI221xp5_ASAP7_75t_L g470 ( 
.A1(n_405),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.C(n_12),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_425),
.B(n_437),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_411),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_371),
.B(n_331),
.Y(n_473)
);

OAI221xp5_ASAP7_75t_L g474 ( 
.A1(n_405),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_411),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

A2O1A1Ixp33_ASAP7_75t_L g477 ( 
.A1(n_423),
.A2(n_331),
.B(n_14),
.C(n_15),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

NAND2xp33_ASAP7_75t_L g479 ( 
.A(n_439),
.B(n_13),
.Y(n_479)
);

AO22x2_ASAP7_75t_L g480 ( 
.A1(n_401),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_375),
.B(n_377),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_398),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_407),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_439),
.B(n_31),
.Y(n_484)
);

OR2x2_ASAP7_75t_SL g485 ( 
.A(n_383),
.B(n_17),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_403),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_377),
.B(n_18),
.Y(n_487)
);

OR2x6_ASAP7_75t_L g488 ( 
.A(n_433),
.B(n_18),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_409),
.B(n_19),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_391),
.B(n_19),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_409),
.B(n_20),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_419),
.Y(n_492)
);

OAI221xp5_ASAP7_75t_L g493 ( 
.A1(n_423),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.C(n_24),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_388),
.Y(n_494)
);

NAND2x1p5_ASAP7_75t_L g495 ( 
.A(n_391),
.B(n_21),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_419),
.B(n_22),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_430),
.B(n_23),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_374),
.B(n_25),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_400),
.B(n_25),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_412),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_400),
.B(n_26),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_415),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_400),
.B(n_32),
.Y(n_503)
);

NAND3xp33_ASAP7_75t_SL g504 ( 
.A(n_393),
.B(n_436),
.C(n_435),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_403),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_420),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_427),
.B(n_33),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_416),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_421),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_374),
.B(n_35),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_396),
.Y(n_511)
);

OAI221xp5_ASAP7_75t_L g512 ( 
.A1(n_433),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.C(n_41),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_SL g513 ( 
.A(n_481),
.B(n_426),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_453),
.B(n_427),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_444),
.B(n_439),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_492),
.B(n_426),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_452),
.B(n_435),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_461),
.B(n_443),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_472),
.B(n_396),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_452),
.B(n_370),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_499),
.B(n_501),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_SL g522 ( 
.A(n_449),
.B(n_399),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_499),
.B(n_370),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_501),
.B(n_370),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_SL g525 ( 
.A(n_487),
.B(n_440),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_465),
.B(n_370),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_462),
.B(n_456),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_447),
.B(n_408),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_SL g529 ( 
.A(n_459),
.B(n_447),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_SL g530 ( 
.A(n_494),
.B(n_438),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_471),
.B(n_408),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_471),
.B(n_408),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_448),
.B(n_424),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_SL g534 ( 
.A(n_489),
.B(n_438),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_448),
.B(n_424),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_466),
.B(n_429),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_SL g537 ( 
.A(n_491),
.B(n_429),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_457),
.B(n_392),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_458),
.B(n_397),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_475),
.B(n_417),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_503),
.B(n_418),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_454),
.B(n_422),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_503),
.B(n_428),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_496),
.B(n_404),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_468),
.B(n_476),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_478),
.B(n_410),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_483),
.B(n_420),
.Y(n_547)
);

AND2x2_ASAP7_75t_SL g548 ( 
.A(n_479),
.B(n_390),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_500),
.B(n_420),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_502),
.B(n_380),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_508),
.B(n_431),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_509),
.B(n_380),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_497),
.B(n_42),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_SL g554 ( 
.A(n_498),
.B(n_43),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_455),
.B(n_44),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_511),
.B(n_45),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_486),
.B(n_47),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_505),
.B(n_48),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_473),
.B(n_49),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_SL g560 ( 
.A(n_510),
.B(n_50),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_451),
.B(n_52),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_467),
.B(n_53),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_446),
.B(n_55),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_482),
.B(n_57),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_441),
.B(n_58),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_445),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_506),
.B(n_59),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_490),
.B(n_62),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_SL g569 ( 
.A(n_507),
.B(n_63),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_495),
.B(n_64),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_464),
.B(n_67),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_464),
.B(n_68),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_519),
.B(n_446),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_518),
.B(n_460),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_566),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_565),
.A2(n_477),
.B(n_493),
.Y(n_576)
);

AOI221xp5_ASAP7_75t_SL g577 ( 
.A1(n_545),
.A2(n_474),
.B1(n_469),
.B2(n_470),
.C(n_542),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_552),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_559),
.A2(n_504),
.B(n_512),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_521),
.B(n_450),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_539),
.A2(n_484),
.B(n_463),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_552),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_551),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_546),
.Y(n_584)
);

OAI21x1_ASAP7_75t_L g585 ( 
.A1(n_544),
.A2(n_484),
.B(n_463),
.Y(n_585)
);

CKINVDCx16_ASAP7_75t_R g586 ( 
.A(n_530),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_537),
.A2(n_488),
.B(n_450),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_552),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_529),
.B(n_485),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_547),
.A2(n_488),
.B(n_484),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_540),
.B(n_442),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_515),
.A2(n_480),
.B(n_442),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_527),
.B(n_70),
.Y(n_593)
);

AND2x4_ASAP7_75t_SL g594 ( 
.A(n_563),
.B(n_480),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_528),
.B(n_71),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_534),
.A2(n_72),
.B(n_75),
.Y(n_596)
);

OA21x2_ASAP7_75t_L g597 ( 
.A1(n_536),
.A2(n_76),
.B(n_77),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_541),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_531),
.Y(n_599)
);

A2O1A1Ixp33_ASAP7_75t_L g600 ( 
.A1(n_525),
.A2(n_553),
.B(n_569),
.C(n_535),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_513),
.A2(n_81),
.B(n_82),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_548),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_532),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_543),
.B(n_571),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_514),
.B(n_84),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_533),
.A2(n_85),
.B(n_88),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_548),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_555),
.A2(n_93),
.B(n_96),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_517),
.B(n_98),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_L g610 ( 
.A1(n_556),
.A2(n_101),
.B(n_102),
.Y(n_610)
);

NOR2xp67_ASAP7_75t_L g611 ( 
.A(n_572),
.B(n_104),
.Y(n_611)
);

NAND2x1_ASAP7_75t_L g612 ( 
.A(n_550),
.B(n_105),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_538),
.B(n_520),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_549),
.A2(n_106),
.B(n_107),
.Y(n_614)
);

AO31x2_ASAP7_75t_L g615 ( 
.A1(n_560),
.A2(n_110),
.A3(n_111),
.B(n_112),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_516),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_523),
.B(n_118),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_522),
.Y(n_618)
);

NAND3xp33_ASAP7_75t_L g619 ( 
.A(n_554),
.B(n_119),
.C(n_120),
.Y(n_619)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_524),
.Y(n_620)
);

OAI22x1_ASAP7_75t_L g621 ( 
.A1(n_526),
.A2(n_121),
.B1(n_126),
.B2(n_128),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_574),
.B(n_570),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_575),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_573),
.B(n_568),
.Y(n_624)
);

AO21x2_ASAP7_75t_L g625 ( 
.A1(n_581),
.A2(n_558),
.B(n_557),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_582),
.B(n_567),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_578),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_582),
.Y(n_628)
);

AOI21x1_ASAP7_75t_L g629 ( 
.A1(n_587),
.A2(n_564),
.B(n_562),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_585),
.A2(n_561),
.B(n_132),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_586),
.B(n_192),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_594),
.A2(n_129),
.B1(n_134),
.B2(n_135),
.Y(n_632)
);

AOI221x1_ASAP7_75t_L g633 ( 
.A1(n_592),
.A2(n_138),
.B1(n_139),
.B2(n_141),
.C(n_144),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_593),
.Y(n_634)
);

O2A1O1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_589),
.A2(n_145),
.B(n_147),
.C(n_148),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_578),
.A2(n_150),
.B1(n_151),
.B2(n_158),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_583),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_596),
.A2(n_160),
.B(n_164),
.Y(n_638)
);

AOI21xp33_ASAP7_75t_L g639 ( 
.A1(n_576),
.A2(n_165),
.B(n_166),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_602),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_584),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_601),
.A2(n_172),
.B(n_173),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_582),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_588),
.B(n_174),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_608),
.A2(n_177),
.B(n_178),
.Y(n_645)
);

OA21x2_ASAP7_75t_L g646 ( 
.A1(n_579),
.A2(n_179),
.B(n_182),
.Y(n_646)
);

INVxp67_ASAP7_75t_SL g647 ( 
.A(n_602),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_588),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_576),
.A2(n_184),
.B(n_185),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_603),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_603),
.Y(n_651)
);

O2A1O1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_600),
.A2(n_186),
.B(n_189),
.C(n_190),
.Y(n_652)
);

NAND3xp33_ASAP7_75t_L g653 ( 
.A(n_577),
.B(n_590),
.C(n_579),
.Y(n_653)
);

NAND2x1_ASAP7_75t_L g654 ( 
.A(n_618),
.B(n_605),
.Y(n_654)
);

OA21x2_ASAP7_75t_L g655 ( 
.A1(n_614),
.A2(n_619),
.B(n_610),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_603),
.Y(n_656)
);

OAI22x1_ASAP7_75t_L g657 ( 
.A1(n_591),
.A2(n_580),
.B1(n_604),
.B2(n_599),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_599),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_620),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_613),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_595),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_611),
.A2(n_607),
.B1(n_620),
.B2(n_621),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_620),
.B(n_617),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_577),
.B(n_609),
.Y(n_664)
);

CKINVDCx8_ASAP7_75t_R g665 ( 
.A(n_597),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_658),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_660),
.B(n_614),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_641),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_647),
.B(n_615),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_641),
.Y(n_670)
);

AND2x6_ASAP7_75t_L g671 ( 
.A(n_663),
.B(n_597),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_627),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_648),
.Y(n_673)
);

INVxp67_ASAP7_75t_SL g674 ( 
.A(n_647),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_623),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_623),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_653),
.B(n_615),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_651),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_630),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_657),
.B(n_615),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_637),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_643),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_661),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_664),
.B(n_622),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_634),
.A2(n_610),
.B1(n_619),
.B2(n_616),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_646),
.Y(n_686)
);

OR2x6_ASAP7_75t_L g687 ( 
.A(n_654),
.B(n_612),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_665),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_650),
.B(n_606),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_646),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_630),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_638),
.A2(n_629),
.B(n_642),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_655),
.A2(n_598),
.B(n_649),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_646),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_625),
.Y(n_695)
);

CKINVDCx6p67_ASAP7_75t_R g696 ( 
.A(n_634),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_625),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_624),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_634),
.B(n_656),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_655),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_655),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_650),
.B(n_659),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_645),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_628),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_645),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_643),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_663),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_663),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_644),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_633),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_652),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_638),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_626),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_643),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_642),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_684),
.B(n_628),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_684),
.B(n_632),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_R g718 ( 
.A(n_699),
.B(n_631),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_678),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_R g720 ( 
.A(n_699),
.B(n_626),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_R g721 ( 
.A(n_702),
.B(n_626),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_713),
.B(n_708),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_681),
.B(n_643),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_681),
.Y(n_724)
);

BUFx10_ASAP7_75t_L g725 ( 
.A(n_672),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_R g726 ( 
.A(n_696),
.B(n_632),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_666),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_689),
.B(n_662),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_696),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_698),
.B(n_662),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_673),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_R g732 ( 
.A(n_678),
.B(n_635),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_698),
.B(n_640),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_R g734 ( 
.A(n_688),
.B(n_713),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_708),
.B(n_636),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_682),
.B(n_639),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_R g737 ( 
.A(n_688),
.B(n_669),
.Y(n_737)
);

XNOR2xp5_ASAP7_75t_L g738 ( 
.A(n_704),
.B(n_707),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_674),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_683),
.B(n_675),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_SL g741 ( 
.A(n_685),
.B(n_711),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_R g742 ( 
.A(n_669),
.B(n_677),
.Y(n_742)
);

NAND2xp33_ASAP7_75t_R g743 ( 
.A(n_669),
.B(n_677),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_683),
.B(n_675),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_R g745 ( 
.A(n_669),
.B(n_707),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_SL g746 ( 
.A(n_711),
.B(n_667),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_682),
.B(n_706),
.Y(n_747)
);

XNOR2xp5_ASAP7_75t_L g748 ( 
.A(n_706),
.B(n_682),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_R g749 ( 
.A(n_714),
.B(n_709),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_668),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_714),
.Y(n_751)
);

CKINVDCx11_ASAP7_75t_R g752 ( 
.A(n_687),
.Y(n_752)
);

NAND2xp33_ASAP7_75t_R g753 ( 
.A(n_709),
.B(n_680),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_676),
.B(n_668),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_670),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_R g756 ( 
.A(n_680),
.B(n_697),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_670),
.Y(n_757)
);

BUFx10_ASAP7_75t_L g758 ( 
.A(n_687),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_724),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_750),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_727),
.B(n_676),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_740),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_739),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_744),
.B(n_701),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_722),
.B(n_700),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_R g766 ( 
.A(n_721),
.B(n_700),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_722),
.B(n_700),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_716),
.B(n_700),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_755),
.Y(n_769)
);

INVx5_ASAP7_75t_L g770 ( 
.A(n_758),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_757),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_731),
.B(n_701),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_754),
.B(n_697),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_723),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_717),
.B(n_679),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_719),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_726),
.B(n_710),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_738),
.B(n_728),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_751),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_735),
.B(n_679),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_730),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_725),
.B(n_694),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_729),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_758),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_725),
.B(n_694),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_752),
.B(n_691),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_733),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_747),
.B(n_710),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_735),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_777),
.A2(n_693),
.B1(n_741),
.B2(n_736),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_787),
.B(n_746),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_763),
.B(n_695),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_763),
.B(n_748),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_778),
.A2(n_736),
.B1(n_687),
.B2(n_691),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_759),
.Y(n_795)
);

OAI211xp5_ASAP7_75t_L g796 ( 
.A1(n_788),
.A2(n_732),
.B(n_712),
.C(n_715),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_780),
.A2(n_687),
.B(n_686),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_780),
.B(n_695),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_759),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_775),
.B(n_712),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_775),
.B(n_715),
.Y(n_801)
);

AOI221xp5_ASAP7_75t_L g802 ( 
.A1(n_778),
.A2(n_686),
.B1(n_690),
.B2(n_715),
.C(n_705),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_771),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_771),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_760),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_760),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_767),
.B(n_715),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_769),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_767),
.B(n_705),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_768),
.B(n_703),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_769),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_805),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_792),
.B(n_774),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_798),
.B(n_786),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_790),
.A2(n_718),
.B1(n_753),
.B2(n_743),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_805),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_793),
.B(n_776),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_791),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_800),
.B(n_776),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_792),
.B(n_774),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_803),
.B(n_772),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_808),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_813),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_818),
.B(n_804),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_820),
.B(n_800),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_821),
.B(n_811),
.Y(n_826)
);

AO221x2_ASAP7_75t_L g827 ( 
.A1(n_821),
.A2(n_794),
.B1(n_799),
.B2(n_806),
.C(n_795),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_823),
.B(n_814),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_827),
.B(n_814),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_824),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_825),
.B(n_819),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_826),
.B(n_822),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_825),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_SL g834 ( 
.A(n_829),
.B(n_815),
.C(n_796),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_830),
.A2(n_817),
.B1(n_801),
.B2(n_802),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_830),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_836),
.B(n_831),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_835),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_837),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_838),
.Y(n_840)
);

BUFx8_ASAP7_75t_SL g841 ( 
.A(n_837),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_839),
.B(n_833),
.Y(n_842)
);

NOR3xp33_ASAP7_75t_L g843 ( 
.A(n_840),
.B(n_834),
.C(n_832),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_L g844 ( 
.A(n_839),
.B(n_828),
.C(n_783),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_841),
.B(n_822),
.Y(n_845)
);

AOI322xp5_ASAP7_75t_L g846 ( 
.A1(n_840),
.A2(n_781),
.A3(n_786),
.B1(n_780),
.B2(n_816),
.C1(n_812),
.C2(n_801),
.Y(n_846)
);

OAI31xp33_ASAP7_75t_L g847 ( 
.A1(n_840),
.A2(n_690),
.A3(n_782),
.B(n_785),
.Y(n_847)
);

AOI222xp33_ASAP7_75t_L g848 ( 
.A1(n_842),
.A2(n_671),
.B1(n_782),
.B2(n_785),
.C1(n_761),
.C2(n_762),
.Y(n_848)
);

OAI221xp5_ASAP7_75t_L g849 ( 
.A1(n_843),
.A2(n_783),
.B1(n_749),
.B2(n_756),
.C(n_734),
.Y(n_849)
);

OAI211xp5_ASAP7_75t_SL g850 ( 
.A1(n_845),
.A2(n_797),
.B(n_808),
.C(n_784),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_844),
.Y(n_851)
);

AOI221xp5_ASAP7_75t_L g852 ( 
.A1(n_847),
.A2(n_772),
.B1(n_766),
.B2(n_810),
.C(n_780),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_846),
.A2(n_671),
.B1(n_742),
.B2(n_779),
.Y(n_853)
);

NOR2x1_ASAP7_75t_L g854 ( 
.A(n_851),
.B(n_687),
.Y(n_854)
);

OAI22x1_ASAP7_75t_L g855 ( 
.A1(n_853),
.A2(n_784),
.B1(n_770),
.B2(n_779),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_849),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_850),
.Y(n_857)
);

NOR2x1p5_ASAP7_75t_L g858 ( 
.A(n_848),
.B(n_807),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_857),
.B(n_852),
.Y(n_859)
);

NAND2xp33_ASAP7_75t_SL g860 ( 
.A(n_858),
.B(n_807),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_R g861 ( 
.A(n_856),
.B(n_720),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_854),
.B(n_810),
.Y(n_862)
);

NAND3xp33_ASAP7_75t_L g863 ( 
.A(n_855),
.B(n_764),
.C(n_768),
.Y(n_863)
);

XNOR2xp5_ASAP7_75t_L g864 ( 
.A(n_856),
.B(n_798),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_R g865 ( 
.A(n_856),
.B(n_737),
.Y(n_865)
);

AOI221x1_ASAP7_75t_L g866 ( 
.A1(n_860),
.A2(n_862),
.B1(n_863),
.B2(n_859),
.C(n_864),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_861),
.A2(n_865),
.B1(n_671),
.B2(n_809),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_864),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_864),
.B(n_809),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_859),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_870),
.A2(n_764),
.B1(n_703),
.B2(n_770),
.Y(n_871)
);

OAI22x1_ASAP7_75t_L g872 ( 
.A1(n_868),
.A2(n_770),
.B1(n_798),
.B2(n_765),
.Y(n_872)
);

OR5x1_ASAP7_75t_L g873 ( 
.A(n_866),
.B(n_765),
.C(n_745),
.D(n_770),
.E(n_671),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_873),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_874),
.A2(n_867),
.B1(n_871),
.B2(n_872),
.Y(n_875)
);

XNOR2xp5_ASAP7_75t_L g876 ( 
.A(n_875),
.B(n_869),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_876),
.B(n_692),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_877),
.Y(n_878)
);

OAI221xp5_ASAP7_75t_R g879 ( 
.A1(n_878),
.A2(n_770),
.B1(n_765),
.B2(n_692),
.C(n_671),
.Y(n_879)
);

AOI211xp5_ASAP7_75t_L g880 ( 
.A1(n_879),
.A2(n_765),
.B(n_789),
.C(n_773),
.Y(n_880)
);


endmodule