module fake_jpeg_16235_n_47 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_47);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_47;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_44;
wire n_24;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_25;
wire n_31;
wire n_37;
wire n_43;
wire n_29;
wire n_32;

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_31),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.C(n_38),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_1),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_23),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_6),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_40),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_41),
.B(n_39),
.Y(n_43)
);

NOR2x1_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_21),
.Y(n_45)
);

AOI322xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_22),
.A3(n_30),
.B1(n_26),
.B2(n_24),
.C1(n_28),
.C2(n_19),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_8),
.B1(n_20),
.B2(n_29),
.Y(n_47)
);


endmodule