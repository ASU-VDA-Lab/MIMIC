module fake_jpeg_15076_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx5_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx5p33_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_11),
.B(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_15),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_5),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_6),
.B1(n_9),
.B2(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_26),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_17),
.C(n_14),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_21),
.B(n_19),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_29),
.Y(n_31)
);

HAxp5_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_24),
.CON(n_30),
.SN(n_30)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B(n_16),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B(n_8),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_17),
.C(n_12),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.B1(n_13),
.B2(n_18),
.Y(n_36)
);

OAI21x1_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_17),
.B(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_10),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_5),
.B(n_20),
.Y(n_38)
);

XNOR2x2_ASAP7_75t_SL g39 ( 
.A(n_38),
.B(n_20),
.Y(n_39)
);


endmodule