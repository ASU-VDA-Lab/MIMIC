module fake_netlist_6_3738_n_1946 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1946);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1946;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_172),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_128),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_181),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_43),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_10),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_112),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_25),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_139),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_178),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_119),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_86),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_34),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_12),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_6),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_101),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_94),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_152),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_175),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_97),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_70),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_127),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_136),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_33),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_69),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_26),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_87),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_49),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_81),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_38),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_72),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_35),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_196),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_59),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_63),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_92),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_78),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_169),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_24),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_51),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_110),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_131),
.Y(n_249)
);

BUFx2_ASAP7_75t_SL g250 ( 
.A(n_39),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_171),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_91),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_41),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_122),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_14),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_60),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_183),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_102),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_0),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_16),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_66),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_13),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_161),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_66),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_163),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_129),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_46),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_93),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_150),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_10),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_83),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_3),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_3),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_157),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_201),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_2),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_75),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_69),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_9),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_156),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_27),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_108),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_151),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_85),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_41),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_59),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_38),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_177),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_0),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_188),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_194),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_130),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_73),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_30),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_191),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_61),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_118),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_180),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_186),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_40),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_158),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_23),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_28),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_31),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_13),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_95),
.Y(n_307)
);

BUFx8_ASAP7_75t_SL g308 ( 
.A(n_40),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_114),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_153),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_8),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_8),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_140),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_170),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_198),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_133),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_5),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_35),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_34),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_147),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_185),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_173),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_120),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_53),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_124),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_148),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_159),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_141),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_49),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_24),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_104),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_107),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_145),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_106),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_179),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_125),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_26),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_19),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_54),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_109),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_50),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_7),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_37),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_182),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_187),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_45),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_18),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_52),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_99),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_36),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_19),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_29),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_100),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_193),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_17),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_146),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_88),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_154),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_134),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_55),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_123),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_96),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_1),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_84),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_48),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_57),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_2),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_61),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_184),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_6),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_25),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_111),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_65),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_56),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_165),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_74),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_57),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_36),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_28),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_17),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_89),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_190),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_77),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_7),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_15),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_52),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_33),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_44),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_68),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_168),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_5),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_4),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_132),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_68),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_71),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_45),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_189),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_44),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_12),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_160),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_20),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_47),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_113),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_62),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_308),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_288),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_305),
.B(n_1),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_255),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_223),
.B(n_4),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_232),
.B(n_316),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_337),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_258),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_224),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_358),
.B(n_9),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_337),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_252),
.Y(n_419)
);

INVxp33_ASAP7_75t_SL g420 ( 
.A(n_280),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_337),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_337),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g423 ( 
.A(n_236),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_264),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_266),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_398),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_268),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_337),
.B(n_11),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_208),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_337),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_251),
.B(n_11),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_269),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_302),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_270),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_301),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_301),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_301),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_272),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_276),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_301),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_281),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_283),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_301),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_284),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_285),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_368),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_302),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_278),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_368),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_368),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_368),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_336),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_368),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_336),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_282),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_L g456 ( 
.A(n_305),
.B(n_14),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_289),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_314),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_292),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_207),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_282),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_344),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_353),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_349),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_369),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_213),
.B(n_15),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_293),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_295),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_295),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_383),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_353),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_298),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_299),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_224),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_373),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_373),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_208),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_300),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_307),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_234),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_315),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_234),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_213),
.B(n_16),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_334),
.B(n_18),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_320),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_321),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_L g487 ( 
.A(n_348),
.B(n_20),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_322),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_389),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_389),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_323),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_231),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_203),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_268),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_240),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_241),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_224),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_246),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_256),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_261),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_205),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_262),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_203),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_271),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_263),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_204),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_265),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_408),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_448),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_499),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_420),
.A2(n_374),
.B1(n_260),
.B2(n_238),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_406),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_500),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_414),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_435),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_424),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_419),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_435),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_425),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_415),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_436),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_432),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_436),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_434),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_439),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_437),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_L g527 ( 
.A(n_448),
.B(n_334),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_448),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_R g529 ( 
.A(n_504),
.B(n_204),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_441),
.B(n_356),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_428),
.A2(n_235),
.B(n_227),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_442),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_444),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_437),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_445),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_471),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_440),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_412),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_438),
.Y(n_539)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_415),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_457),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_440),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_443),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_459),
.B(n_356),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_467),
.Y(n_545)
);

NOR2xp67_ASAP7_75t_L g546 ( 
.A(n_448),
.B(n_211),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_443),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_423),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_480),
.B(n_348),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_411),
.B(n_309),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_458),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_473),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_446),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_446),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_449),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_449),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_478),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_479),
.B(n_227),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_450),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_474),
.B(n_206),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_410),
.A2(n_313),
.B(n_235),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_450),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_488),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_451),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_491),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_451),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_453),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_462),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_472),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_453),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_481),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_464),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_476),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_485),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_476),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_410),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_486),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_413),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_413),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_417),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_417),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_493),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_483),
.B(n_403),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_433),
.B(n_313),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_418),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_418),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_447),
.B(n_397),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_503),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_460),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_529),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_585),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_576),
.Y(n_592)
);

AND2x2_ASAP7_75t_SL g593 ( 
.A(n_550),
.B(n_409),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_583),
.A2(n_506),
.B1(n_416),
.B2(n_431),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_538),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_558),
.B(n_501),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_L g597 ( 
.A(n_584),
.B(n_278),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_536),
.B(n_452),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_536),
.B(n_549),
.Y(n_599)
);

INVx4_ASAP7_75t_SL g600 ( 
.A(n_585),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_536),
.B(n_454),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_589),
.B(n_463),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_585),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_576),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_549),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_530),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_SL g607 ( 
.A(n_544),
.B(n_371),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_578),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_587),
.B(n_278),
.Y(n_609)
);

NAND3x1_ASAP7_75t_L g610 ( 
.A(n_511),
.B(n_484),
.C(n_466),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_578),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_515),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_580),
.B(n_474),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_585),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_580),
.A2(n_371),
.B1(n_456),
.B2(n_407),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_586),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_586),
.B(n_579),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_579),
.B(n_471),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_515),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_555),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_585),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_585),
.Y(n_622)
);

OAI22xp33_ASAP7_75t_L g623 ( 
.A1(n_511),
.A2(n_254),
.B1(n_257),
.B2(n_217),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_512),
.B(n_427),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_560),
.A2(n_489),
.B1(n_426),
.B2(n_470),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_520),
.B(n_426),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_508),
.B(n_397),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_547),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_520),
.B(n_429),
.Y(n_629)
);

NOR2x1p5_ASAP7_75t_L g630 ( 
.A(n_514),
.B(n_497),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_581),
.B(n_471),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_540),
.B(n_429),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_555),
.Y(n_633)
);

INVx4_ASAP7_75t_SL g634 ( 
.A(n_547),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_581),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_548),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_547),
.Y(n_637)
);

AND3x1_ASAP7_75t_L g638 ( 
.A(n_510),
.B(n_297),
.C(n_279),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_518),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_518),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_540),
.B(n_497),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_509),
.B(n_421),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_561),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_582),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_521),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_L g646 ( 
.A(n_509),
.B(n_278),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_521),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_523),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_509),
.B(n_421),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_561),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_513),
.B(n_494),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_516),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_531),
.A2(n_456),
.B1(n_407),
.B2(n_487),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_547),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_509),
.B(n_528),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_547),
.Y(n_656)
);

CKINVDCx16_ASAP7_75t_R g657 ( 
.A(n_517),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_588),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_523),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_528),
.Y(n_660)
);

AND2x2_ASAP7_75t_SL g661 ( 
.A(n_573),
.B(n_278),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_526),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_559),
.Y(n_663)
);

INVx5_ASAP7_75t_L g664 ( 
.A(n_559),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_528),
.B(n_422),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_526),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_531),
.B(n_507),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_528),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_519),
.B(n_477),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_522),
.B(n_291),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_534),
.B(n_422),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_534),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_SL g673 ( 
.A(n_524),
.B(n_247),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_525),
.B(n_477),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_532),
.B(n_482),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_537),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_533),
.B(n_291),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_537),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_542),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_542),
.B(n_291),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_543),
.A2(n_487),
.B1(n_304),
.B2(n_352),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_527),
.B(n_507),
.Y(n_682)
);

INVxp33_ASAP7_75t_L g683 ( 
.A(n_573),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_543),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_553),
.A2(n_342),
.B1(n_391),
.B2(n_388),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_569),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_553),
.B(n_430),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_559),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_527),
.B(n_505),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_559),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_559),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_562),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_571),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_554),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_554),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_556),
.Y(n_696)
);

AND2x6_ASAP7_75t_L g697 ( 
.A(n_556),
.B(n_291),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_535),
.B(n_291),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_541),
.B(n_354),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_545),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_564),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_564),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_566),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_566),
.Y(n_704)
);

INVx4_ASAP7_75t_SL g705 ( 
.A(n_562),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_567),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_567),
.B(n_430),
.Y(n_707)
);

AND2x2_ASAP7_75t_SL g708 ( 
.A(n_575),
.B(n_354),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_570),
.B(n_212),
.Y(n_709)
);

AND2x6_ASAP7_75t_L g710 ( 
.A(n_570),
.B(n_354),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_552),
.B(n_557),
.Y(n_711)
);

INVx5_ASAP7_75t_L g712 ( 
.A(n_562),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_562),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_562),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_563),
.B(n_482),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_539),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_575),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_546),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_565),
.B(n_490),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_546),
.Y(n_720)
);

BUFx10_ASAP7_75t_L g721 ( 
.A(n_577),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_574),
.Y(n_722)
);

BUFx8_ASAP7_75t_SL g723 ( 
.A(n_551),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_568),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_572),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_550),
.B(n_354),
.Y(n_726)
);

AND2x2_ASAP7_75t_SL g727 ( 
.A(n_550),
.B(n_354),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_583),
.A2(n_365),
.B1(n_318),
.B2(n_339),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_550),
.B(n_490),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_550),
.B(n_492),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_538),
.B(n_250),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_583),
.B(n_215),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_550),
.A2(n_465),
.B1(n_376),
.B2(n_335),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_515),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_585),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_515),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_582),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_583),
.B(n_220),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_576),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_727),
.B(n_225),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_730),
.B(n_405),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_727),
.B(n_237),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_593),
.B(n_606),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_639),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_730),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_643),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_593),
.B(n_243),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_660),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_608),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_599),
.B(n_245),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_675),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_605),
.B(n_206),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_608),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_596),
.B(n_338),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_599),
.B(n_253),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_599),
.B(n_259),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_667),
.B(n_267),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_667),
.B(n_275),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_723),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_618),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_660),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_643),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_729),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_729),
.B(n_294),
.Y(n_764)
);

NAND2x1p5_ASAP7_75t_L g765 ( 
.A(n_667),
.B(n_296),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_602),
.B(n_268),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_631),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_592),
.B(n_310),
.Y(n_768)
);

BUFx8_ASAP7_75t_L g769 ( 
.A(n_711),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_613),
.A2(n_209),
.B1(n_214),
.B2(n_219),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_604),
.B(n_325),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_732),
.A2(n_355),
.B1(n_346),
.B2(n_328),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_611),
.B(n_326),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_668),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_674),
.B(n_277),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_616),
.B(n_739),
.Y(n_776)
);

O2A1O1Ixp5_ASAP7_75t_L g777 ( 
.A1(n_726),
.A2(n_393),
.B(n_331),
.C(n_340),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_643),
.B(n_327),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_668),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_717),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_643),
.Y(n_781)
);

AND2x4_ASAP7_75t_SL g782 ( 
.A(n_721),
.B(n_277),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_661),
.B(n_345),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_653),
.B(n_357),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_629),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_717),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_661),
.B(n_708),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_726),
.A2(n_402),
.B(n_343),
.C(n_379),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_653),
.B(n_362),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_613),
.B(n_277),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_651),
.B(n_306),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_738),
.B(n_364),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_728),
.A2(n_385),
.B1(n_392),
.B2(n_303),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_669),
.B(n_306),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_598),
.B(n_381),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_715),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_632),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_708),
.B(n_382),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_594),
.B(n_400),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_717),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_601),
.A2(n_505),
.B(n_502),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_650),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_650),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_SL g804 ( 
.A1(n_700),
.A2(n_306),
.B1(n_218),
.B2(n_216),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_669),
.B(n_209),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_SL g806 ( 
.A1(n_652),
.A2(n_218),
.B1(n_216),
.B2(n_210),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_617),
.B(n_214),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_639),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_626),
.B(n_492),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_683),
.A2(n_502),
.B(n_498),
.C(n_496),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_640),
.B(n_219),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_655),
.B(n_221),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_719),
.B(n_221),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_719),
.B(n_273),
.C(n_404),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_645),
.B(n_222),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_683),
.B(n_222),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_642),
.B(n_226),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_610),
.A2(n_226),
.B1(n_395),
.B2(n_390),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_648),
.B(n_228),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_627),
.B(n_228),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_649),
.B(n_665),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_659),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_662),
.B(n_233),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_666),
.B(n_233),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_672),
.B(n_239),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_SL g826 ( 
.A(n_652),
.B(n_590),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_728),
.A2(n_681),
.B1(n_615),
.B2(n_623),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_681),
.A2(n_210),
.B1(n_401),
.B2(n_399),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_647),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_676),
.B(n_684),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_694),
.B(n_239),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_610),
.A2(n_242),
.B1(n_244),
.B2(n_248),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_647),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_695),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_702),
.B(n_242),
.Y(n_835)
);

O2A1O1Ixp5_ASAP7_75t_L g836 ( 
.A1(n_706),
.A2(n_498),
.B(n_496),
.C(n_495),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_678),
.B(n_244),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_615),
.A2(n_360),
.B1(n_229),
.B2(n_230),
.Y(n_838)
);

OAI221xp5_ASAP7_75t_L g839 ( 
.A1(n_685),
.A2(n_495),
.B1(n_274),
.B2(n_286),
.C(n_287),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_678),
.B(n_248),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_624),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_679),
.B(n_696),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_652),
.B(n_475),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_641),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_679),
.B(n_249),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_682),
.B(n_455),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_696),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_701),
.B(n_249),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_627),
.B(n_332),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_600),
.Y(n_850)
);

NOR2xp67_ASAP7_75t_L g851 ( 
.A(n_733),
.B(n_332),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_625),
.B(n_475),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_SL g853 ( 
.A(n_630),
.B(n_636),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_701),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_703),
.B(n_333),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_SL g856 ( 
.A(n_644),
.B(n_333),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_703),
.B(n_335),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_704),
.Y(n_858)
);

NOR3xp33_ASAP7_75t_L g859 ( 
.A(n_623),
.B(n_290),
.C(n_311),
.Y(n_859)
);

OR2x6_ASAP7_75t_L g860 ( 
.A(n_725),
.B(n_455),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_612),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_595),
.B(n_469),
.Y(n_862)
);

BUFx5_ASAP7_75t_L g863 ( 
.A(n_714),
.Y(n_863)
);

INVx4_ASAP7_75t_L g864 ( 
.A(n_600),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_725),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_624),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_731),
.B(n_469),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_731),
.B(n_461),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_L g869 ( 
.A(n_670),
.B(n_359),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_635),
.A2(n_376),
.B(n_375),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_682),
.Y(n_871)
);

INVx8_ASAP7_75t_L g872 ( 
.A(n_731),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_685),
.A2(n_366),
.B1(n_229),
.B2(n_401),
.Y(n_873)
);

NAND2x1p5_ASAP7_75t_L g874 ( 
.A(n_682),
.B(n_461),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_677),
.B(n_361),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_638),
.A2(n_699),
.B1(n_698),
.B2(n_677),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_622),
.B(n_361),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_597),
.A2(n_366),
.B1(n_399),
.B2(n_396),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_698),
.B(n_372),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_671),
.A2(n_390),
.B(n_372),
.C(n_395),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_619),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_624),
.B(n_468),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_619),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_689),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_689),
.B(n_468),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_620),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_622),
.B(n_375),
.Y(n_887)
);

NOR3xp33_ASAP7_75t_L g888 ( 
.A(n_673),
.B(n_312),
.C(n_317),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_699),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_620),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_600),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_633),
.Y(n_892)
);

NOR2xp67_ASAP7_75t_SL g893 ( 
.A(n_603),
.B(n_207),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_628),
.B(n_319),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_720),
.B(n_324),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_718),
.B(n_230),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_718),
.B(n_687),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_597),
.A2(n_396),
.B1(n_394),
.B2(n_386),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_663),
.B(n_691),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_633),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_607),
.B(n_329),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_734),
.Y(n_902)
);

NAND2xp33_ASAP7_75t_SL g903 ( 
.A(n_722),
.B(n_330),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_734),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_736),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_736),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_743),
.B(n_658),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_744),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_861),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_882),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_805),
.B(n_673),
.C(n_607),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_787),
.A2(n_707),
.B(n_735),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_743),
.B(n_737),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_775),
.Y(n_914)
);

BUFx8_ASAP7_75t_L g915 ( 
.A(n_797),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_787),
.A2(n_735),
.B(n_591),
.Y(n_916)
);

NOR2xp67_ASAP7_75t_L g917 ( 
.A(n_751),
.B(n_686),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_744),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_897),
.A2(n_621),
.B(n_591),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_784),
.A2(n_621),
.B(n_591),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_749),
.B(n_724),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_745),
.B(n_721),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_789),
.A2(n_621),
.B(n_735),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_763),
.B(n_709),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_805),
.B(n_693),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_762),
.A2(n_690),
.B(n_654),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_813),
.B(n_741),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_757),
.A2(n_609),
.B(n_654),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_754),
.A2(n_609),
.B(n_692),
.C(n_691),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_762),
.A2(n_690),
.B(n_656),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_808),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_799),
.A2(n_646),
.B(n_713),
.C(n_692),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_754),
.B(n_794),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_876),
.B(n_721),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_757),
.A2(n_690),
.B(n_654),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_813),
.B(n_657),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_881),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_760),
.B(n_713),
.Y(n_938)
);

NOR3xp33_ASAP7_75t_L g939 ( 
.A(n_799),
.B(n_378),
.C(n_347),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_796),
.B(n_716),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_803),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_758),
.A2(n_656),
.B(n_688),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_781),
.A2(n_656),
.B(n_688),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_843),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_785),
.B(n_341),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_803),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_808),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_791),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_781),
.A2(n_688),
.B(n_603),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_766),
.B(n_716),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_883),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_747),
.B(n_723),
.Y(n_952)
);

NAND3xp33_ASAP7_75t_SL g953 ( 
.A(n_818),
.B(n_341),
.C(n_347),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_746),
.A2(n_603),
.B(n_614),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_747),
.A2(n_646),
.B(n_351),
.C(n_360),
.Y(n_955)
);

OR2x6_ASAP7_75t_L g956 ( 
.A(n_872),
.B(n_21),
.Y(n_956)
);

BUFx12f_ASAP7_75t_L g957 ( 
.A(n_769),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_816),
.B(n_350),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_746),
.A2(n_603),
.B(n_614),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_SL g960 ( 
.A1(n_790),
.A2(n_350),
.B1(n_351),
.B2(n_363),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_746),
.A2(n_614),
.B(n_712),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_833),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_767),
.B(n_764),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_854),
.Y(n_964)
);

BUFx12f_ASAP7_75t_L g965 ( 
.A(n_769),
.Y(n_965)
);

AO21x1_ASAP7_75t_L g966 ( 
.A1(n_740),
.A2(n_680),
.B(n_697),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_889),
.A2(n_386),
.B1(n_367),
.B2(n_370),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_821),
.A2(n_614),
.B(n_712),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_816),
.B(n_634),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_822),
.B(n_634),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_746),
.A2(n_712),
.B(n_637),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_821),
.A2(n_758),
.B(n_842),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_883),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_750),
.A2(n_712),
.B(n_637),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_742),
.A2(n_363),
.B(n_367),
.C(n_370),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_803),
.Y(n_976)
);

O2A1O1Ixp5_ASAP7_75t_L g977 ( 
.A1(n_783),
.A2(n_710),
.B(n_697),
.C(n_680),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_803),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_899),
.A2(n_637),
.B(n_664),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_854),
.Y(n_980)
);

AOI21x1_ASAP7_75t_L g981 ( 
.A1(n_795),
.A2(n_705),
.B(n_634),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_834),
.B(n_705),
.Y(n_982)
);

BUFx4f_ASAP7_75t_L g983 ( 
.A(n_872),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_792),
.B(n_705),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_776),
.B(n_680),
.Y(n_985)
);

AOI21x1_ASAP7_75t_L g986 ( 
.A1(n_847),
.A2(n_664),
.B(n_697),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_802),
.A2(n_664),
.B(n_697),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_880),
.A2(n_377),
.B(n_378),
.C(n_380),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_755),
.A2(n_710),
.B(n_697),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_829),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_827),
.A2(n_394),
.B1(n_384),
.B2(n_380),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_756),
.A2(n_710),
.B(n_680),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_753),
.B(n_79),
.Y(n_993)
);

AOI21xp33_ASAP7_75t_L g994 ( 
.A1(n_820),
.A2(n_377),
.B(n_384),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_830),
.A2(n_710),
.B(n_680),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_846),
.B(n_200),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_860),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_780),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_856),
.B(n_22),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_748),
.A2(n_195),
.B(n_174),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_875),
.B(n_22),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_748),
.A2(n_167),
.B(n_164),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_786),
.A2(n_155),
.B(n_149),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_820),
.B(n_849),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_761),
.A2(n_144),
.B(n_143),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_849),
.B(n_27),
.Y(n_1006)
);

BUFx4f_ASAP7_75t_L g1007 ( 
.A(n_872),
.Y(n_1007)
);

BUFx8_ASAP7_75t_L g1008 ( 
.A(n_865),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_860),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_800),
.A2(n_142),
.B(n_138),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_862),
.B(n_29),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_826),
.B(n_30),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_890),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_879),
.A2(n_870),
.B(n_827),
.C(n_871),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_783),
.A2(n_32),
.B(n_37),
.C(n_39),
.Y(n_1015)
);

AO22x1_ASAP7_75t_L g1016 ( 
.A1(n_859),
.A2(n_32),
.B1(n_42),
.B2(n_43),
.Y(n_1016)
);

INVx11_ASAP7_75t_L g1017 ( 
.A(n_853),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_809),
.B(n_46),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_884),
.B(n_47),
.Y(n_1019)
);

INVx6_ASAP7_75t_L g1020 ( 
.A(n_865),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_852),
.B(n_48),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_774),
.B(n_50),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_890),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_779),
.B(n_51),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_844),
.B(n_53),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_846),
.B(n_54),
.Y(n_1026)
);

INVx5_ASAP7_75t_L g1027 ( 
.A(n_850),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_761),
.A2(n_891),
.B(n_864),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_851),
.A2(n_55),
.B(n_56),
.C(n_58),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_850),
.A2(n_90),
.B(n_135),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_864),
.A2(n_82),
.B(n_126),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_867),
.B(n_58),
.Y(n_1032)
);

NOR2xp67_ASAP7_75t_L g1033 ( 
.A(n_814),
.B(n_98),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_885),
.B(n_858),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_891),
.A2(n_80),
.B(n_121),
.Y(n_1035)
);

OAI321xp33_ASAP7_75t_L g1036 ( 
.A1(n_772),
.A2(n_60),
.A3(n_62),
.B1(n_63),
.B2(n_64),
.C(n_65),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_885),
.B(n_64),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_765),
.A2(n_115),
.B1(n_76),
.B2(n_103),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_770),
.B(n_67),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_868),
.B(n_105),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_894),
.A2(n_116),
.B(n_117),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_895),
.A2(n_137),
.B1(n_812),
.B2(n_817),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_896),
.A2(n_788),
.B(n_901),
.C(n_895),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_896),
.A2(n_901),
.B(n_798),
.C(n_773),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_874),
.B(n_855),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_798),
.A2(n_771),
.B(n_768),
.C(n_869),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_765),
.A2(n_904),
.B(n_900),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_877),
.A2(n_887),
.B(n_837),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_848),
.B(n_900),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_904),
.B(n_906),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_860),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_SL g1052 ( 
.A1(n_810),
.A2(n_857),
.B(n_845),
.C(n_840),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_811),
.B(n_824),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_817),
.A2(n_905),
.B(n_902),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_886),
.A2(n_892),
.B(n_807),
.Y(n_1055)
);

OAI21xp33_ASAP7_75t_L g1056 ( 
.A1(n_838),
.A2(n_793),
.B(n_828),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_782),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_807),
.A2(n_840),
.B(n_857),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_845),
.A2(n_835),
.B(n_823),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_815),
.B(n_831),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_819),
.B(n_825),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_801),
.A2(n_752),
.B(n_777),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_863),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_841),
.A2(n_866),
.B1(n_793),
.B2(n_804),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_836),
.A2(n_903),
.B(n_832),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_893),
.B(n_863),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_839),
.A2(n_888),
.B(n_863),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_863),
.A2(n_898),
.B(n_878),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_878),
.A2(n_898),
.B1(n_806),
.B2(n_838),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_828),
.A2(n_873),
.B(n_863),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_863),
.B(n_782),
.Y(n_1071)
);

OAI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_759),
.A2(n_745),
.B1(n_763),
.B2(n_594),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_873),
.A2(n_787),
.B(n_778),
.Y(n_1073)
);

NAND2x1p5_ASAP7_75t_L g1074 ( 
.A(n_762),
.B(n_781),
.Y(n_1074)
);

AO22x1_ASAP7_75t_L g1075 ( 
.A1(n_805),
.A2(n_813),
.B1(n_859),
.B2(n_849),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_745),
.A2(n_727),
.B1(n_763),
.B2(n_593),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_745),
.A2(n_727),
.B1(n_763),
.B2(n_593),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_778),
.A2(n_897),
.B(n_789),
.Y(n_1078)
);

AOI21x1_ASAP7_75t_L g1079 ( 
.A1(n_897),
.A2(n_778),
.B(n_821),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_743),
.A2(n_593),
.B1(n_727),
.B2(n_876),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_778),
.A2(n_897),
.B(n_789),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_778),
.A2(n_897),
.B(n_789),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1027),
.A2(n_1081),
.B(n_1078),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1004),
.A2(n_1068),
.B(n_1073),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_927),
.B(n_925),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_1006),
.A2(n_1056),
.B(n_958),
.C(n_1080),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1068),
.A2(n_1014),
.B(n_972),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1075),
.A2(n_933),
.B1(n_1069),
.B2(n_1076),
.Y(n_1088)
);

NOR2xp67_ASAP7_75t_L g1089 ( 
.A(n_914),
.B(n_948),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_963),
.B(n_1060),
.Y(n_1090)
);

NAND2x1p5_ASAP7_75t_L g1091 ( 
.A(n_1027),
.B(n_941),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_924),
.B(n_1077),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_1070),
.A2(n_1058),
.B(n_1043),
.C(n_1001),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1059),
.B(n_1049),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1027),
.A2(n_1081),
.B(n_1078),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_1072),
.B(n_944),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_915),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_915),
.Y(n_1098)
);

NOR2x1_ASAP7_75t_SL g1099 ( 
.A(n_1027),
.B(n_1063),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_1020),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_919),
.A2(n_968),
.B(n_972),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_909),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_919),
.A2(n_968),
.B(n_930),
.Y(n_1103)
);

AO22x1_ASAP7_75t_L g1104 ( 
.A1(n_1039),
.A2(n_1012),
.B1(n_999),
.B2(n_936),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_934),
.A2(n_911),
.B1(n_907),
.B2(n_913),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_926),
.A2(n_943),
.B(n_981),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_953),
.A2(n_994),
.B1(n_939),
.B2(n_1021),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1040),
.B(n_917),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1082),
.A2(n_1047),
.B(n_1048),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_921),
.B(n_1040),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1048),
.A2(n_928),
.B(n_1046),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_921),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1058),
.A2(n_1044),
.B(n_1059),
.C(n_1042),
.Y(n_1113)
);

NOR2x1_ASAP7_75t_L g1114 ( 
.A(n_1071),
.B(n_922),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_910),
.B(n_950),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1053),
.B(n_1061),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1045),
.B(n_998),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1067),
.A2(n_1065),
.B(n_912),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_935),
.A2(n_942),
.B(n_923),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_1008),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_SL g1121 ( 
.A1(n_1003),
.A2(n_1010),
.B(n_1015),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_908),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1018),
.B(n_1011),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_920),
.A2(n_923),
.B(n_916),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1067),
.A2(n_975),
.B(n_1055),
.C(n_988),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_920),
.A2(n_1054),
.B(n_1055),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1032),
.B(n_960),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1054),
.A2(n_949),
.B(n_979),
.Y(n_1128)
);

INVxp67_ASAP7_75t_SL g1129 ( 
.A(n_1074),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_938),
.B(n_918),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_945),
.B(n_997),
.Y(n_1131)
);

NAND2x1_ASAP7_75t_L g1132 ( 
.A(n_941),
.B(n_946),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_929),
.A2(n_966),
.A3(n_1062),
.B(n_1019),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_1020),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_977),
.A2(n_1062),
.B(n_1050),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_996),
.B(n_1034),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_931),
.A2(n_980),
.B(n_947),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_940),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_974),
.A2(n_971),
.B(n_954),
.Y(n_1139)
);

O2A1O1Ixp5_ASAP7_75t_L g1140 ( 
.A1(n_984),
.A2(n_1022),
.B(n_1024),
.C(n_985),
.Y(n_1140)
);

BUFx2_ASAP7_75t_SL g1141 ( 
.A(n_996),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_SL g1142 ( 
.A1(n_1074),
.A2(n_1066),
.B(n_932),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1020),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1028),
.A2(n_1066),
.B(n_970),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_982),
.A2(n_1052),
.B(n_946),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_1029),
.A2(n_992),
.A3(n_989),
.B(n_995),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_959),
.A2(n_961),
.B(n_986),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_987),
.A2(n_964),
.B(n_962),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1026),
.A2(n_1037),
.B1(n_1064),
.B2(n_993),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1009),
.B(n_1051),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_937),
.A2(n_951),
.B(n_973),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_1038),
.A2(n_1041),
.A3(n_1013),
.B(n_1023),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_955),
.A2(n_990),
.B(n_1033),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1000),
.A2(n_1005),
.B(n_1002),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_976),
.A2(n_978),
.B(n_993),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_976),
.A2(n_978),
.B(n_1030),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1025),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1031),
.A2(n_1035),
.B(n_1007),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_983),
.A2(n_1007),
.B(n_1057),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_991),
.B(n_1016),
.Y(n_1160)
);

AOI21x1_ASAP7_75t_L g1161 ( 
.A1(n_967),
.A2(n_956),
.B(n_1036),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_952),
.B(n_956),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_956),
.A2(n_983),
.B1(n_1008),
.B2(n_957),
.Y(n_1163)
);

AO21x1_ASAP7_75t_L g1164 ( 
.A1(n_1017),
.A2(n_1004),
.B(n_1006),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_965),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1004),
.A2(n_927),
.B(n_1006),
.C(n_1056),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_919),
.A2(n_968),
.B(n_972),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1027),
.A2(n_781),
.B(n_762),
.Y(n_1168)
);

OAI22x1_ASAP7_75t_L g1169 ( 
.A1(n_927),
.A2(n_1004),
.B1(n_511),
.B2(n_925),
.Y(n_1169)
);

AOI21xp33_ASAP7_75t_L g1170 ( 
.A1(n_1004),
.A2(n_927),
.B(n_1006),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1027),
.A2(n_781),
.B(n_762),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1004),
.A2(n_927),
.B1(n_1075),
.B2(n_933),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1006),
.A2(n_929),
.A3(n_1014),
.B(n_1004),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_921),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1004),
.B(n_745),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_944),
.B(n_921),
.Y(n_1176)
);

OA22x2_ASAP7_75t_L g1177 ( 
.A1(n_1056),
.A2(n_1069),
.B1(n_511),
.B2(n_745),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1004),
.A2(n_1068),
.B(n_1073),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_919),
.A2(n_968),
.B(n_972),
.Y(n_1179)
);

AO21x1_ASAP7_75t_L g1180 ( 
.A1(n_1004),
.A2(n_1006),
.B(n_1001),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_919),
.A2(n_968),
.B(n_972),
.Y(n_1181)
);

AOI21x1_ASAP7_75t_L g1182 ( 
.A1(n_969),
.A2(n_1079),
.B(n_1078),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1004),
.B(n_745),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_919),
.A2(n_968),
.B(n_972),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_908),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_919),
.A2(n_968),
.B(n_972),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1004),
.B(n_745),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1027),
.A2(n_781),
.B(n_762),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1004),
.B(n_927),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1027),
.A2(n_781),
.B(n_762),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_944),
.B(n_921),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_921),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_908),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1004),
.A2(n_927),
.B(n_1006),
.C(n_1056),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1004),
.B(n_745),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1004),
.B(n_745),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_915),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_910),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1004),
.A2(n_1068),
.B(n_1073),
.Y(n_1199)
);

INVxp67_ASAP7_75t_L g1200 ( 
.A(n_910),
.Y(n_1200)
);

NOR2xp67_ASAP7_75t_L g1201 ( 
.A(n_914),
.B(n_590),
.Y(n_1201)
);

AOI21x1_ASAP7_75t_L g1202 ( 
.A1(n_969),
.A2(n_1079),
.B(n_1078),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1078),
.A2(n_1082),
.B(n_1081),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_L g1204 ( 
.A1(n_969),
.A2(n_1079),
.B(n_1078),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_919),
.A2(n_968),
.B(n_972),
.Y(n_1205)
);

BUFx8_ASAP7_75t_L g1206 ( 
.A(n_957),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1004),
.A2(n_1080),
.B1(n_1056),
.B2(n_827),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1004),
.A2(n_1068),
.B(n_1073),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_908),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1004),
.B(n_927),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1004),
.B(n_927),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_919),
.A2(n_968),
.B(n_972),
.Y(n_1212)
);

AOI21xp33_ASAP7_75t_L g1213 ( 
.A1(n_1004),
.A2(n_927),
.B(n_1006),
.Y(n_1213)
);

BUFx10_ASAP7_75t_L g1214 ( 
.A(n_952),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1027),
.A2(n_781),
.B(n_762),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1008),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_950),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_933),
.B(n_745),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1004),
.A2(n_1068),
.B(n_1073),
.Y(n_1219)
);

AND3x4_ASAP7_75t_L g1220 ( 
.A(n_917),
.B(n_859),
.C(n_888),
.Y(n_1220)
);

INVx8_ASAP7_75t_L g1221 ( 
.A(n_1027),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_944),
.B(n_921),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1078),
.A2(n_1082),
.B(n_1081),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1006),
.A2(n_929),
.A3(n_1014),
.B(n_1004),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1004),
.B(n_745),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1004),
.A2(n_927),
.B(n_1006),
.C(n_1056),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_1027),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1221),
.Y(n_1228)
);

AO22x1_ASAP7_75t_L g1229 ( 
.A1(n_1085),
.A2(n_1220),
.B1(n_1110),
.B2(n_1191),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1206),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1115),
.Y(n_1231)
);

NAND2xp33_ASAP7_75t_L g1232 ( 
.A(n_1166),
.B(n_1194),
.Y(n_1232)
);

NOR2x1_ASAP7_75t_SL g1233 ( 
.A(n_1227),
.B(n_1136),
.Y(n_1233)
);

INVxp67_ASAP7_75t_SL g1234 ( 
.A(n_1090),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1119),
.A2(n_1094),
.B(n_1111),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1221),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1090),
.A2(n_1226),
.B1(n_1086),
.B2(n_1207),
.Y(n_1237)
);

NAND2x1p5_ASAP7_75t_L g1238 ( 
.A(n_1227),
.B(n_1100),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1175),
.B(n_1183),
.Y(n_1239)
);

CKINVDCx8_ASAP7_75t_R g1240 ( 
.A(n_1097),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1218),
.B(n_1123),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1122),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_1206),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1110),
.B(n_1176),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1150),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1172),
.B(n_1138),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1176),
.B(n_1191),
.Y(n_1247)
);

INVx5_ASAP7_75t_L g1248 ( 
.A(n_1221),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1185),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1100),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1170),
.B(n_1213),
.Y(n_1251)
);

NAND2x1p5_ASAP7_75t_L g1252 ( 
.A(n_1227),
.B(n_1100),
.Y(n_1252)
);

NAND2x1p5_ASAP7_75t_L g1253 ( 
.A(n_1227),
.B(n_1143),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1094),
.A2(n_1111),
.B(n_1109),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1169),
.A2(n_1207),
.B1(n_1104),
.B2(n_1170),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1213),
.B(n_1189),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1084),
.A2(n_1199),
.B(n_1178),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1175),
.B(n_1183),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1091),
.Y(n_1259)
);

AND2x6_ASAP7_75t_L g1260 ( 
.A(n_1105),
.B(n_1114),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1187),
.B(n_1195),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1143),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1187),
.B(n_1195),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_SL g1264 ( 
.A(n_1141),
.B(n_1084),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1210),
.B(n_1211),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1143),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1193),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1222),
.B(n_1134),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1127),
.B(n_1131),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1209),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_SL g1271 ( 
.A1(n_1093),
.A2(n_1219),
.B(n_1199),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1222),
.B(n_1112),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1109),
.A2(n_1113),
.B(n_1124),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1196),
.B(n_1225),
.Y(n_1274)
);

OR2x6_ASAP7_75t_L g1275 ( 
.A(n_1159),
.B(n_1108),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1117),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1196),
.B(n_1225),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_1217),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1088),
.A2(n_1178),
.B(n_1219),
.C(n_1208),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1174),
.B(n_1192),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1216),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1117),
.Y(n_1282)
);

CKINVDCx8_ASAP7_75t_R g1283 ( 
.A(n_1098),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1089),
.B(n_1198),
.Y(n_1284)
);

INVx8_ASAP7_75t_L g1285 ( 
.A(n_1162),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1214),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1177),
.B(n_1157),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1148),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1116),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1130),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1092),
.B(n_1096),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1092),
.B(n_1116),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1151),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1149),
.A2(n_1160),
.B(n_1121),
.C(n_1208),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1177),
.A2(n_1107),
.B1(n_1160),
.B2(n_1149),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1164),
.A2(n_1180),
.B1(n_1200),
.B2(n_1118),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1091),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1173),
.B(n_1224),
.Y(n_1298)
);

NAND2x1p5_ASAP7_75t_L g1299 ( 
.A(n_1132),
.B(n_1155),
.Y(n_1299)
);

OAI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1161),
.A2(n_1201),
.B1(n_1197),
.B2(n_1120),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1214),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1129),
.B(n_1153),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1083),
.A2(n_1095),
.B(n_1142),
.Y(n_1303)
);

OR2x6_ASAP7_75t_L g1304 ( 
.A(n_1158),
.B(n_1168),
.Y(n_1304)
);

OAI321xp33_ASAP7_75t_L g1305 ( 
.A1(n_1087),
.A2(n_1125),
.A3(n_1154),
.B1(n_1153),
.B2(n_1163),
.C(n_1203),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1137),
.B(n_1099),
.Y(n_1306)
);

CKINVDCx11_ASAP7_75t_R g1307 ( 
.A(n_1165),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1146),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1173),
.B(n_1224),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1203),
.A2(n_1223),
.B1(n_1135),
.B2(n_1145),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1146),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1173),
.B(n_1224),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1152),
.Y(n_1313)
);

AND2x4_ASAP7_75t_SL g1314 ( 
.A(n_1156),
.B(n_1140),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1126),
.A2(n_1181),
.B1(n_1101),
.B2(n_1212),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1133),
.B(n_1182),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1133),
.B(n_1186),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1202),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1144),
.A2(n_1215),
.B(n_1190),
.C(n_1188),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1204),
.Y(n_1320)
);

INVx5_ASAP7_75t_L g1321 ( 
.A(n_1171),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1167),
.A2(n_1179),
.B(n_1205),
.Y(n_1322)
);

NOR2xp67_ASAP7_75t_L g1323 ( 
.A(n_1139),
.B(n_1147),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1184),
.A2(n_1103),
.B(n_1128),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1106),
.A2(n_1004),
.B1(n_1085),
.B2(n_1169),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1218),
.B(n_1123),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1206),
.Y(n_1327)
);

A2O1A1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1085),
.A2(n_1004),
.B(n_927),
.C(n_1170),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1085),
.A2(n_1004),
.B1(n_1090),
.B2(n_1166),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1085),
.B(n_1090),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1131),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1110),
.B(n_1176),
.Y(n_1332)
);

CKINVDCx6p67_ASAP7_75t_R g1333 ( 
.A(n_1216),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1085),
.A2(n_1004),
.B(n_927),
.C(n_1170),
.Y(n_1334)
);

BUFx4_ASAP7_75t_SL g1335 ( 
.A(n_1216),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1206),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1100),
.Y(n_1337)
);

BUFx12f_ASAP7_75t_L g1338 ( 
.A(n_1206),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1085),
.B(n_1090),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1141),
.B(n_1221),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1150),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1085),
.A2(n_1004),
.B1(n_1056),
.B2(n_927),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1115),
.Y(n_1343)
);

INVxp67_ASAP7_75t_SL g1344 ( 
.A(n_1085),
.Y(n_1344)
);

NAND2x1_ASAP7_75t_L g1345 ( 
.A(n_1142),
.B(n_762),
.Y(n_1345)
);

NAND2x1p5_ASAP7_75t_L g1346 ( 
.A(n_1227),
.B(n_746),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1102),
.Y(n_1347)
);

BUFx10_ASAP7_75t_L g1348 ( 
.A(n_1176),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1090),
.B(n_1225),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1085),
.B(n_927),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1085),
.B(n_1090),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1085),
.B(n_1090),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1115),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1102),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1150),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1221),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1119),
.A2(n_781),
.B(n_762),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1115),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1119),
.A2(n_781),
.B(n_762),
.Y(n_1359)
);

INVx4_ASAP7_75t_L g1360 ( 
.A(n_1221),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1085),
.A2(n_1004),
.B1(n_1090),
.B2(n_1166),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1085),
.B(n_1090),
.Y(n_1362)
);

INVx4_ASAP7_75t_L g1363 ( 
.A(n_1221),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1085),
.B(n_1090),
.Y(n_1364)
);

NOR2x1_ASAP7_75t_SL g1365 ( 
.A(n_1227),
.B(n_1027),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1115),
.Y(n_1366)
);

NAND2x1p5_ASAP7_75t_L g1367 ( 
.A(n_1227),
.B(n_746),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1085),
.A2(n_1004),
.B1(n_1090),
.B2(n_1166),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1110),
.B(n_1176),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1085),
.A2(n_1004),
.B(n_927),
.C(n_1170),
.Y(n_1370)
);

AO21x1_ASAP7_75t_L g1371 ( 
.A1(n_1232),
.A2(n_1237),
.B(n_1329),
.Y(n_1371)
);

CKINVDCx6p67_ASAP7_75t_R g1372 ( 
.A(n_1338),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1273),
.A2(n_1235),
.B(n_1254),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1242),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1275),
.B(n_1340),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1249),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1267),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_SL g1378 ( 
.A1(n_1350),
.A2(n_1344),
.B1(n_1251),
.B2(n_1295),
.Y(n_1378)
);

AOI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1256),
.A2(n_1265),
.B1(n_1342),
.B2(n_1246),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1245),
.Y(n_1380)
);

CKINVDCx6p67_ASAP7_75t_R g1381 ( 
.A(n_1243),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1255),
.A2(n_1295),
.B1(n_1361),
.B2(n_1368),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1330),
.A2(n_1362),
.B1(n_1339),
.B2(n_1364),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_SL g1384 ( 
.A(n_1281),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1270),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1255),
.B(n_1234),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1355),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1335),
.Y(n_1388)
);

BUFx2_ASAP7_75t_R g1389 ( 
.A(n_1230),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1285),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1346),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_1346),
.Y(n_1392)
);

INVxp33_ASAP7_75t_L g1393 ( 
.A(n_1241),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1367),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1287),
.B(n_1291),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1276),
.B(n_1282),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1345),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1329),
.A2(n_1361),
.B1(n_1368),
.B2(n_1237),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1328),
.A2(n_1370),
.B(n_1334),
.Y(n_1399)
);

AO21x1_ASAP7_75t_SL g1400 ( 
.A1(n_1298),
.A2(n_1309),
.B(n_1311),
.Y(n_1400)
);

INVx6_ASAP7_75t_L g1401 ( 
.A(n_1248),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1353),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1248),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1248),
.Y(n_1404)
);

OR2x6_ASAP7_75t_L g1405 ( 
.A(n_1271),
.B(n_1294),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1257),
.A2(n_1269),
.B1(n_1260),
.B2(n_1352),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1347),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1302),
.B(n_1325),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1358),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1285),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1354),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1348),
.Y(n_1412)
);

NAND3xp33_ASAP7_75t_L g1413 ( 
.A(n_1325),
.B(n_1351),
.C(n_1296),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1289),
.B(n_1290),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1304),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1349),
.B(n_1239),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1274),
.A2(n_1263),
.B1(n_1261),
.B2(n_1277),
.Y(n_1417)
);

AOI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1357),
.A2(n_1359),
.B(n_1310),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1258),
.B(n_1326),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1257),
.A2(n_1260),
.B1(n_1275),
.B2(n_1231),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1289),
.Y(n_1421)
);

INVx4_ASAP7_75t_L g1422 ( 
.A(n_1340),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1304),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1319),
.A2(n_1315),
.B(n_1288),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1260),
.A2(n_1275),
.B1(n_1366),
.B2(n_1231),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1312),
.B(n_1292),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1305),
.A2(n_1316),
.B(n_1320),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1260),
.A2(n_1366),
.B1(n_1343),
.B2(n_1300),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1343),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1293),
.Y(n_1430)
);

OAI22xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1264),
.A2(n_1286),
.B1(n_1331),
.B2(n_1301),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1340),
.B(n_1259),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1278),
.A2(n_1341),
.B1(n_1284),
.B2(n_1279),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1317),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1264),
.A2(n_1233),
.B1(n_1284),
.B2(n_1247),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1247),
.B(n_1229),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1240),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1308),
.Y(n_1438)
);

BUFx12f_ASAP7_75t_L g1439 ( 
.A(n_1327),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1297),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1318),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1238),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1244),
.A2(n_1332),
.B1(n_1369),
.B2(n_1272),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1306),
.Y(n_1444)
);

BUFx4f_ASAP7_75t_SL g1445 ( 
.A(n_1333),
.Y(n_1445)
);

CKINVDCx8_ASAP7_75t_R g1446 ( 
.A(n_1244),
.Y(n_1446)
);

BUFx12f_ASAP7_75t_L g1447 ( 
.A(n_1336),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1306),
.B(n_1259),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1332),
.A2(n_1369),
.B1(n_1272),
.B2(n_1348),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1252),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1313),
.A2(n_1322),
.B(n_1299),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1252),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1280),
.A2(n_1268),
.B1(n_1281),
.B2(n_1304),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1268),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1253),
.Y(n_1455)
);

INVx11_ASAP7_75t_L g1456 ( 
.A(n_1283),
.Y(n_1456)
);

NAND2x1p5_ASAP7_75t_L g1457 ( 
.A(n_1360),
.B(n_1363),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1253),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1228),
.B(n_1236),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1337),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1280),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_SL g1462 ( 
.A1(n_1281),
.A2(n_1314),
.B1(n_1365),
.B2(n_1363),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1322),
.Y(n_1463)
);

INVxp33_ASAP7_75t_L g1464 ( 
.A(n_1307),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1250),
.A2(n_1262),
.B1(n_1266),
.B2(n_1228),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1299),
.A2(n_1236),
.B(n_1356),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1356),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1360),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1321),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1346),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_SL g1471 ( 
.A1(n_1292),
.A2(n_1294),
.B(n_1164),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1350),
.B(n_1085),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1255),
.B(n_1234),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1234),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1350),
.A2(n_1004),
.B1(n_1085),
.B2(n_927),
.Y(n_1475)
);

AOI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1323),
.A2(n_1119),
.B(n_1324),
.Y(n_1476)
);

AO21x2_ASAP7_75t_L g1477 ( 
.A1(n_1324),
.A2(n_1118),
.B(n_1303),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1350),
.A2(n_1004),
.B1(n_1085),
.B2(n_927),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1234),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1245),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1245),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1348),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1245),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1242),
.Y(n_1484)
);

BUFx12f_ASAP7_75t_L g1485 ( 
.A(n_1230),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1242),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1242),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1298),
.B(n_1309),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1350),
.A2(n_1004),
.B1(n_1085),
.B2(n_927),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1255),
.B(n_1234),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1350),
.B(n_1085),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1346),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1350),
.A2(n_1085),
.B1(n_927),
.B2(n_1004),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_SL g1494 ( 
.A(n_1281),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1350),
.A2(n_1085),
.B1(n_1004),
.B2(n_1330),
.Y(n_1495)
);

BUFx10_ASAP7_75t_L g1496 ( 
.A(n_1301),
.Y(n_1496)
);

INVx8_ASAP7_75t_L g1497 ( 
.A(n_1384),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1426),
.B(n_1386),
.Y(n_1498)
);

INVx3_ASAP7_75t_SL g1499 ( 
.A(n_1388),
.Y(n_1499)
);

BUFx2_ASAP7_75t_SL g1500 ( 
.A(n_1384),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1437),
.Y(n_1501)
);

OR2x6_ASAP7_75t_L g1502 ( 
.A(n_1405),
.B(n_1415),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_SL g1503 ( 
.A1(n_1495),
.A2(n_1399),
.B1(n_1413),
.B2(n_1405),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1417),
.B(n_1383),
.Y(n_1504)
);

INVx5_ASAP7_75t_L g1505 ( 
.A(n_1405),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1488),
.B(n_1434),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1388),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1415),
.B(n_1423),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1438),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1488),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1386),
.B(n_1473),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1480),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1426),
.B(n_1473),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1416),
.B(n_1419),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1430),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1375),
.B(n_1448),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1463),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1490),
.B(n_1395),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1463),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1441),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1476),
.A2(n_1424),
.B(n_1418),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1481),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1490),
.B(n_1408),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1427),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1395),
.B(n_1408),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1374),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1378),
.B(n_1379),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1387),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1427),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1427),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1375),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1466),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1382),
.B(n_1398),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1376),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1377),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1472),
.B(n_1491),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1466),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1385),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1414),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1415),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1474),
.B(n_1479),
.Y(n_1541)
);

OR2x6_ASAP7_75t_L g1542 ( 
.A(n_1405),
.B(n_1375),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1414),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1421),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1437),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1448),
.B(n_1444),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1402),
.Y(n_1547)
);

INVx8_ASAP7_75t_L g1548 ( 
.A(n_1384),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1444),
.B(n_1432),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1396),
.B(n_1400),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1409),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1493),
.A2(n_1489),
.B1(n_1475),
.B2(n_1478),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1396),
.B(n_1400),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1393),
.B(n_1454),
.Y(n_1554)
);

AO21x2_ASAP7_75t_L g1555 ( 
.A1(n_1471),
.A2(n_1477),
.B(n_1371),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1451),
.A2(n_1397),
.B(n_1373),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1484),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1371),
.B(n_1406),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1486),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1487),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1429),
.Y(n_1561)
);

NAND2xp33_ASAP7_75t_SL g1562 ( 
.A(n_1494),
.B(n_1464),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1420),
.B(n_1393),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1380),
.B(n_1483),
.Y(n_1564)
);

INVx8_ASAP7_75t_L g1565 ( 
.A(n_1494),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1471),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1477),
.Y(n_1567)
);

AO21x2_ASAP7_75t_L g1568 ( 
.A1(n_1469),
.A2(n_1436),
.B(n_1440),
.Y(n_1568)
);

INVxp67_ASAP7_75t_R g1569 ( 
.A(n_1433),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1407),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1411),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1387),
.Y(n_1572)
);

OR2x6_ASAP7_75t_L g1573 ( 
.A(n_1422),
.B(n_1401),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1425),
.B(n_1428),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1422),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1392),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1432),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1461),
.B(n_1432),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1492),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1467),
.Y(n_1580)
);

NAND2xp33_ASAP7_75t_SL g1581 ( 
.A(n_1533),
.B(n_1494),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1550),
.B(n_1435),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1517),
.B(n_1453),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1553),
.B(n_1460),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1567),
.B(n_1460),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1568),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1519),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1510),
.B(n_1431),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1524),
.B(n_1458),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1541),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1515),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1505),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1529),
.B(n_1482),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1529),
.B(n_1459),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1510),
.B(n_1462),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1508),
.B(n_1390),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1530),
.B(n_1412),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1509),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1530),
.B(n_1459),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1555),
.B(n_1459),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1527),
.A2(n_1464),
.B1(n_1449),
.B2(n_1381),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1508),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1504),
.B(n_1455),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1555),
.B(n_1470),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1552),
.A2(n_1533),
.B1(n_1503),
.B2(n_1558),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1498),
.B(n_1394),
.Y(n_1606)
);

NAND2x1p5_ASAP7_75t_L g1607 ( 
.A(n_1505),
.B(n_1403),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1506),
.B(n_1498),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1506),
.B(n_1513),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1508),
.B(n_1532),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1532),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1568),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1541),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1513),
.B(n_1450),
.Y(n_1614)
);

AOI21xp33_ASAP7_75t_L g1615 ( 
.A1(n_1558),
.A2(n_1442),
.B(n_1452),
.Y(n_1615)
);

BUFx2_ASAP7_75t_SL g1616 ( 
.A(n_1505),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1509),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1525),
.B(n_1391),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1518),
.B(n_1391),
.Y(n_1619)
);

OAI221xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1605),
.A2(n_1601),
.B1(n_1523),
.B2(n_1574),
.C(n_1588),
.Y(n_1620)
);

NAND4xp25_ASAP7_75t_L g1621 ( 
.A(n_1605),
.B(n_1536),
.C(n_1514),
.D(n_1564),
.Y(n_1621)
);

NAND3xp33_ASAP7_75t_SL g1622 ( 
.A(n_1601),
.B(n_1562),
.C(n_1545),
.Y(n_1622)
);

NOR2xp67_ASAP7_75t_L g1623 ( 
.A(n_1586),
.B(n_1537),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1608),
.B(n_1523),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1603),
.B(n_1501),
.Y(n_1625)
);

OAI221xp5_ASAP7_75t_SL g1626 ( 
.A1(n_1588),
.A2(n_1574),
.B1(n_1511),
.B2(n_1563),
.C(n_1542),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1582),
.A2(n_1563),
.B1(n_1542),
.B2(n_1549),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1594),
.B(n_1518),
.Y(n_1628)
);

INVxp67_ASAP7_75t_L g1629 ( 
.A(n_1590),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1603),
.A2(n_1569),
.B1(n_1446),
.B2(n_1505),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1608),
.B(n_1609),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1594),
.B(n_1540),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1599),
.B(n_1540),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1609),
.B(n_1512),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1598),
.B(n_1522),
.Y(n_1635)
);

OAI221xp5_ASAP7_75t_SL g1636 ( 
.A1(n_1595),
.A2(n_1542),
.B1(n_1502),
.B2(n_1554),
.C(n_1566),
.Y(n_1636)
);

OAI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1581),
.A2(n_1443),
.B1(n_1572),
.B2(n_1551),
.C(n_1547),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1598),
.B(n_1539),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1581),
.B(n_1531),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1617),
.B(n_1543),
.Y(n_1640)
);

OA21x2_ASAP7_75t_L g1641 ( 
.A1(n_1586),
.A2(n_1521),
.B(n_1556),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1595),
.A2(n_1569),
.B1(n_1446),
.B2(n_1505),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1583),
.A2(n_1502),
.B1(n_1531),
.B2(n_1573),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_SL g1644 ( 
.A1(n_1582),
.A2(n_1516),
.B(n_1549),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1618),
.B(n_1546),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1618),
.B(n_1546),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1617),
.B(n_1544),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1602),
.B(n_1546),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1602),
.B(n_1568),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1602),
.B(n_1502),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1590),
.B(n_1561),
.Y(n_1651)
);

NOR3xp33_ASAP7_75t_L g1652 ( 
.A(n_1615),
.B(n_1575),
.C(n_1566),
.Y(n_1652)
);

AOI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1615),
.A2(n_1580),
.B1(n_1520),
.B2(n_1559),
.C(n_1557),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1613),
.B(n_1520),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1613),
.B(n_1526),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1607),
.A2(n_1577),
.B(n_1578),
.Y(n_1656)
);

OAI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1583),
.A2(n_1528),
.B1(n_1465),
.B2(n_1500),
.C(n_1575),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1614),
.B(n_1526),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_R g1659 ( 
.A(n_1583),
.B(n_1507),
.Y(n_1659)
);

OAI21xp33_ASAP7_75t_L g1660 ( 
.A1(n_1614),
.A2(n_1559),
.B(n_1560),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1616),
.A2(n_1565),
.B1(n_1497),
.B2(n_1548),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1606),
.B(n_1534),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1591),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1596),
.B(n_1545),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1606),
.B(n_1534),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1612),
.B(n_1570),
.C(n_1571),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1606),
.B(n_1535),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1602),
.B(n_1502),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1596),
.A2(n_1410),
.B1(n_1390),
.B2(n_1548),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1619),
.B(n_1535),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1607),
.A2(n_1573),
.B(n_1565),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1619),
.B(n_1538),
.Y(n_1672)
);

AOI21xp33_ASAP7_75t_L g1673 ( 
.A1(n_1604),
.A2(n_1579),
.B(n_1576),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1663),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1663),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1623),
.B(n_1610),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1641),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1629),
.B(n_1587),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1624),
.B(n_1587),
.Y(n_1679)
);

INVx4_ASAP7_75t_L g1680 ( 
.A(n_1650),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1628),
.B(n_1600),
.Y(n_1681)
);

INVx5_ASAP7_75t_L g1682 ( 
.A(n_1649),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1649),
.Y(n_1683)
);

OR2x2_ASAP7_75t_SL g1684 ( 
.A(n_1622),
.B(n_1592),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1655),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1641),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1623),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1654),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1666),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1659),
.B(n_1592),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1666),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1651),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_1647),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1631),
.B(n_1604),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1632),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1632),
.Y(n_1696)
);

AND2x4_ASAP7_75t_SL g1697 ( 
.A(n_1650),
.B(n_1592),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1633),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1638),
.B(n_1593),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1668),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1668),
.B(n_1610),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1640),
.B(n_1593),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1662),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1645),
.B(n_1585),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1665),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1660),
.B(n_1589),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1667),
.B(n_1593),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1670),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1671),
.B(n_1611),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1674),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1689),
.B(n_1635),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1697),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1692),
.B(n_1634),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1690),
.B(n_1661),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1693),
.B(n_1625),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1692),
.B(n_1646),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1674),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1675),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1674),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1680),
.B(n_1648),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1680),
.B(n_1648),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1689),
.B(n_1672),
.Y(n_1722)
);

NAND2x1p5_ASAP7_75t_L g1723 ( 
.A(n_1690),
.B(n_1592),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1675),
.Y(n_1724)
);

AOI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1691),
.A2(n_1620),
.B1(n_1621),
.B2(n_1626),
.C(n_1673),
.Y(n_1725)
);

BUFx3_ASAP7_75t_L g1726 ( 
.A(n_1693),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1691),
.B(n_1658),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1680),
.B(n_1644),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1675),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1680),
.B(n_1681),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1675),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1680),
.B(n_1644),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1676),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1677),
.Y(n_1734)
);

NAND3xp33_ASAP7_75t_L g1735 ( 
.A(n_1688),
.B(n_1621),
.C(n_1653),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1681),
.B(n_1584),
.Y(n_1736)
);

AOI32xp33_ASAP7_75t_L g1737 ( 
.A1(n_1697),
.A2(n_1652),
.A3(n_1642),
.B1(n_1630),
.B2(n_1657),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1688),
.B(n_1685),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1681),
.B(n_1584),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1694),
.B(n_1597),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1695),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1695),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1694),
.B(n_1703),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1683),
.B(n_1584),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1703),
.B(n_1597),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1677),
.Y(n_1746)
);

NAND2x1p5_ASAP7_75t_L g1747 ( 
.A(n_1682),
.B(n_1592),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1696),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1683),
.B(n_1656),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1696),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1698),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1707),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1683),
.B(n_1656),
.Y(n_1753)
);

INVxp67_ASAP7_75t_SL g1754 ( 
.A(n_1726),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1728),
.B(n_1683),
.Y(n_1755)
);

NAND2x1p5_ASAP7_75t_L g1756 ( 
.A(n_1726),
.B(n_1639),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1710),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1712),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1735),
.A2(n_1685),
.B1(n_1705),
.B2(n_1708),
.C(n_1679),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1725),
.B(n_1705),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1710),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1752),
.B(n_1699),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1727),
.B(n_1699),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1717),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1717),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1711),
.B(n_1708),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1728),
.B(n_1701),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1727),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1719),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1711),
.B(n_1703),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1722),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1715),
.B(n_1700),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1712),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1713),
.B(n_1700),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1719),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1722),
.B(n_1700),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1718),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1748),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1748),
.Y(n_1779)
);

OAI21xp33_ASAP7_75t_L g1780 ( 
.A1(n_1737),
.A2(n_1636),
.B(n_1706),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1750),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1714),
.A2(n_1664),
.B(n_1643),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1741),
.B(n_1699),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1732),
.B(n_1749),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1716),
.B(n_1738),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1718),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1750),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1741),
.B(n_1702),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1732),
.B(n_1701),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1736),
.B(n_1704),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1742),
.B(n_1702),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1751),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1742),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1751),
.Y(n_1794)
);

NOR2x1_ASAP7_75t_L g1795 ( 
.A(n_1749),
.B(n_1678),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1736),
.B(n_1704),
.Y(n_1796)
);

INVxp67_ASAP7_75t_L g1797 ( 
.A(n_1720),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1724),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1730),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1758),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1765),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1777),
.Y(n_1802)
);

AO21x2_ASAP7_75t_L g1803 ( 
.A1(n_1798),
.A2(n_1746),
.B(n_1734),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1763),
.B(n_1743),
.Y(n_1804)
);

BUFx3_ASAP7_75t_L g1805 ( 
.A(n_1758),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1756),
.B(n_1753),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1777),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1780),
.A2(n_1753),
.B1(n_1637),
.B2(n_1730),
.Y(n_1808)
);

INVxp67_ASAP7_75t_SL g1809 ( 
.A(n_1754),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1759),
.B(n_1743),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1786),
.Y(n_1811)
);

INVx3_ASAP7_75t_SL g1812 ( 
.A(n_1773),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1756),
.B(n_1733),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1786),
.Y(n_1814)
);

AND2x2_ASAP7_75t_SL g1815 ( 
.A(n_1760),
.B(n_1684),
.Y(n_1815)
);

INVx1_ASAP7_75t_SL g1816 ( 
.A(n_1773),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1793),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1765),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1756),
.B(n_1733),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1769),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1769),
.Y(n_1821)
);

CKINVDCx14_ASAP7_75t_R g1822 ( 
.A(n_1784),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1757),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1768),
.B(n_1740),
.Y(n_1824)
);

NOR2x1_ASAP7_75t_L g1825 ( 
.A(n_1795),
.B(n_1733),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1763),
.B(n_1724),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_1784),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1761),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1764),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1771),
.B(n_1740),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1775),
.Y(n_1831)
);

INVx1_ASAP7_75t_SL g1832 ( 
.A(n_1772),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1762),
.B(n_1783),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1785),
.B(n_1745),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1762),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1767),
.B(n_1747),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1755),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1809),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1809),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1822),
.B(n_1755),
.Y(n_1840)
);

AOI221xp5_ASAP7_75t_L g1841 ( 
.A1(n_1810),
.A2(n_1782),
.B1(n_1797),
.B2(n_1799),
.C(n_1774),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1815),
.A2(n_1776),
.B1(n_1789),
.B2(n_1767),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1815),
.A2(n_1766),
.B(n_1770),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1801),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1805),
.Y(n_1845)
);

OAI32xp33_ASAP7_75t_L g1846 ( 
.A1(n_1810),
.A2(n_1747),
.A3(n_1723),
.B1(n_1783),
.B2(n_1791),
.Y(n_1846)
);

O2A1O1Ixp33_ASAP7_75t_L g1847 ( 
.A1(n_1817),
.A2(n_1812),
.B(n_1832),
.C(n_1816),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1827),
.B(n_1789),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1801),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1815),
.A2(n_1709),
.B1(n_1723),
.B2(n_1697),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1825),
.A2(n_1723),
.B(n_1747),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1805),
.Y(n_1852)
);

AOI21xp33_ASAP7_75t_SL g1853 ( 
.A1(n_1812),
.A2(n_1499),
.B(n_1507),
.Y(n_1853)
);

O2A1O1Ixp5_ASAP7_75t_L g1854 ( 
.A1(n_1806),
.A2(n_1791),
.B(n_1788),
.C(n_1778),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1806),
.B(n_1788),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1827),
.B(n_1372),
.Y(n_1856)
);

OAI211xp5_ASAP7_75t_SL g1857 ( 
.A1(n_1832),
.A2(n_1737),
.B(n_1798),
.C(n_1781),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1837),
.B(n_1790),
.Y(n_1858)
);

OAI221xp5_ASAP7_75t_L g1859 ( 
.A1(n_1808),
.A2(n_1794),
.B1(n_1792),
.B2(n_1787),
.C(n_1779),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1817),
.Y(n_1860)
);

OAI21xp33_ASAP7_75t_L g1861 ( 
.A1(n_1808),
.A2(n_1627),
.B(n_1796),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1837),
.B(n_1739),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1812),
.B(n_1800),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1806),
.B(n_1720),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1820),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_SL g1866 ( 
.A1(n_1840),
.A2(n_1805),
.B1(n_1836),
.B2(n_1816),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1856),
.B(n_1800),
.Y(n_1867)
);

AOI222xp33_ASAP7_75t_L g1868 ( 
.A1(n_1857),
.A2(n_1825),
.B1(n_1824),
.B2(n_1830),
.C1(n_1835),
.C2(n_1834),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1853),
.B(n_1824),
.Y(n_1869)
);

NOR2xp67_ASAP7_75t_SL g1870 ( 
.A(n_1860),
.B(n_1439),
.Y(n_1870)
);

OAI222xp33_ASAP7_75t_L g1871 ( 
.A1(n_1842),
.A2(n_1833),
.B1(n_1830),
.B2(n_1835),
.C1(n_1804),
.C2(n_1813),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1856),
.B(n_1838),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1860),
.B(n_1852),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1863),
.B(n_1835),
.Y(n_1874)
);

HB1xp67_ASAP7_75t_L g1875 ( 
.A(n_1845),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1863),
.B(n_1833),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1855),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1859),
.A2(n_1684),
.B1(n_1833),
.B2(n_1682),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1864),
.B(n_1836),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1839),
.B(n_1823),
.Y(n_1880)
);

INVxp67_ASAP7_75t_L g1881 ( 
.A(n_1845),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1855),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1847),
.B(n_1439),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1864),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1848),
.B(n_1836),
.Y(n_1885)
);

NAND2x1_ASAP7_75t_L g1886 ( 
.A(n_1850),
.B(n_1813),
.Y(n_1886)
);

AND2x4_ASAP7_75t_SL g1887 ( 
.A(n_1865),
.B(n_1381),
.Y(n_1887)
);

OAI21xp5_ASAP7_75t_SL g1888 ( 
.A1(n_1868),
.A2(n_1841),
.B(n_1843),
.Y(n_1888)
);

OAI211xp5_ASAP7_75t_L g1889 ( 
.A1(n_1866),
.A2(n_1846),
.B(n_1861),
.C(n_1851),
.Y(n_1889)
);

AOI21xp33_ASAP7_75t_SL g1890 ( 
.A1(n_1883),
.A2(n_1499),
.B(n_1858),
.Y(n_1890)
);

OAI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1886),
.A2(n_1862),
.B1(n_1804),
.B2(n_1682),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1881),
.B(n_1844),
.Y(n_1892)
);

OAI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1871),
.A2(n_1854),
.B(n_1819),
.Y(n_1893)
);

AOI211xp5_ASAP7_75t_SL g1894 ( 
.A1(n_1883),
.A2(n_1849),
.B(n_1819),
.C(n_1813),
.Y(n_1894)
);

OAI322xp33_ASAP7_75t_L g1895 ( 
.A1(n_1873),
.A2(n_1820),
.A3(n_1831),
.B1(n_1829),
.B2(n_1828),
.C1(n_1823),
.C2(n_1804),
.Y(n_1895)
);

AOI311xp33_ASAP7_75t_L g1896 ( 
.A1(n_1872),
.A2(n_1831),
.A3(n_1829),
.B(n_1828),
.C(n_1834),
.Y(n_1896)
);

AOI211x1_ASAP7_75t_SL g1897 ( 
.A1(n_1869),
.A2(n_1821),
.B(n_1818),
.C(n_1807),
.Y(n_1897)
);

AOI211xp5_ASAP7_75t_SL g1898 ( 
.A1(n_1867),
.A2(n_1819),
.B(n_1445),
.C(n_1807),
.Y(n_1898)
);

NOR3xp33_ASAP7_75t_L g1899 ( 
.A(n_1872),
.B(n_1821),
.C(n_1818),
.Y(n_1899)
);

AOI222xp33_ASAP7_75t_L g1900 ( 
.A1(n_1874),
.A2(n_1821),
.B1(n_1818),
.B2(n_1807),
.C1(n_1814),
.C2(n_1811),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1893),
.A2(n_1867),
.B1(n_1882),
.B2(n_1877),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1888),
.B(n_1875),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1894),
.B(n_1875),
.Y(n_1903)
);

NOR3x1_ASAP7_75t_L g1904 ( 
.A(n_1889),
.B(n_1876),
.C(n_1880),
.Y(n_1904)
);

NAND3xp33_ASAP7_75t_L g1905 ( 
.A(n_1899),
.B(n_1870),
.C(n_1884),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1890),
.B(n_1887),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1892),
.B(n_1885),
.Y(n_1907)
);

NOR2x1_ASAP7_75t_L g1908 ( 
.A(n_1895),
.B(n_1878),
.Y(n_1908)
);

NAND3xp33_ASAP7_75t_L g1909 ( 
.A(n_1899),
.B(n_1879),
.C(n_1811),
.Y(n_1909)
);

NAND3xp33_ASAP7_75t_L g1910 ( 
.A(n_1896),
.B(n_1811),
.C(n_1802),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1900),
.Y(n_1911)
);

NOR5xp2_ASAP7_75t_L g1912 ( 
.A(n_1910),
.B(n_1897),
.C(n_1898),
.D(n_1891),
.E(n_1687),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_L g1913 ( 
.A1(n_1911),
.A2(n_1802),
.B1(n_1814),
.B2(n_1826),
.Y(n_1913)
);

NOR2x1_ASAP7_75t_L g1914 ( 
.A(n_1902),
.B(n_1802),
.Y(n_1914)
);

NAND3xp33_ASAP7_75t_SL g1915 ( 
.A(n_1901),
.B(n_1389),
.C(n_1814),
.Y(n_1915)
);

AOI221xp5_ASAP7_75t_L g1916 ( 
.A1(n_1903),
.A2(n_1905),
.B1(n_1909),
.B2(n_1907),
.C(n_1906),
.Y(n_1916)
);

XOR2x2_ASAP7_75t_L g1917 ( 
.A(n_1908),
.B(n_1499),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1915),
.B(n_1447),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1914),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1917),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1913),
.Y(n_1921)
);

AOI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1916),
.A2(n_1904),
.B1(n_1485),
.B2(n_1447),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1912),
.B(n_1826),
.Y(n_1923)
);

NOR2xp67_ASAP7_75t_L g1924 ( 
.A(n_1915),
.B(n_1485),
.Y(n_1924)
);

NAND4xp25_ASAP7_75t_SL g1925 ( 
.A(n_1922),
.B(n_1826),
.C(n_1456),
.D(n_1721),
.Y(n_1925)
);

INVxp33_ASAP7_75t_L g1926 ( 
.A(n_1918),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1919),
.Y(n_1927)
);

AND3x4_ASAP7_75t_L g1928 ( 
.A(n_1924),
.B(n_1456),
.C(n_1496),
.Y(n_1928)
);

NOR2x1_ASAP7_75t_L g1929 ( 
.A(n_1921),
.B(n_1803),
.Y(n_1929)
);

NAND3xp33_ASAP7_75t_L g1930 ( 
.A(n_1920),
.B(n_1687),
.C(n_1734),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1927),
.B(n_1923),
.Y(n_1931)
);

NOR3xp33_ASAP7_75t_SL g1932 ( 
.A(n_1925),
.B(n_1496),
.C(n_1669),
.Y(n_1932)
);

INVx4_ASAP7_75t_L g1933 ( 
.A(n_1928),
.Y(n_1933)
);

NOR3xp33_ASAP7_75t_L g1934 ( 
.A(n_1930),
.B(n_1929),
.C(n_1926),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1931),
.A2(n_1933),
.B1(n_1934),
.B2(n_1932),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1931),
.B(n_1803),
.Y(n_1936)
);

AOI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1935),
.A2(n_1803),
.B1(n_1746),
.B2(n_1721),
.C(n_1729),
.Y(n_1937)
);

OAI211xp5_ASAP7_75t_L g1938 ( 
.A1(n_1937),
.A2(n_1936),
.B(n_1496),
.C(n_1497),
.Y(n_1938)
);

OA21x2_ASAP7_75t_L g1939 ( 
.A1(n_1937),
.A2(n_1731),
.B(n_1729),
.Y(n_1939)
);

AOI21x1_ASAP7_75t_L g1940 ( 
.A1(n_1938),
.A2(n_1803),
.B(n_1731),
.Y(n_1940)
);

AOI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1939),
.A2(n_1744),
.B1(n_1709),
.B2(n_1497),
.Y(n_1941)
);

OAI21xp5_ASAP7_75t_SL g1942 ( 
.A1(n_1940),
.A2(n_1404),
.B(n_1457),
.Y(n_1942)
);

AOI222xp33_ASAP7_75t_L g1943 ( 
.A1(n_1942),
.A2(n_1941),
.B1(n_1744),
.B2(n_1548),
.C1(n_1497),
.C2(n_1565),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1943),
.A2(n_1565),
.B1(n_1548),
.B2(n_1497),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1944),
.A2(n_1565),
.B1(n_1548),
.B2(n_1686),
.Y(n_1945)
);

AOI211xp5_ASAP7_75t_L g1946 ( 
.A1(n_1945),
.A2(n_1404),
.B(n_1468),
.C(n_1678),
.Y(n_1946)
);


endmodule