module fake_netlist_1_2580_n_669 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_669);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_669;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_535;
wire n_225;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_75), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_68), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_8), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_43), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_58), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_61), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_72), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_27), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_47), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_15), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_54), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_62), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_41), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_44), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_18), .Y(n_91) );
INVxp33_ASAP7_75t_SL g92 ( .A(n_17), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_11), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_55), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_30), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_51), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_66), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_65), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_2), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_38), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_16), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_6), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_15), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_0), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_34), .Y(n_105) );
INVx3_ASAP7_75t_L g106 ( .A(n_32), .Y(n_106) );
XNOR2xp5_ASAP7_75t_L g107 ( .A(n_71), .B(n_29), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_31), .Y(n_108) );
OR2x2_ASAP7_75t_L g109 ( .A(n_64), .B(n_36), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_59), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_9), .Y(n_111) );
BUFx2_ASAP7_75t_SL g112 ( .A(n_56), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_63), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_17), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_70), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_74), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_48), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_26), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_35), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_69), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_23), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_33), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_11), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_106), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_88), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_88), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_90), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_121), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_106), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_106), .B(n_0), .Y(n_131) );
BUFx2_ASAP7_75t_L g132 ( .A(n_79), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_82), .B(n_1), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_90), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_123), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_121), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_123), .B(n_1), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_122), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_92), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_97), .Y(n_140) );
BUFx8_ASAP7_75t_L g141 ( .A(n_109), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_121), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_86), .B(n_3), .Y(n_143) );
NAND2xp33_ASAP7_75t_SL g144 ( .A(n_87), .B(n_4), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_122), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_77), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_78), .Y(n_147) );
NOR2xp33_ASAP7_75t_SL g148 ( .A(n_105), .B(n_25), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_86), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_80), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_93), .B(n_5), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_81), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_93), .B(n_5), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_83), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_95), .Y(n_157) );
OAI22xp5_ASAP7_75t_L g158 ( .A1(n_92), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_96), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_98), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_101), .B(n_7), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_121), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_100), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_108), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_103), .B(n_9), .Y(n_165) );
INVx5_ASAP7_75t_L g166 ( .A(n_162), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_129), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_129), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_129), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_132), .B(n_105), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_124), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_124), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_130), .Y(n_174) );
INVx1_ASAP7_75t_SL g175 ( .A(n_132), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_140), .B(n_89), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_129), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_136), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_140), .B(n_111), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_136), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_146), .B(n_89), .Y(n_182) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_143), .B(n_109), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_139), .A2(n_102), .B1(n_87), .B2(n_91), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_149), .B(n_104), .Y(n_185) );
OR2x2_ASAP7_75t_L g186 ( .A(n_128), .B(n_99), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_130), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_146), .B(n_94), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_143), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_143), .Y(n_190) );
INVx1_ASAP7_75t_SL g191 ( .A(n_135), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_125), .B(n_126), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_136), .Y(n_195) );
OR2x2_ASAP7_75t_L g196 ( .A(n_137), .B(n_114), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_136), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_154), .A2(n_102), .B1(n_94), .B2(n_107), .Y(n_198) );
OR2x6_ASAP7_75t_L g199 ( .A(n_158), .B(n_112), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_154), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_147), .B(n_115), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_142), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_154), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_147), .B(n_113), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_142), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_133), .B(n_112), .Y(n_206) );
AND2x2_ASAP7_75t_SL g207 ( .A(n_161), .B(n_116), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_142), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_161), .B(n_119), .Y(n_209) );
BUFx10_ASAP7_75t_L g210 ( .A(n_161), .Y(n_210) );
OAI21xp33_ASAP7_75t_L g211 ( .A1(n_125), .A2(n_118), .B(n_117), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_126), .B(n_84), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_162), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_151), .B(n_110), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_161), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_142), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_134), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_165), .B(n_120), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_165), .Y(n_219) );
INVxp67_ASAP7_75t_SL g220 ( .A(n_141), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_165), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_142), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_134), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_127), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_162), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_187), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_175), .Y(n_227) );
INVx5_ASAP7_75t_L g228 ( .A(n_210), .Y(n_228) );
BUFx3_ASAP7_75t_L g229 ( .A(n_187), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_188), .B(n_141), .Y(n_230) );
INVx1_ASAP7_75t_SL g231 ( .A(n_175), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_187), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_178), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_215), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_203), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_182), .B(n_141), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_215), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_198), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_217), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_189), .A2(n_138), .B(n_145), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_215), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_217), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_218), .B(n_165), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_178), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_178), .Y(n_245) );
OR2x6_ASAP7_75t_L g246 ( .A(n_183), .B(n_152), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_212), .B(n_152), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_207), .A2(n_151), .B1(n_159), .B2(n_157), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_178), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_221), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_218), .B(n_156), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_223), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_191), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_207), .A2(n_159), .B1(n_157), .B2(n_156), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_210), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_221), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_191), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_212), .B(n_138), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_218), .B(n_145), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_207), .B(n_127), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_170), .B(n_153), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_223), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_218), .B(n_164), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_190), .Y(n_264) );
AND2x4_ASAP7_75t_SL g265 ( .A(n_210), .B(n_164), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_176), .B(n_163), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_190), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_221), .A2(n_209), .B1(n_192), .B2(n_200), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_209), .B(n_163), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_183), .B(n_160), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_203), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_190), .Y(n_272) );
AOI21xp33_ASAP7_75t_L g273 ( .A1(n_206), .A2(n_148), .B(n_107), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_190), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_210), .Y(n_275) );
BUFx4f_ASAP7_75t_L g276 ( .A(n_183), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_198), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_220), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_185), .B(n_160), .Y(n_279) );
INVx3_ASAP7_75t_L g280 ( .A(n_203), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_184), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_224), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_224), .Y(n_283) );
OAI21xp33_ASAP7_75t_L g284 ( .A1(n_193), .A2(n_155), .B(n_153), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_213), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_206), .B(n_155), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_193), .B(n_131), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_203), .Y(n_288) );
INVx4_ASAP7_75t_L g289 ( .A(n_228), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_246), .A2(n_199), .B1(n_219), .B2(n_209), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_227), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_257), .B(n_185), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_275), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_231), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_282), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_233), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_233), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_260), .B(n_196), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_263), .A2(n_186), .B(n_196), .C(n_199), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_253), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_257), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_282), .Y(n_302) );
INVx4_ASAP7_75t_L g303 ( .A(n_228), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_246), .B(n_219), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_283), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_283), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_246), .A2(n_199), .B1(n_219), .B2(n_209), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_246), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_228), .Y(n_309) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_286), .A2(n_189), .B(n_192), .C(n_200), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_246), .B(n_219), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_236), .B(n_180), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_227), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_278), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_244), .Y(n_315) );
INVx4_ASAP7_75t_L g316 ( .A(n_228), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_260), .B(n_180), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_264), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_238), .A2(n_184), .B1(n_277), .B2(n_247), .C(n_279), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_228), .Y(n_320) );
INVx4_ASAP7_75t_SL g321 ( .A(n_275), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_270), .B(n_199), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_264), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_278), .Y(n_324) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_276), .B(n_171), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_270), .B(n_204), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_240), .A2(n_214), .B(n_171), .Y(n_327) );
BUFx4f_ASAP7_75t_SL g328 ( .A(n_281), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_276), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g330 ( .A1(n_238), .A2(n_199), .B1(n_186), .B2(n_174), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_244), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_251), .B(n_201), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_251), .B(n_211), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_237), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_237), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_266), .A2(n_211), .B(n_173), .C(n_174), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_251), .B(n_173), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_301), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_295), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_295), .Y(n_340) );
BUFx12f_ASAP7_75t_SL g341 ( .A(n_304), .Y(n_341) );
AOI21xp33_ASAP7_75t_L g342 ( .A1(n_312), .A2(n_230), .B(n_299), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_319), .A2(n_277), .B1(n_276), .B2(n_243), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_301), .A2(n_243), .B1(n_273), .B2(n_144), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_291), .A2(n_258), .B1(n_259), .B2(n_251), .Y(n_345) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_294), .A2(n_243), .B1(n_287), .B2(n_242), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_324), .Y(n_347) );
INVx4_ASAP7_75t_SL g348 ( .A(n_309), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_298), .B(n_247), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_322), .A2(n_243), .B1(n_254), .B2(n_248), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_309), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_304), .Y(n_352) );
AO32x2_ASAP7_75t_L g353 ( .A1(n_289), .A2(n_284), .A3(n_255), .B1(n_261), .B2(n_269), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_329), .B(n_228), .Y(n_354) );
AOI211xp5_ASAP7_75t_L g355 ( .A1(n_330), .A2(n_279), .B(n_284), .C(n_269), .Y(n_355) );
OAI222xp33_ASAP7_75t_L g356 ( .A1(n_294), .A2(n_252), .B1(n_239), .B2(n_262), .C1(n_242), .C2(n_269), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_290), .A2(n_268), .B1(n_269), .B2(n_265), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_292), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_314), .A2(n_265), .B1(n_255), .B2(n_280), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_322), .A2(n_234), .B1(n_288), .B2(n_280), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_329), .Y(n_362) );
INVx4_ASAP7_75t_SL g363 ( .A(n_309), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_313), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_302), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_305), .Y(n_366) );
BUFx12f_ASAP7_75t_L g367 ( .A(n_304), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_289), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_349), .B(n_317), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_340), .B(n_317), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_358), .B(n_292), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_355), .A2(n_308), .B1(n_307), .B2(n_305), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_340), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_366), .A2(n_327), .B(n_306), .Y(n_374) );
A2O1A1Ixp33_ASAP7_75t_L g375 ( .A1(n_342), .A2(n_310), .B(n_304), .C(n_311), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_338), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_348), .B(n_363), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_343), .A2(n_328), .B1(n_308), .B2(n_311), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_338), .B(n_300), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_366), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_345), .B(n_326), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_339), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_357), .A2(n_311), .B1(n_326), .B2(n_306), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g384 ( .A1(n_356), .A2(n_332), .B(n_336), .C(n_337), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_344), .B(n_333), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_367), .A2(n_311), .B1(n_325), .B2(n_320), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_339), .Y(n_387) );
OR2x6_ASAP7_75t_L g388 ( .A(n_367), .B(n_325), .Y(n_388) );
AOI21x1_ASAP7_75t_L g389 ( .A1(n_360), .A2(n_327), .B(n_252), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_352), .A2(n_234), .B1(n_323), .B2(n_318), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_347), .A2(n_337), .B1(n_239), .B2(n_262), .C(n_323), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_364), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_360), .A2(n_325), .B1(n_296), .B2(n_331), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_365), .A2(n_296), .B1(n_297), .B2(n_331), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_365), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_369), .B(n_364), .Y(n_396) );
OA21x2_ASAP7_75t_L g397 ( .A1(n_374), .A2(n_353), .B(n_318), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_382), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_373), .B(n_352), .Y(n_399) );
NAND4xp25_ASAP7_75t_L g400 ( .A(n_378), .B(n_350), .C(n_361), .D(n_359), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
AOI33xp33_ASAP7_75t_L g402 ( .A1(n_383), .A2(n_346), .A3(n_12), .B1(n_13), .B2(n_14), .B3(n_16), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_376), .A2(n_362), .B(n_368), .C(n_351), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_381), .A2(n_341), .B1(n_354), .B2(n_362), .Y(n_404) );
OAI211xp5_ASAP7_75t_SL g405 ( .A1(n_379), .A2(n_368), .B(n_222), .C(n_216), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_370), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g407 ( .A1(n_372), .A2(n_354), .B1(n_368), .B2(n_351), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_371), .A2(n_267), .B1(n_274), .B2(n_354), .C(n_249), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_382), .Y(n_409) );
OAI221xp5_ASAP7_75t_SL g410 ( .A1(n_375), .A2(n_341), .B1(n_274), .B2(n_267), .C(n_320), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_391), .B(n_150), .C(n_202), .Y(n_411) );
OAI211xp5_ASAP7_75t_SL g412 ( .A1(n_385), .A2(n_195), .B(n_194), .C(n_181), .Y(n_412) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_372), .B(n_10), .C(n_12), .D(n_13), .Y(n_413) );
OAI21x1_ASAP7_75t_L g414 ( .A1(n_374), .A2(n_335), .B(n_334), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_392), .A2(n_289), .B1(n_303), .B2(n_316), .Y(n_415) );
AOI221xp5_ASAP7_75t_SL g416 ( .A1(n_384), .A2(n_331), .B1(n_297), .B2(n_315), .C(n_296), .Y(n_416) );
OA21x2_ASAP7_75t_L g417 ( .A1(n_389), .A2(n_353), .B(n_297), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_393), .A2(n_293), .B(n_315), .Y(n_418) );
AND3x2_ASAP7_75t_L g419 ( .A(n_377), .B(n_363), .C(n_348), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_370), .A2(n_245), .B1(n_249), .B2(n_272), .C(n_315), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_393), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_388), .A2(n_320), .B1(n_289), .B2(n_303), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_387), .Y(n_423) );
OAI21xp33_ASAP7_75t_L g424 ( .A1(n_373), .A2(n_150), .B(n_229), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_388), .A2(n_303), .B1(n_316), .B2(n_241), .Y(n_425) );
NAND3xp33_ASAP7_75t_L g426 ( .A(n_394), .B(n_150), .C(n_167), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_388), .A2(n_303), .B1(n_316), .B2(n_241), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_387), .B(n_334), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_380), .B(n_348), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g430 ( .A1(n_394), .A2(n_272), .B(n_245), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_398), .B(n_380), .Y(n_431) );
INVx4_ASAP7_75t_L g432 ( .A(n_419), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_407), .A2(n_386), .B1(n_388), .B2(n_390), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_398), .B(n_395), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_409), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_406), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_421), .A2(n_388), .B1(n_395), .B2(n_377), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_423), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_397), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_402), .B(n_377), .Y(n_440) );
AND2x4_ASAP7_75t_L g441 ( .A(n_429), .B(n_377), .Y(n_441) );
AOI33xp33_ASAP7_75t_L g442 ( .A1(n_404), .A2(n_10), .A3(n_14), .B1(n_18), .B2(n_19), .B3(n_194), .Y(n_442) );
AOI33xp33_ASAP7_75t_L g443 ( .A1(n_415), .A2(n_19), .A3(n_195), .B1(n_197), .B2(n_168), .B3(n_169), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_401), .B(n_389), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_397), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_397), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_429), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_417), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_396), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_413), .A2(n_400), .B1(n_421), .B2(n_408), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_410), .A2(n_316), .B1(n_293), .B2(n_335), .Y(n_451) );
OAI33xp33_ASAP7_75t_L g452 ( .A1(n_399), .A2(n_195), .A3(n_168), .B1(n_169), .B2(n_172), .B3(n_222), .Y(n_452) );
INVx6_ASAP7_75t_L g453 ( .A(n_428), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_422), .A2(n_293), .B1(n_335), .B2(n_334), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_417), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_399), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_405), .A2(n_335), .B1(n_334), .B2(n_348), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_403), .A2(n_293), .B1(n_353), .B2(n_363), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_428), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_402), .Y(n_460) );
BUFx3_ASAP7_75t_L g461 ( .A(n_414), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_417), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_414), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_426), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_430), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_411), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_420), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_418), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_425), .B(n_293), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_416), .B(n_363), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_427), .B(n_293), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_424), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_412), .B(n_321), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_401), .B(n_226), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_398), .B(n_353), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_419), .Y(n_476) );
AOI222xp33_ASAP7_75t_L g477 ( .A1(n_396), .A2(n_321), .B1(n_150), .B2(n_234), .C1(n_232), .C2(n_226), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_419), .B(n_321), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_398), .B(n_353), .Y(n_479) );
NAND3xp33_ASAP7_75t_L g480 ( .A(n_460), .B(n_150), .C(n_167), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_435), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_436), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_442), .B(n_167), .C(n_202), .Y(n_483) );
OAI322xp33_ASAP7_75t_L g484 ( .A1(n_440), .A2(n_177), .A3(n_172), .B1(n_169), .B2(n_168), .C1(n_179), .C2(n_181), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_462), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_450), .A2(n_321), .B1(n_256), .B2(n_250), .Y(n_486) );
INVx2_ASAP7_75t_SL g487 ( .A(n_476), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_456), .B(n_232), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_475), .B(n_20), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_438), .Y(n_490) );
NOR3xp33_ASAP7_75t_L g491 ( .A(n_443), .B(n_179), .C(n_172), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_475), .B(n_21), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_479), .B(n_22), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_462), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_438), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_479), .B(n_24), .Y(n_496) );
NAND4xp25_ASAP7_75t_L g497 ( .A(n_449), .B(n_194), .C(n_177), .D(n_179), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_434), .B(n_321), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_448), .Y(n_499) );
INVx5_ASAP7_75t_L g500 ( .A(n_432), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_473), .A2(n_452), .B(n_464), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_434), .B(n_229), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_476), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_444), .B(n_28), .Y(n_504) );
AOI211xp5_ASAP7_75t_L g505 ( .A1(n_433), .A2(n_181), .B(n_177), .C(n_197), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_431), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_459), .B(n_37), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_431), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_448), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_444), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_447), .B(n_39), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_453), .B(n_40), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_467), .B(n_42), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_453), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_453), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_455), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_474), .B(n_45), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_432), .B(n_46), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_474), .B(n_49), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_439), .B(n_50), .Y(n_520) );
OAI221xp5_ASAP7_75t_SL g521 ( .A1(n_467), .A2(n_288), .B1(n_280), .B2(n_271), .C(n_235), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_437), .A2(n_237), .B1(n_241), .B2(n_256), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_439), .B(n_52), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_445), .B(n_53), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_455), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_445), .B(n_57), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_446), .Y(n_527) );
OAI211xp5_ASAP7_75t_L g528 ( .A1(n_432), .A2(n_458), .B(n_477), .C(n_470), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_446), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_441), .B(n_60), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_468), .Y(n_531) );
NAND4xp75_ASAP7_75t_SL g532 ( .A(n_478), .B(n_67), .C(n_73), .D(n_76), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_441), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_441), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_478), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_508), .B(n_465), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_482), .B(n_465), .Y(n_537) );
OAI31xp33_ASAP7_75t_L g538 ( .A1(n_528), .A2(n_478), .A3(n_466), .B(n_451), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_506), .B(n_468), .Y(n_539) );
INVx1_ASAP7_75t_SL g540 ( .A(n_503), .Y(n_540) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_485), .Y(n_541) );
INVx2_ASAP7_75t_SL g542 ( .A(n_487), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_481), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_490), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_495), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_510), .B(n_464), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_533), .B(n_469), .Y(n_547) );
AND4x1_ASAP7_75t_L g548 ( .A(n_505), .B(n_457), .C(n_471), .D(n_472), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_527), .Y(n_549) );
OAI31xp33_ASAP7_75t_L g550 ( .A1(n_521), .A2(n_454), .A3(n_461), .B(n_469), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_534), .B(n_461), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_525), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_487), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_529), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_511), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_529), .Y(n_556) );
AND2x4_ASAP7_75t_SL g557 ( .A(n_518), .B(n_463), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_514), .B(n_216), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_499), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_499), .Y(n_560) );
NOR2x1_ASAP7_75t_L g561 ( .A(n_497), .B(n_205), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_515), .B(n_208), .Y(n_562) );
OAI21xp5_ASAP7_75t_SL g563 ( .A1(n_518), .A2(n_235), .B(n_280), .Y(n_563) );
NOR2xp33_ASAP7_75t_SL g564 ( .A(n_500), .B(n_256), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_509), .B(n_216), .Y(n_565) );
NAND4xp25_ASAP7_75t_L g566 ( .A(n_513), .B(n_222), .C(n_208), .D(n_197), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_509), .B(n_208), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_516), .B(n_205), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_535), .B(n_241), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_500), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_513), .B(n_167), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_531), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_494), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_500), .B(n_275), .Y(n_574) );
NAND3xp33_ASAP7_75t_SL g575 ( .A(n_511), .B(n_275), .C(n_241), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_504), .B(n_237), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_504), .B(n_202), .Y(n_577) );
OAI21xp33_ASAP7_75t_L g578 ( .A1(n_486), .A2(n_202), .B(n_167), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_535), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_494), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_489), .B(n_237), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_542), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_570), .B(n_500), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_543), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_536), .B(n_546), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_554), .B(n_492), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_553), .A2(n_501), .B1(n_483), .B2(n_492), .C(n_496), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_554), .B(n_493), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_573), .B(n_493), .Y(n_589) );
NOR4xp25_ASAP7_75t_L g590 ( .A(n_540), .B(n_507), .C(n_496), .D(n_489), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_544), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_570), .Y(n_592) );
OAI322xp33_ASAP7_75t_L g593 ( .A1(n_555), .A2(n_488), .A3(n_502), .B1(n_530), .B2(n_519), .C1(n_517), .C2(n_498), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_545), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_563), .A2(n_518), .B1(n_500), .B2(n_524), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g596 ( .A1(n_575), .A2(n_480), .B(n_522), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_552), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_539), .B(n_524), .Y(n_598) );
INVx2_ASAP7_75t_SL g599 ( .A(n_573), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_579), .B(n_523), .Y(n_600) );
INVxp33_ASAP7_75t_L g601 ( .A(n_574), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_538), .B(n_526), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_549), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_557), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_561), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_557), .Y(n_606) );
AOI222xp33_ASAP7_75t_L g607 ( .A1(n_537), .A2(n_520), .B1(n_526), .B2(n_512), .C1(n_532), .C2(n_488), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_572), .B(n_491), .Y(n_608) );
NAND2x1_ASAP7_75t_L g609 ( .A(n_556), .B(n_484), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_541), .B(n_167), .Y(n_610) );
NOR2xp67_ASAP7_75t_L g611 ( .A(n_575), .B(n_202), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_560), .Y(n_612) );
OAI211xp5_ASAP7_75t_L g613 ( .A1(n_550), .A2(n_202), .B(n_288), .C(n_271), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_559), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_559), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_SL g616 ( .A1(n_574), .A2(n_288), .B(n_235), .C(n_271), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_541), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_547), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_580), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_576), .A2(n_250), .B1(n_256), .B2(n_271), .Y(n_620) );
AND2x4_ASAP7_75t_L g621 ( .A(n_551), .B(n_250), .Y(n_621) );
XNOR2x2_ASAP7_75t_L g622 ( .A(n_566), .B(n_256), .Y(n_622) );
XOR2xp5_ASAP7_75t_L g623 ( .A(n_569), .B(n_235), .Y(n_623) );
OAI221xp5_ASAP7_75t_L g624 ( .A1(n_548), .A2(n_285), .B1(n_213), .B2(n_225), .C(n_275), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_565), .Y(n_625) );
AO22x2_ASAP7_75t_L g626 ( .A1(n_581), .A2(n_213), .B1(n_225), .B2(n_285), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_567), .B(n_213), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_571), .A2(n_166), .B1(n_225), .B2(n_562), .C(n_577), .Y(n_628) );
OA21x2_ASAP7_75t_L g629 ( .A1(n_568), .A2(n_225), .B(n_166), .Y(n_629) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_571), .B(n_166), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_558), .B(n_166), .Y(n_631) );
NAND2xp33_ASAP7_75t_R g632 ( .A(n_564), .B(n_166), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_578), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_542), .B(n_166), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_590), .B(n_618), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g636 ( .A1(n_602), .A2(n_613), .B(n_595), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_L g637 ( .A1(n_602), .A2(n_601), .B(n_582), .C(n_592), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_606), .A2(n_604), .B1(n_592), .B2(n_601), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_583), .A2(n_630), .B1(n_605), .B2(n_611), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_594), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_634), .Y(n_641) );
AOI222xp33_ASAP7_75t_L g642 ( .A1(n_587), .A2(n_584), .B1(n_608), .B2(n_586), .C1(n_588), .C2(n_597), .Y(n_642) );
INVx1_ASAP7_75t_SL g643 ( .A(n_585), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_583), .A2(n_616), .B(n_609), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_591), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_599), .A2(n_626), .B(n_596), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_599), .B(n_603), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_640), .Y(n_648) );
XNOR2x1_ASAP7_75t_L g649 ( .A(n_638), .B(n_622), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_645), .Y(n_650) );
AOI211xp5_ASAP7_75t_SL g651 ( .A1(n_646), .A2(n_593), .B(n_624), .C(n_633), .Y(n_651) );
AOI211xp5_ASAP7_75t_SL g652 ( .A1(n_636), .A2(n_628), .B(n_620), .C(n_625), .Y(n_652) );
AOI21xp33_ASAP7_75t_L g653 ( .A1(n_635), .A2(n_607), .B(n_626), .Y(n_653) );
AO22x2_ASAP7_75t_L g654 ( .A1(n_643), .A2(n_617), .B1(n_612), .B2(n_619), .Y(n_654) );
OAI31xp33_ASAP7_75t_L g655 ( .A1(n_637), .A2(n_623), .A3(n_588), .B(n_586), .Y(n_655) );
OAI22xp5_ASAP7_75t_SL g656 ( .A1(n_649), .A2(n_641), .B1(n_639), .B2(n_644), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_654), .A2(n_647), .B1(n_642), .B2(n_589), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_652), .B(n_647), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_651), .B(n_632), .C(n_631), .D(n_621), .Y(n_659) );
OR3x1_ASAP7_75t_L g660 ( .A(n_659), .B(n_653), .C(n_655), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_656), .A2(n_654), .B1(n_650), .B2(n_648), .Y(n_661) );
OR4x2_ASAP7_75t_L g662 ( .A(n_657), .B(n_655), .C(n_600), .D(n_589), .Y(n_662) );
BUFx2_ASAP7_75t_SL g663 ( .A(n_661), .Y(n_663) );
NOR2x1p5_ASAP7_75t_L g664 ( .A(n_660), .B(n_658), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_664), .B(n_615), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_663), .Y(n_666) );
AOI222xp33_ASAP7_75t_SL g667 ( .A1(n_666), .A2(n_662), .B1(n_620), .B2(n_614), .C1(n_629), .C2(n_621), .Y(n_667) );
OAI22xp33_ASAP7_75t_L g668 ( .A1(n_667), .A2(n_665), .B1(n_627), .B2(n_598), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g669 ( .A1(n_668), .A2(n_610), .B1(n_629), .B2(n_627), .Y(n_669) );
endmodule