module fake_jpeg_6025_n_251 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx10_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_19),
.B1(n_30),
.B2(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_21),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_47),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_50),
.B1(n_40),
.B2(n_20),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_33),
.B(n_35),
.C(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_53),
.Y(n_71)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_59),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_19),
.B1(n_24),
.B2(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_21),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_20),
.Y(n_74)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_31),
.C(n_22),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_62),
.B1(n_25),
.B2(n_23),
.Y(n_80)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_19),
.B1(n_15),
.B2(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_69),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_76),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_74),
.B(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_44),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_26),
.Y(n_106)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_79),
.Y(n_95)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_17),
.B1(n_22),
.B2(n_64),
.Y(n_104)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_100),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_52),
.B(n_60),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_98),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_67),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_16),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_51),
.B(n_16),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_23),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_98),
.B1(n_85),
.B2(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_17),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_114),
.Y(n_147)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_80),
.B1(n_43),
.B2(n_57),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_122),
.B1(n_78),
.B2(n_65),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_127),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_104),
.B1(n_93),
.B2(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_86),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_99),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_85),
.A2(n_57),
.B1(n_43),
.B2(n_73),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_77),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_124),
.B(n_128),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_92),
.A2(n_73),
.B1(n_68),
.B2(n_79),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_136),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_90),
.B(n_92),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_139),
.B1(n_140),
.B2(n_143),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_27),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_94),
.C(n_106),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_142),
.C(n_27),
.Y(n_157)
);

AOI32xp33_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_94),
.A3(n_68),
.B1(n_101),
.B2(n_105),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_125),
.C(n_110),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_65),
.B1(n_54),
.B2(n_39),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_26),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_34),
.C(n_96),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_111),
.B1(n_113),
.B2(n_116),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_39),
.B1(n_28),
.B2(n_84),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_144),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_111),
.B(n_96),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_34),
.B(n_96),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_88),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_34),
.B1(n_28),
.B2(n_72),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_108),
.A2(n_28),
.B1(n_87),
.B2(n_88),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_152),
.B(n_167),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_129),
.B(n_109),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_156),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_141),
.C(n_136),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_143),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_163),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_168),
.Y(n_185)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_114),
.Y(n_165)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_166),
.B(n_112),
.Y(n_173)
);

NOR4xp25_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_88),
.C(n_1),
.D(n_2),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_27),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_171),
.A2(n_160),
.B1(n_155),
.B2(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_132),
.B(n_130),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_183),
.B(n_154),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_190),
.Y(n_196)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_87),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_139),
.C(n_140),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_187),
.Y(n_197)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_131),
.C(n_138),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_146),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_135),
.B1(n_150),
.B2(n_112),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_189),
.A2(n_170),
.B1(n_169),
.B2(n_135),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_181),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_182),
.C(n_26),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_156),
.C(n_168),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_200),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_161),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_183),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_154),
.B1(n_87),
.B2(n_27),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_204),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_178),
.A2(n_0),
.B(n_3),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_188),
.B(n_180),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_213),
.B(n_215),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_196),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_174),
.C(n_184),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_211),
.C(n_205),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_198),
.C(n_201),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_196),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_212),
.B(n_219),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_182),
.B(n_4),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_218),
.C(n_216),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_223),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_204),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_225),
.B(n_228),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_200),
.C(n_26),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_227),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_4),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_5),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_5),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_222),
.A2(n_214),
.B1(n_6),
.B2(n_8),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_233),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_234),
.Y(n_241)
);

NOR2x1_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_8),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_237),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_242),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g242 ( 
.A(n_235),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_236),
.A3(n_232),
.B1(n_234),
.B2(n_231),
.C1(n_226),
.C2(n_8),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_9),
.C(n_10),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.C1(n_14),
.C2(n_235),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_244),
.C(n_246),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_248),
.C(n_11),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_9),
.C(n_13),
.Y(n_251)
);


endmodule