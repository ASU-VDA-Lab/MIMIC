module real_jpeg_14052_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_307, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_307;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_300;
wire n_221;
wire n_292;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_293;
wire n_164;
wire n_275;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_285;
wire n_45;
wire n_160;
wire n_304;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_295;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g109 ( 
.A(n_0),
.Y(n_109)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_2),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_2),
.A2(n_29),
.B1(n_47),
.B2(n_48),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_2),
.A2(n_29),
.B1(n_41),
.B2(n_45),
.Y(n_234)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_4),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_4),
.A2(n_41),
.B1(n_45),
.B2(n_114),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_114),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_4),
.A2(n_26),
.B1(n_28),
.B2(n_114),
.Y(n_208)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_7),
.A2(n_26),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_34),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_7),
.A2(n_34),
.B1(n_41),
.B2(n_45),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_7),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_10),
.A2(n_41),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_53),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_10),
.A2(n_26),
.B1(n_28),
.B2(n_53),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_10),
.B(n_59),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_10),
.B(n_44),
.C(n_48),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_10),
.B(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_10),
.B(n_46),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_10),
.A2(n_24),
.B(n_61),
.C(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_10),
.B(n_20),
.Y(n_187)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_93),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_91),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_83),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_15),
.B(n_83),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_69),
.C(n_75),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_16),
.A2(n_17),
.B1(n_69),
.B2(n_77),
.Y(n_301)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_35),
.B1(n_36),
.B2(n_68),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_18),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_25),
.B(n_30),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_19),
.A2(n_73),
.B(n_74),
.Y(n_278)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_20),
.B(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_20),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_20),
.B(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_22),
.B1(n_26),
.B2(n_28),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_21),
.B(n_24),
.C(n_53),
.Y(n_199)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_23),
.A2(n_24),
.B1(n_61),
.B2(n_62),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_25),
.A2(n_70),
.B(n_73),
.Y(n_88)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_26),
.B(n_199),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_30),
.B(n_207),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_31),
.B(n_208),
.Y(n_218)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_54),
.B1(n_55),
.B2(n_67),
.Y(n_36)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_37),
.B(n_77),
.C(n_78),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_37),
.B(n_55),
.C(n_68),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_37),
.A2(n_67),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_37),
.A2(n_67),
.B1(n_78),
.B2(n_295),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_51),
.B(n_52),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_38),
.A2(n_118),
.B(n_234),
.Y(n_264)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_39),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_39),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_39),
.B(n_119),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_45),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_41),
.B(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AO22x1_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_45),
.A2(n_53),
.B(n_62),
.Y(n_170)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_46),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_46),
.B(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_46),
.B(n_133),
.Y(n_177)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_48),
.B(n_109),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_48),
.B(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_51),
.A2(n_165),
.B(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_52),
.Y(n_133)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_63),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_57),
.B(n_220),
.Y(n_219)
);

NAND2x1_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_59),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_58),
.B(n_86),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_59),
.B(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_59),
.A2(n_63),
.B(n_80),
.Y(n_282)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_66),
.Y(n_82)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_63),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_79),
.B(n_81),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_64),
.B(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_67),
.B(n_205),
.C(n_211),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_69),
.A2(n_77),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_70),
.B(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_72),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_74),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_75),
.A2(n_76),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_78),
.Y(n_295)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_82),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_82),
.B(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_90),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_85),
.A2(n_89),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_85),
.B(n_224),
.C(n_230),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_285),
.B(n_302),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_268),
.B(n_284),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_247),
.B(n_267),
.Y(n_96)
);

AOI321xp33_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_214),
.A3(n_240),
.B1(n_245),
.B2(n_246),
.C(n_307),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_190),
.B(n_213),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_173),
.B(n_189),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_156),
.B(n_172),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_134),
.B(n_155),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_126),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_126),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_115),
.B1(n_116),
.B2(n_125),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_110),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_105),
.B(n_152),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_112),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_107),
.A2(n_109),
.B(n_112),
.Y(n_168)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_109),
.A2(n_152),
.B(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_145),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_112),
.A2(n_201),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_118),
.B(n_132),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_120),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_123),
.C(n_125),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_128),
.B1(n_130),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_148),
.B(n_154),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_142),
.B(n_147),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_144),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_146),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_158),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_166),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_164),
.C(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_163),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_165),
.B(n_177),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_171),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_167),
.A2(n_168),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_167),
.A2(n_168),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_169),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_168),
.B(n_264),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_168),
.A2(n_275),
.B(n_277),
.Y(n_289)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_188),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_188),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_181),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_179),
.C(n_181),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_186),
.C(n_187),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_192),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_203),
.B2(n_204),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_196),
.C(n_203),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_202),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_209),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_235),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_235),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_222),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_223),
.C(n_231),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.C(n_221),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_219),
.CI(n_221),
.CON(n_237),
.SN(n_237)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_231),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_227),
.Y(n_238)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_233),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.C(n_239),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_237),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_237),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_244),
.Y(n_245)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_249),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_266),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_262),
.B2(n_263),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_263),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_255),
.C(n_260),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_264),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_270),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_273),
.C(n_280),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_279),
.B2(n_280),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B(n_283),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_282),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_283),
.A2(n_291),
.B1(n_292),
.B2(n_296),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_283),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_289),
.C(n_291),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_297),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_288),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_299),
.Y(n_304)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);


endmodule