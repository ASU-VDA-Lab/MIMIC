module fake_ariane_3061_n_5378 (n_913, n_589, n_1174, n_691, n_423, n_603, n_373, n_1250, n_1169, n_789, n_850, n_610, n_245, n_96, n_319, n_49, n_690, n_416, n_1109, n_525, n_187, n_1238, n_817, n_924, n_781, n_189, n_717, n_72, n_952, n_864, n_1096, n_57, n_117, n_524, n_1214, n_634, n_1246, n_1138, n_214, n_764, n_462, n_1196, n_1181, n_32, n_410, n_1187, n_1131, n_1225, n_737, n_137, n_232, n_52, n_568, n_1088, n_77, n_766, n_377, n_520, n_870, n_279, n_945, n_958, n_813, n_419, n_146, n_270, n_338, n_995, n_285, n_1184, n_202, n_500, n_665, n_754, n_903, n_871, n_1073, n_239, n_402, n_54, n_829, n_1062, n_339, n_738, n_672, n_740, n_167, n_1018, n_69, n_259, n_953, n_143, n_1224, n_625, n_557, n_1107, n_989, n_242, n_645, n_331, n_559, n_267, n_495, n_350, n_381, n_795, n_721, n_1084, n_200, n_1241, n_821, n_561, n_770, n_507, n_486, n_901, n_569, n_1145, n_971, n_787, n_31, n_1195, n_518, n_1207, n_222, n_786, n_868, n_884, n_1034, n_1085, n_277, n_432, n_293, n_823, n_620, n_93, n_1074, n_859, n_108, n_587, n_693, n_863, n_303, n_1254, n_929, n_206, n_352, n_899, n_611, n_238, n_365, n_1013, n_136, n_334, n_192, n_661, n_300, n_533, n_104, n_438, n_16, n_440, n_273, n_1230, n_612, n_333, n_376, n_512, n_579, n_844, n_1012, n_149, n_1213, n_237, n_780, n_1021, n_491, n_1142, n_1140, n_705, n_570, n_260, n_942, n_7, n_461, n_1121, n_209, n_490, n_17, n_225, n_1006, n_575, n_546, n_503, n_1112, n_700, n_1159, n_772, n_1216, n_1245, n_676, n_42, n_680, n_287, n_302, n_380, n_94, n_4, n_249, n_1108, n_355, n_212, n_65, n_123, n_444, n_851, n_257, n_652, n_475, n_135, n_947, n_930, n_1260, n_1179, n_468, n_102, n_182, n_696, n_482, n_798, n_577, n_407, n_27, n_916, n_912, n_460, n_366, n_762, n_1253, n_555, n_804, n_966, n_992, n_955, n_1182, n_794, n_78, n_514, n_418, n_513, n_288, n_179, n_1178, n_1026, n_306, n_92, n_203, n_436, n_150, n_324, n_669, n_931, n_619, n_337, n_437, n_111, n_21, n_274, n_967, n_1083, n_746, n_292, n_1079, n_615, n_1139, n_76, n_517, n_0, n_824, n_428, n_159, n_892, n_959, n_30, n_1101, n_563, n_144, n_990, n_867, n_1226, n_944, n_749, n_815, n_542, n_470, n_1240, n_1087, n_632, n_477, n_650, n_425, n_1155, n_1071, n_712, n_976, n_909, n_767, n_964, n_382, n_489, n_80, n_251, n_974, n_506, n_799, n_1147, n_397, n_471, n_351, n_965, n_155, n_934, n_1220, n_356, n_698, n_124, n_307, n_1209, n_1020, n_646, n_34, n_404, n_172, n_1058, n_347, n_1042, n_183, n_1234, n_479, n_299, n_836, n_564, n_133, n_66, n_205, n_1029, n_1247, n_760, n_522, n_20, n_367, n_1111, n_970, n_713, n_1255, n_598, n_345, n_1237, n_927, n_261, n_1095, n_370, n_706, n_286, n_776, n_424, n_85, n_130, n_466, n_1263, n_346, n_348, n_552, n_670, n_379, n_138, n_162, n_264, n_441, n_1032, n_1217, n_637, n_73, n_327, n_1259, n_1177, n_1231, n_980, n_905, n_207, n_720, n_926, n_41, n_194, n_1163, n_186, n_145, n_59, n_1173, n_1068, n_1198, n_487, n_90, n_855, n_158, n_808, n_553, n_814, n_578, n_405, n_120, n_320, n_1134, n_647, n_481, n_600, n_1053, n_529, n_502, n_218, n_247, n_1105, n_547, n_439, n_604, n_677, n_478, n_703, n_1061, n_326, n_681, n_227, n_874, n_707, n_11, n_129, n_126, n_983, n_590, n_699, n_727, n_301, n_545, n_1015, n_1162, n_536, n_325, n_688, n_636, n_427, n_1098, n_442, n_777, n_1080, n_920, n_1086, n_1092, n_986, n_1104, n_729, n_887, n_1122, n_1205, n_163, n_1132, n_390, n_1156, n_501, n_314, n_1120, n_1202, n_627, n_1188, n_233, n_957, n_388, n_1242, n_1218, n_221, n_321, n_86, n_861, n_877, n_1119, n_616, n_1055, n_1189, n_1089, n_281, n_262, n_735, n_297, n_1005, n_527, n_46, n_84, n_845, n_888, n_178, n_551, n_417, n_70, n_343, n_1222, n_582, n_755, n_1097, n_1219, n_710, n_534, n_1239, n_278, n_560, n_890, n_842, n_148, n_451, n_745, n_61, n_742, n_1081, n_1266, n_769, n_13, n_476, n_832, n_55, n_535, n_744, n_982, n_915, n_215, n_1075, n_454, n_298, n_1227, n_655, n_403, n_1007, n_657, n_837, n_812, n_606, n_951, n_862, n_659, n_509, n_666, n_430, n_1206, n_722, n_1171, n_1030, n_785, n_999, n_456, n_852, n_704, n_1060, n_1044, n_521, n_873, n_1243, n_342, n_358, n_608, n_1037, n_317, n_134, n_1257, n_1078, n_266, n_157, n_1161, n_811, n_624, n_791, n_876, n_618, n_1191, n_736, n_1025, n_1215, n_241, n_687, n_797, n_480, n_211, n_642, n_97, n_408, n_595, n_602, n_592, n_854, n_393, n_474, n_805, n_295, n_190, n_1072, n_695, n_64, n_180, n_730, n_386, n_516, n_1137, n_1258, n_197, n_640, n_463, n_943, n_1118, n_678, n_651, n_961, n_469, n_1046, n_726, n_1123, n_878, n_771, n_752, n_71, n_985, n_421, n_906, n_1180, n_283, n_806, n_649, n_374, n_643, n_226, n_682, n_36, n_819, n_586, n_686, n_605, n_1154, n_584, n_1130, n_349, n_756, n_1016, n_1149, n_979, n_2, n_897, n_949, n_515, n_807, n_891, n_885, n_198, n_1208, n_396, n_802, n_23, n_1151, n_554, n_960, n_1256, n_87, n_714, n_790, n_354, n_140, n_725, n_151, n_28, n_1009, n_230, n_1133, n_154, n_883, n_142, n_473, n_801, n_818, n_779, n_594, n_35, n_1052, n_272, n_833, n_879, n_1117, n_38, n_422, n_597, n_75, n_1047, n_95, n_1050, n_566, n_152, n_169, n_106, n_1201, n_173, n_858, n_1185, n_335, n_1035, n_1143, n_344, n_426, n_433, n_398, n_62, n_210, n_1090, n_166, n_253, n_928, n_1153, n_271, n_465, n_825, n_1103, n_732, n_1192, n_128, n_224, n_82, n_894, n_420, n_562, n_748, n_510, n_1045, n_256, n_1160, n_1023, n_988, n_330, n_914, n_400, n_689, n_1116, n_282, n_328, n_368, n_467, n_644, n_1197, n_276, n_497, n_1165, n_168, n_81, n_538, n_576, n_843, n_511, n_455, n_429, n_588, n_638, n_1128, n_1048, n_775, n_667, n_1049, n_14, n_869, n_141, n_846, n_305, n_312, n_56, n_60, n_728, n_413, n_715, n_889, n_1066, n_935, n_685, n_911, n_361, n_89, n_623, n_1065, n_453, n_74, n_810, n_19, n_40, n_181, n_617, n_543, n_236, n_601, n_683, n_565, n_628, n_743, n_1194, n_907, n_660, n_464, n_962, n_941, n_1210, n_847, n_747, n_1135, n_918, n_107, n_639, n_452, n_673, n_1038, n_414, n_571, n_6, n_284, n_593, n_1164, n_37, n_58, n_609, n_1193, n_613, n_1022, n_1033, n_409, n_171, n_519, n_384, n_1166, n_1056, n_526, n_1040, n_674, n_1158, n_316, n_125, n_820, n_43, n_872, n_254, n_1157, n_234, n_848, n_280, n_629, n_161, n_532, n_763, n_99, n_540, n_216, n_692, n_5, n_984, n_223, n_750, n_834, n_800, n_395, n_621, n_213, n_67, n_1014, n_724, n_493, n_114, n_1100, n_585, n_875, n_827, n_697, n_622, n_296, n_880, n_793, n_1175, n_132, n_751, n_1027, n_1070, n_739, n_1028, n_1221, n_530, n_792, n_1262, n_580, n_494, n_434, n_975, n_229, n_394, n_923, n_1124, n_932, n_1183, n_981, n_1110, n_243, n_185, n_1204, n_994, n_973, n_268, n_972, n_164, n_184, n_856, n_1248, n_1176, n_1054, n_508, n_118, n_121, n_353, n_1057, n_191, n_978, n_1011, n_828, n_322, n_558, n_116, n_39, n_653, n_783, n_556, n_1127, n_170, n_160, n_119, n_1008, n_332, n_581, n_294, n_1024, n_830, n_176, n_987, n_936, n_541, n_499, n_788, n_12, n_908, n_1036, n_341, n_109, n_1167, n_549, n_591, n_969, n_919, n_50, n_318, n_103, n_244, n_679, n_220, n_663, n_443, n_528, n_1200, n_387, n_406, n_826, n_139, n_391, n_940, n_1077, n_607, n_956, n_445, n_765, n_122, n_385, n_917, n_372, n_15, n_631, n_399, n_1170, n_1261, n_702, n_857, n_898, n_363, n_968, n_1067, n_1235, n_1064, n_633, n_900, n_1093, n_193, n_733, n_761, n_731, n_336, n_315, n_311, n_8, n_668, n_758, n_1106, n_47, n_153, n_18, n_648, n_784, n_269, n_816, n_835, n_446, n_1076, n_753, n_701, n_1003, n_1125, n_309, n_115, n_401, n_485, n_504, n_483, n_435, n_1141, n_291, n_822, n_1094, n_840, n_1099, n_839, n_79, n_3, n_759, n_567, n_91, n_240, n_369, n_44, n_1172, n_614, n_1212, n_831, n_778, n_48, n_188, n_323, n_550, n_997, n_635, n_694, n_1113, n_248, n_1152, n_921, n_1236, n_228, n_1265, n_671, n_1, n_1148, n_654, n_488, n_904, n_505, n_88, n_498, n_1059, n_684, n_1039, n_539, n_1150, n_977, n_449, n_392, n_459, n_1136, n_458, n_1190, n_1144, n_383, n_838, n_175, n_950, n_1017, n_711, n_734, n_723, n_658, n_630, n_53, n_362, n_310, n_709, n_24, n_809, n_235, n_881, n_1019, n_662, n_641, n_910, n_290, n_741, n_939, n_371, n_199, n_217, n_1114, n_708, n_308, n_1223, n_201, n_572, n_1199, n_865, n_10, n_1041, n_993, n_948, n_922, n_1004, n_448, n_860, n_1043, n_255, n_450, n_896, n_902, n_1031, n_853, n_716, n_196, n_774, n_933, n_596, n_954, n_1168, n_219, n_231, n_656, n_492, n_574, n_252, n_664, n_1229, n_68, n_415, n_63, n_544, n_1186, n_599, n_768, n_1091, n_537, n_1063, n_25, n_991, n_83, n_389, n_1126, n_195, n_938, n_895, n_110, n_304, n_583, n_1000, n_313, n_626, n_378, n_98, n_946, n_757, n_375, n_113, n_33, n_1146, n_1203, n_998, n_472, n_937, n_265, n_208, n_156, n_174, n_275, n_100, n_147, n_204, n_1232, n_996, n_1211, n_963, n_1264, n_51, n_1082, n_496, n_866, n_26, n_246, n_925, n_1001, n_1115, n_1002, n_105, n_1051, n_719, n_131, n_263, n_1102, n_360, n_1129, n_1252, n_250, n_773, n_165, n_1010, n_882, n_1249, n_101, n_803, n_329, n_718, n_340, n_289, n_9, n_112, n_45, n_548, n_523, n_457, n_177, n_782, n_364, n_258, n_431, n_1228, n_1244, n_411, n_484, n_849, n_22, n_29, n_357, n_412, n_1251, n_447, n_1233, n_893, n_841, n_886, n_1069, n_359, n_573, n_796, n_127, n_531, n_675, n_5378);

input n_913;
input n_589;
input n_1174;
input n_691;
input n_423;
input n_603;
input n_373;
input n_1250;
input n_1169;
input n_789;
input n_850;
input n_610;
input n_245;
input n_96;
input n_319;
input n_49;
input n_690;
input n_416;
input n_1109;
input n_525;
input n_187;
input n_1238;
input n_817;
input n_924;
input n_781;
input n_189;
input n_717;
input n_72;
input n_952;
input n_864;
input n_1096;
input n_57;
input n_117;
input n_524;
input n_1214;
input n_634;
input n_1246;
input n_1138;
input n_214;
input n_764;
input n_462;
input n_1196;
input n_1181;
input n_32;
input n_410;
input n_1187;
input n_1131;
input n_1225;
input n_737;
input n_137;
input n_232;
input n_52;
input n_568;
input n_1088;
input n_77;
input n_766;
input n_377;
input n_520;
input n_870;
input n_279;
input n_945;
input n_958;
input n_813;
input n_419;
input n_146;
input n_270;
input n_338;
input n_995;
input n_285;
input n_1184;
input n_202;
input n_500;
input n_665;
input n_754;
input n_903;
input n_871;
input n_1073;
input n_239;
input n_402;
input n_54;
input n_829;
input n_1062;
input n_339;
input n_738;
input n_672;
input n_740;
input n_167;
input n_1018;
input n_69;
input n_259;
input n_953;
input n_143;
input n_1224;
input n_625;
input n_557;
input n_1107;
input n_989;
input n_242;
input n_645;
input n_331;
input n_559;
input n_267;
input n_495;
input n_350;
input n_381;
input n_795;
input n_721;
input n_1084;
input n_200;
input n_1241;
input n_821;
input n_561;
input n_770;
input n_507;
input n_486;
input n_901;
input n_569;
input n_1145;
input n_971;
input n_787;
input n_31;
input n_1195;
input n_518;
input n_1207;
input n_222;
input n_786;
input n_868;
input n_884;
input n_1034;
input n_1085;
input n_277;
input n_432;
input n_293;
input n_823;
input n_620;
input n_93;
input n_1074;
input n_859;
input n_108;
input n_587;
input n_693;
input n_863;
input n_303;
input n_1254;
input n_929;
input n_206;
input n_352;
input n_899;
input n_611;
input n_238;
input n_365;
input n_1013;
input n_136;
input n_334;
input n_192;
input n_661;
input n_300;
input n_533;
input n_104;
input n_438;
input n_16;
input n_440;
input n_273;
input n_1230;
input n_612;
input n_333;
input n_376;
input n_512;
input n_579;
input n_844;
input n_1012;
input n_149;
input n_1213;
input n_237;
input n_780;
input n_1021;
input n_491;
input n_1142;
input n_1140;
input n_705;
input n_570;
input n_260;
input n_942;
input n_7;
input n_461;
input n_1121;
input n_209;
input n_490;
input n_17;
input n_225;
input n_1006;
input n_575;
input n_546;
input n_503;
input n_1112;
input n_700;
input n_1159;
input n_772;
input n_1216;
input n_1245;
input n_676;
input n_42;
input n_680;
input n_287;
input n_302;
input n_380;
input n_94;
input n_4;
input n_249;
input n_1108;
input n_355;
input n_212;
input n_65;
input n_123;
input n_444;
input n_851;
input n_257;
input n_652;
input n_475;
input n_135;
input n_947;
input n_930;
input n_1260;
input n_1179;
input n_468;
input n_102;
input n_182;
input n_696;
input n_482;
input n_798;
input n_577;
input n_407;
input n_27;
input n_916;
input n_912;
input n_460;
input n_366;
input n_762;
input n_1253;
input n_555;
input n_804;
input n_966;
input n_992;
input n_955;
input n_1182;
input n_794;
input n_78;
input n_514;
input n_418;
input n_513;
input n_288;
input n_179;
input n_1178;
input n_1026;
input n_306;
input n_92;
input n_203;
input n_436;
input n_150;
input n_324;
input n_669;
input n_931;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_967;
input n_1083;
input n_746;
input n_292;
input n_1079;
input n_615;
input n_1139;
input n_76;
input n_517;
input n_0;
input n_824;
input n_428;
input n_159;
input n_892;
input n_959;
input n_30;
input n_1101;
input n_563;
input n_144;
input n_990;
input n_867;
input n_1226;
input n_944;
input n_749;
input n_815;
input n_542;
input n_470;
input n_1240;
input n_1087;
input n_632;
input n_477;
input n_650;
input n_425;
input n_1155;
input n_1071;
input n_712;
input n_976;
input n_909;
input n_767;
input n_964;
input n_382;
input n_489;
input n_80;
input n_251;
input n_974;
input n_506;
input n_799;
input n_1147;
input n_397;
input n_471;
input n_351;
input n_965;
input n_155;
input n_934;
input n_1220;
input n_356;
input n_698;
input n_124;
input n_307;
input n_1209;
input n_1020;
input n_646;
input n_34;
input n_404;
input n_172;
input n_1058;
input n_347;
input n_1042;
input n_183;
input n_1234;
input n_479;
input n_299;
input n_836;
input n_564;
input n_133;
input n_66;
input n_205;
input n_1029;
input n_1247;
input n_760;
input n_522;
input n_20;
input n_367;
input n_1111;
input n_970;
input n_713;
input n_1255;
input n_598;
input n_345;
input n_1237;
input n_927;
input n_261;
input n_1095;
input n_370;
input n_706;
input n_286;
input n_776;
input n_424;
input n_85;
input n_130;
input n_466;
input n_1263;
input n_346;
input n_348;
input n_552;
input n_670;
input n_379;
input n_138;
input n_162;
input n_264;
input n_441;
input n_1032;
input n_1217;
input n_637;
input n_73;
input n_327;
input n_1259;
input n_1177;
input n_1231;
input n_980;
input n_905;
input n_207;
input n_720;
input n_926;
input n_41;
input n_194;
input n_1163;
input n_186;
input n_145;
input n_59;
input n_1173;
input n_1068;
input n_1198;
input n_487;
input n_90;
input n_855;
input n_158;
input n_808;
input n_553;
input n_814;
input n_578;
input n_405;
input n_120;
input n_320;
input n_1134;
input n_647;
input n_481;
input n_600;
input n_1053;
input n_529;
input n_502;
input n_218;
input n_247;
input n_1105;
input n_547;
input n_439;
input n_604;
input n_677;
input n_478;
input n_703;
input n_1061;
input n_326;
input n_681;
input n_227;
input n_874;
input n_707;
input n_11;
input n_129;
input n_126;
input n_983;
input n_590;
input n_699;
input n_727;
input n_301;
input n_545;
input n_1015;
input n_1162;
input n_536;
input n_325;
input n_688;
input n_636;
input n_427;
input n_1098;
input n_442;
input n_777;
input n_1080;
input n_920;
input n_1086;
input n_1092;
input n_986;
input n_1104;
input n_729;
input n_887;
input n_1122;
input n_1205;
input n_163;
input n_1132;
input n_390;
input n_1156;
input n_501;
input n_314;
input n_1120;
input n_1202;
input n_627;
input n_1188;
input n_233;
input n_957;
input n_388;
input n_1242;
input n_1218;
input n_221;
input n_321;
input n_86;
input n_861;
input n_877;
input n_1119;
input n_616;
input n_1055;
input n_1189;
input n_1089;
input n_281;
input n_262;
input n_735;
input n_297;
input n_1005;
input n_527;
input n_46;
input n_84;
input n_845;
input n_888;
input n_178;
input n_551;
input n_417;
input n_70;
input n_343;
input n_1222;
input n_582;
input n_755;
input n_1097;
input n_1219;
input n_710;
input n_534;
input n_1239;
input n_278;
input n_560;
input n_890;
input n_842;
input n_148;
input n_451;
input n_745;
input n_61;
input n_742;
input n_1081;
input n_1266;
input n_769;
input n_13;
input n_476;
input n_832;
input n_55;
input n_535;
input n_744;
input n_982;
input n_915;
input n_215;
input n_1075;
input n_454;
input n_298;
input n_1227;
input n_655;
input n_403;
input n_1007;
input n_657;
input n_837;
input n_812;
input n_606;
input n_951;
input n_862;
input n_659;
input n_509;
input n_666;
input n_430;
input n_1206;
input n_722;
input n_1171;
input n_1030;
input n_785;
input n_999;
input n_456;
input n_852;
input n_704;
input n_1060;
input n_1044;
input n_521;
input n_873;
input n_1243;
input n_342;
input n_358;
input n_608;
input n_1037;
input n_317;
input n_134;
input n_1257;
input n_1078;
input n_266;
input n_157;
input n_1161;
input n_811;
input n_624;
input n_791;
input n_876;
input n_618;
input n_1191;
input n_736;
input n_1025;
input n_1215;
input n_241;
input n_687;
input n_797;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_602;
input n_592;
input n_854;
input n_393;
input n_474;
input n_805;
input n_295;
input n_190;
input n_1072;
input n_695;
input n_64;
input n_180;
input n_730;
input n_386;
input n_516;
input n_1137;
input n_1258;
input n_197;
input n_640;
input n_463;
input n_943;
input n_1118;
input n_678;
input n_651;
input n_961;
input n_469;
input n_1046;
input n_726;
input n_1123;
input n_878;
input n_771;
input n_752;
input n_71;
input n_985;
input n_421;
input n_906;
input n_1180;
input n_283;
input n_806;
input n_649;
input n_374;
input n_643;
input n_226;
input n_682;
input n_36;
input n_819;
input n_586;
input n_686;
input n_605;
input n_1154;
input n_584;
input n_1130;
input n_349;
input n_756;
input n_1016;
input n_1149;
input n_979;
input n_2;
input n_897;
input n_949;
input n_515;
input n_807;
input n_891;
input n_885;
input n_198;
input n_1208;
input n_396;
input n_802;
input n_23;
input n_1151;
input n_554;
input n_960;
input n_1256;
input n_87;
input n_714;
input n_790;
input n_354;
input n_140;
input n_725;
input n_151;
input n_28;
input n_1009;
input n_230;
input n_1133;
input n_154;
input n_883;
input n_142;
input n_473;
input n_801;
input n_818;
input n_779;
input n_594;
input n_35;
input n_1052;
input n_272;
input n_833;
input n_879;
input n_1117;
input n_38;
input n_422;
input n_597;
input n_75;
input n_1047;
input n_95;
input n_1050;
input n_566;
input n_152;
input n_169;
input n_106;
input n_1201;
input n_173;
input n_858;
input n_1185;
input n_335;
input n_1035;
input n_1143;
input n_344;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_1090;
input n_166;
input n_253;
input n_928;
input n_1153;
input n_271;
input n_465;
input n_825;
input n_1103;
input n_732;
input n_1192;
input n_128;
input n_224;
input n_82;
input n_894;
input n_420;
input n_562;
input n_748;
input n_510;
input n_1045;
input n_256;
input n_1160;
input n_1023;
input n_988;
input n_330;
input n_914;
input n_400;
input n_689;
input n_1116;
input n_282;
input n_328;
input n_368;
input n_467;
input n_644;
input n_1197;
input n_276;
input n_497;
input n_1165;
input n_168;
input n_81;
input n_538;
input n_576;
input n_843;
input n_511;
input n_455;
input n_429;
input n_588;
input n_638;
input n_1128;
input n_1048;
input n_775;
input n_667;
input n_1049;
input n_14;
input n_869;
input n_141;
input n_846;
input n_305;
input n_312;
input n_56;
input n_60;
input n_728;
input n_413;
input n_715;
input n_889;
input n_1066;
input n_935;
input n_685;
input n_911;
input n_361;
input n_89;
input n_623;
input n_1065;
input n_453;
input n_74;
input n_810;
input n_19;
input n_40;
input n_181;
input n_617;
input n_543;
input n_236;
input n_601;
input n_683;
input n_565;
input n_628;
input n_743;
input n_1194;
input n_907;
input n_660;
input n_464;
input n_962;
input n_941;
input n_1210;
input n_847;
input n_747;
input n_1135;
input n_918;
input n_107;
input n_639;
input n_452;
input n_673;
input n_1038;
input n_414;
input n_571;
input n_6;
input n_284;
input n_593;
input n_1164;
input n_37;
input n_58;
input n_609;
input n_1193;
input n_613;
input n_1022;
input n_1033;
input n_409;
input n_171;
input n_519;
input n_384;
input n_1166;
input n_1056;
input n_526;
input n_1040;
input n_674;
input n_1158;
input n_316;
input n_125;
input n_820;
input n_43;
input n_872;
input n_254;
input n_1157;
input n_234;
input n_848;
input n_280;
input n_629;
input n_161;
input n_532;
input n_763;
input n_99;
input n_540;
input n_216;
input n_692;
input n_5;
input n_984;
input n_223;
input n_750;
input n_834;
input n_800;
input n_395;
input n_621;
input n_213;
input n_67;
input n_1014;
input n_724;
input n_493;
input n_114;
input n_1100;
input n_585;
input n_875;
input n_827;
input n_697;
input n_622;
input n_296;
input n_880;
input n_793;
input n_1175;
input n_132;
input n_751;
input n_1027;
input n_1070;
input n_739;
input n_1028;
input n_1221;
input n_530;
input n_792;
input n_1262;
input n_580;
input n_494;
input n_434;
input n_975;
input n_229;
input n_394;
input n_923;
input n_1124;
input n_932;
input n_1183;
input n_981;
input n_1110;
input n_243;
input n_185;
input n_1204;
input n_994;
input n_973;
input n_268;
input n_972;
input n_164;
input n_184;
input n_856;
input n_1248;
input n_1176;
input n_1054;
input n_508;
input n_118;
input n_121;
input n_353;
input n_1057;
input n_191;
input n_978;
input n_1011;
input n_828;
input n_322;
input n_558;
input n_116;
input n_39;
input n_653;
input n_783;
input n_556;
input n_1127;
input n_170;
input n_160;
input n_119;
input n_1008;
input n_332;
input n_581;
input n_294;
input n_1024;
input n_830;
input n_176;
input n_987;
input n_936;
input n_541;
input n_499;
input n_788;
input n_12;
input n_908;
input n_1036;
input n_341;
input n_109;
input n_1167;
input n_549;
input n_591;
input n_969;
input n_919;
input n_50;
input n_318;
input n_103;
input n_244;
input n_679;
input n_220;
input n_663;
input n_443;
input n_528;
input n_1200;
input n_387;
input n_406;
input n_826;
input n_139;
input n_391;
input n_940;
input n_1077;
input n_607;
input n_956;
input n_445;
input n_765;
input n_122;
input n_385;
input n_917;
input n_372;
input n_15;
input n_631;
input n_399;
input n_1170;
input n_1261;
input n_702;
input n_857;
input n_898;
input n_363;
input n_968;
input n_1067;
input n_1235;
input n_1064;
input n_633;
input n_900;
input n_1093;
input n_193;
input n_733;
input n_761;
input n_731;
input n_336;
input n_315;
input n_311;
input n_8;
input n_668;
input n_758;
input n_1106;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_816;
input n_835;
input n_446;
input n_1076;
input n_753;
input n_701;
input n_1003;
input n_1125;
input n_309;
input n_115;
input n_401;
input n_485;
input n_504;
input n_483;
input n_435;
input n_1141;
input n_291;
input n_822;
input n_1094;
input n_840;
input n_1099;
input n_839;
input n_79;
input n_3;
input n_759;
input n_567;
input n_91;
input n_240;
input n_369;
input n_44;
input n_1172;
input n_614;
input n_1212;
input n_831;
input n_778;
input n_48;
input n_188;
input n_323;
input n_550;
input n_997;
input n_635;
input n_694;
input n_1113;
input n_248;
input n_1152;
input n_921;
input n_1236;
input n_228;
input n_1265;
input n_671;
input n_1;
input n_1148;
input n_654;
input n_488;
input n_904;
input n_505;
input n_88;
input n_498;
input n_1059;
input n_684;
input n_1039;
input n_539;
input n_1150;
input n_977;
input n_449;
input n_392;
input n_459;
input n_1136;
input n_458;
input n_1190;
input n_1144;
input n_383;
input n_838;
input n_175;
input n_950;
input n_1017;
input n_711;
input n_734;
input n_723;
input n_658;
input n_630;
input n_53;
input n_362;
input n_310;
input n_709;
input n_24;
input n_809;
input n_235;
input n_881;
input n_1019;
input n_662;
input n_641;
input n_910;
input n_290;
input n_741;
input n_939;
input n_371;
input n_199;
input n_217;
input n_1114;
input n_708;
input n_308;
input n_1223;
input n_201;
input n_572;
input n_1199;
input n_865;
input n_10;
input n_1041;
input n_993;
input n_948;
input n_922;
input n_1004;
input n_448;
input n_860;
input n_1043;
input n_255;
input n_450;
input n_896;
input n_902;
input n_1031;
input n_853;
input n_716;
input n_196;
input n_774;
input n_933;
input n_596;
input n_954;
input n_1168;
input n_219;
input n_231;
input n_656;
input n_492;
input n_574;
input n_252;
input n_664;
input n_1229;
input n_68;
input n_415;
input n_63;
input n_544;
input n_1186;
input n_599;
input n_768;
input n_1091;
input n_537;
input n_1063;
input n_25;
input n_991;
input n_83;
input n_389;
input n_1126;
input n_195;
input n_938;
input n_895;
input n_110;
input n_304;
input n_583;
input n_1000;
input n_313;
input n_626;
input n_378;
input n_98;
input n_946;
input n_757;
input n_375;
input n_113;
input n_33;
input n_1146;
input n_1203;
input n_998;
input n_472;
input n_937;
input n_265;
input n_208;
input n_156;
input n_174;
input n_275;
input n_100;
input n_147;
input n_204;
input n_1232;
input n_996;
input n_1211;
input n_963;
input n_1264;
input n_51;
input n_1082;
input n_496;
input n_866;
input n_26;
input n_246;
input n_925;
input n_1001;
input n_1115;
input n_1002;
input n_105;
input n_1051;
input n_719;
input n_131;
input n_263;
input n_1102;
input n_360;
input n_1129;
input n_1252;
input n_250;
input n_773;
input n_165;
input n_1010;
input n_882;
input n_1249;
input n_101;
input n_803;
input n_329;
input n_718;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_548;
input n_523;
input n_457;
input n_177;
input n_782;
input n_364;
input n_258;
input n_431;
input n_1228;
input n_1244;
input n_411;
input n_484;
input n_849;
input n_22;
input n_29;
input n_357;
input n_412;
input n_1251;
input n_447;
input n_1233;
input n_893;
input n_841;
input n_886;
input n_1069;
input n_359;
input n_573;
input n_796;
input n_127;
input n_531;
input n_675;

output n_5378;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_2182;
wire n_2680;
wire n_3264;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_2729;
wire n_4302;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_5302;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_2646;
wire n_2653;
wire n_4610;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_2482;
wire n_1682;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_4260;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_2322;
wire n_2663;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_4143;
wire n_4273;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_4567;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_3015;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_3482;
wire n_1900;
wire n_4268;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_5247;
wire n_4476;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_2382;
wire n_5292;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_3458;
wire n_3511;
wire n_2077;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_3549;
wire n_3914;
wire n_1692;
wire n_2611;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5056;
wire n_2015;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_2257;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5179;
wire n_2435;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_3814;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_2019;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2649;
wire n_1568;
wire n_2919;
wire n_3108;
wire n_2632;
wire n_4314;
wire n_2980;
wire n_1728;
wire n_4315;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_2697;
wire n_1817;
wire n_3704;
wire n_4296;
wire n_2677;
wire n_2483;
wire n_5088;
wire n_1592;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_5149;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_5089;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_5296;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1349;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_4292;
wire n_2118;
wire n_1490;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_3025;
wire n_3051;
wire n_2802;
wire n_2125;
wire n_4974;
wire n_5123;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1498;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_2707;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_3713;
wire n_1863;
wire n_4798;
wire n_1500;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_3944;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_2448;
wire n_2211;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_2958;
wire n_1714;
wire n_4429;
wire n_3340;
wire n_5053;
wire n_3486;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_2520;
wire n_3864;
wire n_4694;
wire n_4664;
wire n_3450;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_1406;
wire n_5073;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_2991;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_4822;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_3740;
wire n_2417;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_3726;
wire n_4419;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_3421;
wire n_1448;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_4966;
wire n_2250;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_2610;
wire n_1593;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_3886;
wire n_2619;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_2613;
wire n_1517;
wire n_2647;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_1671;
wire n_5027;
wire n_2343;
wire n_3380;
wire n_2826;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_4631;
wire n_1504;
wire n_2110;
wire n_5377;
wire n_3822;
wire n_4355;
wire n_3818;
wire n_3587;
wire n_2608;
wire n_1948;
wire n_4155;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_4685;
wire n_3927;
wire n_2068;
wire n_3595;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_3396;
wire n_4093;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_2963;
wire n_2561;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_5125;
wire n_4922;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_3630;
wire n_1612;
wire n_1910;
wire n_2189;
wire n_4194;
wire n_2672;
wire n_2018;
wire n_2602;
wire n_2931;
wire n_3433;
wire n_3597;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_3786;
wire n_2828;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_3645;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_5011;
wire n_1554;
wire n_3279;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_1679;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_4053;
wire n_3963;
wire n_3091;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_1775;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_3225;
wire n_3621;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_3633;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_2009;
wire n_4339;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_3457;
wire n_2324;
wire n_5283;
wire n_3454;
wire n_2139;
wire n_2521;
wire n_2740;
wire n_1991;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_5040;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_3628;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_3872;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_3555;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_4574;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_4663;
wire n_3296;
wire n_3794;
wire n_3762;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_3707;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_5304;
wire n_1581;
wire n_3058;
wire n_2047;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_5355;
wire n_3592;
wire n_5321;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_1368;
wire n_4120;
wire n_2880;
wire n_1313;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_1339;
wire n_5116;
wire n_3771;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_2830;
wire n_4622;
wire n_4757;
wire n_1871;
wire n_4016;
wire n_3334;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_4591;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_2259;
wire n_5337;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_4493;
wire n_1808;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_3181;
wire n_1916;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_1566;
wire n_2837;
wire n_2446;
wire n_4116;
wire n_5360;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_4439;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_2248;
wire n_4660;
wire n_3081;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_2844;
wire n_1979;
wire n_4814;
wire n_2221;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_2634;
wire n_2746;
wire n_5098;
wire n_1276;
wire n_5145;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_1528;
wire n_3315;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_5213;
wire n_3474;
wire n_2458;
wire n_3150;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1652;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_2685;
wire n_2061;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_4995;
wire n_4498;
wire n_2743;
wire n_2969;
wire n_3429;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_4850;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_3391;
wire n_4786;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_3240;
wire n_5066;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_5130;
wire n_4175;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_2172;
wire n_2601;
wire n_2365;
wire n_1880;
wire n_1399;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_3257;
wire n_3730;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_4003;
wire n_1832;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5159;
wire n_4022;
wire n_2495;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_1279;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_3031;
wire n_2335;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_5287;
wire n_4719;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_2296;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_2059;
wire n_4713;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_4916;
wire n_4323;
wire n_1899;
wire n_5376;
wire n_3508;
wire n_4129;
wire n_3599;
wire n_4480;
wire n_3734;
wire n_3401;
wire n_3542;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_2218;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_3995;
wire n_3908;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_2266;
wire n_4324;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_3671;
wire n_2366;
wire n_1753;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_3791;
wire n_2008;
wire n_4989;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_1332;
wire n_1747;
wire n_3990;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5256;
wire n_4779;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_1400;
wire n_3735;
wire n_1513;
wire n_1527;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1954;
wire n_3964;
wire n_5364;
wire n_3302;
wire n_2486;
wire n_1897;
wire n_2137;
wire n_3685;
wire n_4977;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_2912;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_2264;
wire n_1950;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_3411;
wire n_5222;
wire n_3463;
wire n_2785;
wire n_4938;
wire n_2574;
wire n_1281;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1697;
wire n_2730;
wire n_5129;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_1561;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5161;
wire n_1557;
wire n_4744;
wire n_4706;
wire n_2022;
wire n_3879;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_4990;
wire n_2986;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_3317;
wire n_4835;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_4372;
wire n_4097;
wire n_4162;
wire n_5293;
wire n_4790;
wire n_4173;
wire n_5309;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_3973;
wire n_4799;
wire n_4534;
wire n_4960;
wire n_3738;
wire n_1380;
wire n_2020;
wire n_2310;
wire n_3600;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_3967;
wire n_4370;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_2234;
wire n_1341;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_2592;
wire n_3490;
wire n_5043;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_1968;
wire n_5020;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_4333;
wire n_5339;
wire n_2007;
wire n_3363;
wire n_1803;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_3481;
wire n_5101;
wire n_2236;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_2406;
wire n_4477;
wire n_4110;
wire n_5182;
wire n_4217;
wire n_5277;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_3873;
wire n_4649;
wire n_2428;
wire n_1360;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_4999;
wire n_4592;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_2385;
wire n_1980;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_3114;
wire n_2092;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_2402;
wire n_1458;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_1550;
wire n_1358;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_3687;
wire n_2787;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_5193;
wire n_4933;
wire n_4144;
wire n_2375;
wire n_3278;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_4726;
wire n_5143;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_5273;
wire n_2469;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_3068;
wire n_1629;
wire n_1510;
wire n_3002;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_3132;
wire n_5002;
wire n_3681;
wire n_3970;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_4579;
wire n_4776;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_4165;
wire n_2056;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1941;
wire n_3637;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_1686;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_2297;
wire n_1410;
wire n_4203;
wire n_1325;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_3674;
wire n_1638;
wire n_1571;
wire n_5349;
wire n_3763;
wire n_3499;
wire n_1821;
wire n_3947;
wire n_3910;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_3088;
wire n_1724;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_5375;
wire n_4958;
wire n_1827;
wire n_4149;
wire n_2361;
wire n_1752;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_3075;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_2304;
wire n_2514;
wire n_1299;
wire n_3430;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_4971;
wire n_2095;
wire n_2738;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_2423;
wire n_2208;
wire n_1421;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_2866;
wire n_3153;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_1383;
wire n_4259;
wire n_2030;
wire n_4299;
wire n_2407;
wire n_5367;
wire n_2243;
wire n_5288;
wire n_2694;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_5294;
wire n_2731;
wire n_3703;
wire n_5265;
wire n_2123;
wire n_2238;
wire n_4802;
wire n_4793;
wire n_3435;
wire n_2380;
wire n_4897;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_3220;
wire n_4581;
wire n_4625;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_5316;
wire n_2735;
wire n_4214;
wire n_1888;
wire n_5290;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_4032;
wire n_2571;
wire n_4929;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_3634;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_4815;
wire n_4665;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_1461;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_4174;
wire n_5131;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_3119;
wire n_4740;
wire n_1274;
wire n_4394;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_2628;
wire n_1491;
wire n_3219;
wire n_5333;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_3479;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_2755;
wire n_5109;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_2220;
wire n_4433;
wire n_2829;
wire n_1914;
wire n_2253;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_3936;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_2473;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_3078;
wire n_3971;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_4751;
wire n_4242;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_4952;
wire n_4426;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_2112;
wire n_2640;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_4506;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_4039;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_3983;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_2338;
wire n_5261;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_2594;
wire n_5298;
wire n_3417;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_4328;
wire n_1854;
wire n_5191;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_4940;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_2280;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_3586;
wire n_4160;
wire n_1668;
wire n_4137;
wire n_4545;
wire n_4758;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_4535;
wire n_4385;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_4766;
wire n_4558;
wire n_1318;
wire n_1769;
wire n_1632;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1733;
wire n_4651;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_1352;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1822;
wire n_1441;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_2907;
wire n_2353;
wire n_1429;
wire n_2528;
wire n_1778;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_3718;
wire n_3390;
wire n_2298;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_3976;
wire n_2813;
wire n_2546;
wire n_3381;
wire n_3736;
wire n_4466;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_5369;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_4377;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5270;
wire n_3468;
wire n_1877;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_2497;
wire n_4561;
wire n_3291;
wire n_1541;
wire n_1472;
wire n_2578;
wire n_2475;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5351;
wire n_5267;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_3358;
wire n_2533;
wire n_2003;
wire n_1307;
wire n_4682;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_1440;
wire n_1370;
wire n_5005;
wire n_1549;
wire n_5207;
wire n_2658;
wire n_3620;
wire n_4601;
wire n_4518;
wire n_2767;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_2862;
wire n_4325;
wire n_2553;
wire n_1420;
wire n_2645;
wire n_4711;
wire n_2749;
wire n_4413;
wire n_3307;
wire n_3251;
wire n_1885;
wire n_3288;
wire n_2833;
wire n_3723;
wire n_4135;
wire n_5223;
wire n_3880;
wire n_3904;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_3532;
wire n_5154;
wire n_2609;
wire n_1767;
wire n_3131;
wire n_4138;
wire n_1973;
wire n_1444;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_4270;
wire n_4620;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_1645;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_2465;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_1834;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_4858;
wire n_1445;
wire n_5370;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_1663;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_3897;
wire n_1735;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_1271;
wire n_2186;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_1285;
wire n_3838;
wire n_4059;
wire n_5194;
wire n_2734;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_3273;
wire n_2918;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3001;
wire n_5260;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_5372;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_2422;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_1393;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_3032;
wire n_4886;
wire n_5172;
wire n_1477;
wire n_1982;
wire n_5311;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1273;
wire n_2982;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_4693;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_4487;
wire n_2674;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_3112;
wire n_2562;
wire n_1779;
wire n_2051;
wire n_3196;
wire n_2673;
wire n_4678;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_1891;
wire n_5348;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_1725;
wire n_2318;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_3045;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_4047;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_2135;
wire n_4475;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_2461;
wire n_1706;
wire n_3719;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_1503;
wire n_5295;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_3383;
wire n_1835;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_2323;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_1988;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_2078;
wire n_4809;
wire n_4012;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_5042;
wire n_4768;
wire n_1889;
wire n_5368;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_2727;
wire n_5234;
wire n_1416;
wire n_1599;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_5253;
wire n_3588;
wire n_3280;
wire n_1590;
wire n_4115;
wire n_5274;
wire n_5019;
wire n_1819;
wire n_3095;
wire n_3698;
wire n_4513;
wire n_1442;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2549;
wire n_2499;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_4264;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_4170;
wire n_2462;
wire n_2155;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_4267;
wire n_2083;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_2378;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_1483;
wire n_1363;
wire n_3467;
wire n_3179;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_3699;
wire n_2120;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_5335;
wire n_2801;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_3246;
wire n_3299;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_3276;
wire n_3682;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_2932;
wire n_2027;
wire n_3118;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_1467;
wire n_5209;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_5099;
wire n_3286;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_3009;
wire n_5219;
wire n_3951;
wire n_3035;
wire n_4261;
wire n_1823;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_1666;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_3224;
wire n_1969;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_1572;
wire n_4463;
wire n_5357;
wire n_3648;
wire n_1975;
wire n_1388;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_1532;
wire n_5181;
wire n_3208;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_2916;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_3650;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_5017;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_2091;
wire n_4312;
wire n_3789;
wire n_1658;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_4537;
wire n_3694;
wire n_3893;
wire n_4847;
wire n_2307;
wire n_3702;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_1971;
wire n_2945;
wire n_3543;
wire n_1324;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_2698;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_5142;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_4595;
wire n_2352;
wire n_5201;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_4054;
wire n_1286;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_4732;
wire n_2203;
wire n_2076;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_4139;
wire n_4769;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_3509;
wire n_1403;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_3790;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_2174;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_5228;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_4720;
wire n_2889;
wire n_2141;
wire n_1758;
wire n_3470;
wire n_5221;
wire n_1407;
wire n_2865;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_3677;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_4131;
wire n_4215;
wire n_2488;
wire n_1509;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_2169;
wire n_5133;
wire n_5305;
wire n_2175;
wire n_1625;
wire n_4578;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_2724;
wire n_2258;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_5343;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_2268;
wire n_3469;
wire n_2835;
wire n_1452;
wire n_2111;
wire n_3743;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_4472;
wire n_2699;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_2710;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_4371;
wire n_1902;
wire n_2784;
wire n_3898;
wire n_4749;
wire n_1845;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_3094;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_5034;
wire n_3312;
wire n_2451;
wire n_2913;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_1764;
wire n_4807;
wire n_5115;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_4095;
wire n_1310;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1699;
wire n_5226;
wire n_2081;
wire n_1474;
wire n_1631;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_4516;
wire n_5235;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_1870;
wire n_4467;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_5258;

INVx1_ASAP7_75t_L g1267 ( 
.A(n_984),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1174),
.Y(n_1268)
);

BUFx10_ASAP7_75t_L g1269 ( 
.A(n_1068),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1163),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_818),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_216),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_973),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1218),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_604),
.Y(n_1275)
);

INVxp67_ASAP7_75t_L g1276 ( 
.A(n_1194),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1073),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_881),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_871),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1247),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1157),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_860),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_523),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_702),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1127),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_15),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_658),
.Y(n_1287)
);

BUFx5_ASAP7_75t_L g1288 ( 
.A(n_191),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1232),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_533),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_130),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_39),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1076),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1254),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_538),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_726),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_966),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_781),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_270),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_363),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1042),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_887),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_563),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_340),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_1158),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1132),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1003),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_913),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_773),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1167),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_672),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_352),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_396),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_731),
.Y(n_1314)
);

BUFx8_ASAP7_75t_SL g1315 ( 
.A(n_12),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1019),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_496),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1120),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1191),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_44),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_273),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1175),
.Y(n_1322)
);

CKINVDCx14_ASAP7_75t_R g1323 ( 
.A(n_923),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_1006),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_644),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_745),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_553),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_760),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_907),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_915),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1138),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1130),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1173),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1093),
.Y(n_1334)
);

BUFx10_ASAP7_75t_L g1335 ( 
.A(n_1134),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_125),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_106),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1236),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1094),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_675),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_968),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1066),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_692),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_588),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1233),
.Y(n_1345)
);

BUFx2_ASAP7_75t_SL g1346 ( 
.A(n_132),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1263),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1077),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_942),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_950),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_819),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_791),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1160),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_631),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1121),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_425),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_461),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1250),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_873),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_167),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1108),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1200),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_535),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_204),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1039),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_488),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_352),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1156),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_801),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_111),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_383),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_558),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_864),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_848),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_535),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_513),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_666),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_906),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_1096),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_86),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_936),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_661),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_391),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_891),
.Y(n_1384)
);

BUFx10_ASAP7_75t_L g1385 ( 
.A(n_454),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_537),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_459),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_971),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1177),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1141),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_496),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_8),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_630),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_207),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_171),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_325),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_304),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_582),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_223),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_805),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_615),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1085),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_943),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_910),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_389),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_236),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1128),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_328),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1083),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_306),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1171),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1165),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1170),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_356),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_642),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1240),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_507),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1208),
.Y(n_1418)
);

CKINVDCx14_ASAP7_75t_R g1419 ( 
.A(n_1017),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_534),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_239),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_951),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_920),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_606),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1059),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1102),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1179),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_220),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_335),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_837),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_879),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_114),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_656),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_878),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_359),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_857),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_544),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_637),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1169),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_159),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1026),
.Y(n_1441)
);

BUFx10_ASAP7_75t_L g1442 ( 
.A(n_890),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_412),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_945),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_932),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_500),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1072),
.Y(n_1447)
);

INVx4_ASAP7_75t_R g1448 ( 
.A(n_1205),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_30),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_427),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1075),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1148),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1154),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1152),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_665),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_806),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_321),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_911),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1235),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_32),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_956),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_536),
.Y(n_1462)
);

BUFx5_ASAP7_75t_L g1463 ( 
.A(n_1264),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_617),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1149),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_986),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_179),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_351),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1029),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_645),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1114),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1110),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_97),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_909),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_689),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1098),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1185),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_754),
.Y(n_1478)
);

BUFx10_ASAP7_75t_L g1479 ( 
.A(n_359),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1207),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_300),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_954),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_957),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_943),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1043),
.Y(n_1485)
);

BUFx10_ASAP7_75t_L g1486 ( 
.A(n_163),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_840),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1181),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_342),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_603),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1000),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1199),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_922),
.Y(n_1493)
);

CKINVDCx20_ASAP7_75t_R g1494 ( 
.A(n_952),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_885),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1078),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_127),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_562),
.Y(n_1498)
);

BUFx10_ASAP7_75t_L g1499 ( 
.A(n_675),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_241),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_532),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1224),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_938),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1221),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_1253),
.Y(n_1505)
);

CKINVDCx16_ASAP7_75t_R g1506 ( 
.A(n_41),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_930),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_238),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_965),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_169),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_934),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_341),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_995),
.Y(n_1513)
);

BUFx10_ASAP7_75t_L g1514 ( 
.A(n_1150),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1084),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_917),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_328),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_981),
.Y(n_1518)
);

INVxp33_ASAP7_75t_L g1519 ( 
.A(n_547),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_872),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_618),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1021),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_557),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1266),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_892),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_700),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1071),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_646),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_740),
.Y(n_1529)
);

BUFx10_ASAP7_75t_L g1530 ( 
.A(n_934),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_996),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_157),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_157),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_257),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_979),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1013),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_582),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_17),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_919),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_429),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_339),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_699),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_640),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_135),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_307),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_857),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1228),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_489),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_188),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1105),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_749),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_163),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_216),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1237),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1054),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_751),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_72),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_98),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_963),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1227),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_901),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_459),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_845),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_148),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_889),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1225),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1213),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_897),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_519),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_940),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1219),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_648),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_881),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_19),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_405),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1057),
.Y(n_1576)
);

BUFx10_ASAP7_75t_L g1577 ( 
.A(n_316),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_763),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1187),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_26),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_558),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_806),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_683),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_810),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_423),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_792),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_532),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_252),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_765),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1126),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_691),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_311),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_906),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_299),
.Y(n_1595)
);

CKINVDCx14_ASAP7_75t_R g1596 ( 
.A(n_1257),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_99),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1100),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_59),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_671),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_749),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_299),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_991),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_695),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1062),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_176),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1113),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1143),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1015),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1220),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1162),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_141),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1089),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1069),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_741),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_347),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_31),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1229),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1111),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_472),
.Y(n_1620)
);

BUFx5_ASAP7_75t_L g1621 ( 
.A(n_678),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1209),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_162),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_738),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_724),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1139),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_90),
.Y(n_1627)
);

CKINVDCx20_ASAP7_75t_R g1628 ( 
.A(n_1265),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_896),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1012),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1135),
.Y(n_1631)
);

BUFx10_ASAP7_75t_L g1632 ( 
.A(n_933),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_16),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_768),
.Y(n_1634)
);

CKINVDCx16_ASAP7_75t_R g1635 ( 
.A(n_961),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1193),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_660),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_187),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_182),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_1212),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1180),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1217),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_967),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_236),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_908),
.Y(n_1645)
);

BUFx5_ASAP7_75t_L g1646 ( 
.A(n_629),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1183),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_631),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1215),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_617),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1260),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_875),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_221),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_892),
.Y(n_1654)
);

BUFx10_ASAP7_75t_L g1655 ( 
.A(n_866),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_373),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_629),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_467),
.Y(n_1658)
);

CKINVDCx20_ASAP7_75t_R g1659 ( 
.A(n_384),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_937),
.Y(n_1660)
);

BUFx10_ASAP7_75t_L g1661 ( 
.A(n_667),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_66),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_135),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1238),
.Y(n_1664)
);

CKINVDCx16_ASAP7_75t_R g1665 ( 
.A(n_550),
.Y(n_1665)
);

CKINVDCx20_ASAP7_75t_R g1666 ( 
.A(n_314),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_706),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_953),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_570),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_725),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_478),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_444),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1206),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_944),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_306),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_605),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_252),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1092),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1222),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_560),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_340),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_627),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_240),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_226),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1234),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_949),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_824),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_11),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_440),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1124),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1258),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1245),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1202),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1107),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1184),
.Y(n_1695)
);

CKINVDCx20_ASAP7_75t_R g1696 ( 
.A(n_214),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_191),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_988),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_676),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_738),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_245),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1081),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_717),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1005),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1117),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_261),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1052),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1140),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_935),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_893),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_476),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1242),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_209),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_894),
.Y(n_1714)
);

BUFx10_ASAP7_75t_L g1715 ( 
.A(n_1091),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1131),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_212),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_205),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_315),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_482),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_413),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1151),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_844),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_307),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_903),
.Y(n_1725)
);

CKINVDCx14_ASAP7_75t_R g1726 ( 
.A(n_423),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_811),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1080),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_488),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_904),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_336),
.Y(n_1731)
);

CKINVDCx14_ASAP7_75t_R g1732 ( 
.A(n_829),
.Y(n_1732)
);

CKINVDCx20_ASAP7_75t_R g1733 ( 
.A(n_886),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_825),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_622),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_448),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1196),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1168),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_657),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_468),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_916),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1027),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_96),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_736),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_227),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1038),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1186),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1025),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1122),
.Y(n_1749)
);

CKINVDCx20_ASAP7_75t_R g1750 ( 
.A(n_743),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1203),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_888),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_874),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1262),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_217),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_898),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_347),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_1197),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_931),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1097),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1155),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_872),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_324),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1190),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_268),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_946),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_25),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_696),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_924),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_642),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_648),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_389),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_97),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_440),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_556),
.Y(n_1775)
);

CKINVDCx20_ASAP7_75t_R g1776 ( 
.A(n_1166),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_623),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_584),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1125),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_551),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_640),
.Y(n_1781)
);

BUFx5_ASAP7_75t_L g1782 ( 
.A(n_72),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_750),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1249),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1079),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_447),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_744),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1244),
.Y(n_1788)
);

CKINVDCx20_ASAP7_75t_R g1789 ( 
.A(n_927),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_457),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1159),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_10),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1189),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_800),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_859),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1256),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_150),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1090),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1095),
.Y(n_1799)
);

CKINVDCx20_ASAP7_75t_R g1800 ( 
.A(n_584),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1070),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_974),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_933),
.Y(n_1803)
);

INVx2_ASAP7_75t_SL g1804 ( 
.A(n_833),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1255),
.Y(n_1805)
);

BUFx10_ASAP7_75t_L g1806 ( 
.A(n_390),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_668),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_569),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_255),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_671),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_225),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_233),
.Y(n_1812)
);

CKINVDCx20_ASAP7_75t_R g1813 ( 
.A(n_166),
.Y(n_1813)
);

BUFx3_ASAP7_75t_L g1814 ( 
.A(n_926),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_784),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_137),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_156),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1261),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_89),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1176),
.Y(n_1820)
);

CKINVDCx20_ASAP7_75t_R g1821 ( 
.A(n_895),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_63),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_1161),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_653),
.Y(n_1824)
);

BUFx2_ASAP7_75t_L g1825 ( 
.A(n_544),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_52),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1211),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_305),
.Y(n_1828)
);

INVx1_ASAP7_75t_SL g1829 ( 
.A(n_348),
.Y(n_1829)
);

CKINVDCx20_ASAP7_75t_R g1830 ( 
.A(n_36),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1087),
.Y(n_1831)
);

BUFx3_ASAP7_75t_L g1832 ( 
.A(n_740),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_654),
.Y(n_1833)
);

INVx2_ASAP7_75t_SL g1834 ( 
.A(n_14),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_85),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_478),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_733),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_232),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_224),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_563),
.Y(n_1840)
);

BUFx2_ASAP7_75t_L g1841 ( 
.A(n_825),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_291),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_421),
.Y(n_1843)
);

INVxp67_ASAP7_75t_L g1844 ( 
.A(n_1182),
.Y(n_1844)
);

BUFx2_ASAP7_75t_L g1845 ( 
.A(n_1210),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1239),
.Y(n_1846)
);

CKINVDCx20_ASAP7_75t_R g1847 ( 
.A(n_371),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_366),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_905),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_2),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_65),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_1032),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_925),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_275),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1023),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1109),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_877),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_51),
.Y(n_1858)
);

BUFx6f_ASAP7_75t_L g1859 ( 
.A(n_588),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1136),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_315),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_170),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_893),
.Y(n_1863)
);

CKINVDCx20_ASAP7_75t_R g1864 ( 
.A(n_206),
.Y(n_1864)
);

BUFx10_ASAP7_75t_L g1865 ( 
.A(n_1041),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_336),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1088),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1074),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_949),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_468),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_322),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_276),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_891),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_207),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_365),
.Y(n_1875)
);

CKINVDCx16_ASAP7_75t_R g1876 ( 
.A(n_874),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_77),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1259),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_162),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1129),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1137),
.Y(n_1881)
);

CKINVDCx20_ASAP7_75t_R g1882 ( 
.A(n_50),
.Y(n_1882)
);

BUFx10_ASAP7_75t_L g1883 ( 
.A(n_1082),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_250),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1142),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_160),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1201),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_723),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_790),
.Y(n_1889)
);

INVx2_ASAP7_75t_SL g1890 ( 
.A(n_1153),
.Y(n_1890)
);

BUFx2_ASAP7_75t_SL g1891 ( 
.A(n_1119),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1230),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_718),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_114),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1243),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_487),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_999),
.Y(n_1897)
);

CKINVDCx20_ASAP7_75t_R g1898 ( 
.A(n_337),
.Y(n_1898)
);

CKINVDCx20_ASAP7_75t_R g1899 ( 
.A(n_167),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_486),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_914),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_281),
.Y(n_1902)
);

CKINVDCx20_ASAP7_75t_R g1903 ( 
.A(n_590),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_123),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_130),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_266),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_811),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1103),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1099),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_369),
.Y(n_1910)
);

CKINVDCx20_ASAP7_75t_R g1911 ( 
.A(n_586),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_721),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_44),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_457),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1118),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_731),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_158),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_282),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_463),
.Y(n_1919)
);

CKINVDCx20_ASAP7_75t_R g1920 ( 
.A(n_353),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_501),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_611),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1011),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_902),
.Y(n_1924)
);

CKINVDCx20_ASAP7_75t_R g1925 ( 
.A(n_899),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_1101),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_13),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_912),
.Y(n_1928)
);

BUFx10_ASAP7_75t_L g1929 ( 
.A(n_193),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_52),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_575),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_662),
.Y(n_1932)
);

BUFx2_ASAP7_75t_L g1933 ( 
.A(n_1251),
.Y(n_1933)
);

BUFx3_ASAP7_75t_L g1934 ( 
.A(n_1248),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1241),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_17),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_921),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_516),
.Y(n_1938)
);

CKINVDCx16_ASAP7_75t_R g1939 ( 
.A(n_929),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1231),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_267),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_876),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_630),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_679),
.Y(n_1944)
);

BUFx10_ASAP7_75t_L g1945 ( 
.A(n_429),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1086),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_900),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_450),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_885),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_267),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_179),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1214),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_701),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_761),
.Y(n_1954)
);

INVxp67_ASAP7_75t_L g1955 ( 
.A(n_1226),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_301),
.Y(n_1956)
);

BUFx3_ASAP7_75t_L g1957 ( 
.A(n_1164),
.Y(n_1957)
);

CKINVDCx14_ASAP7_75t_R g1958 ( 
.A(n_650),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_787),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_6),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_140),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1146),
.Y(n_1962)
);

CKINVDCx20_ASAP7_75t_R g1963 ( 
.A(n_1198),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_L g1964 ( 
.A(n_1195),
.Y(n_1964)
);

INVx2_ASAP7_75t_SL g1965 ( 
.A(n_637),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_474),
.Y(n_1966)
);

INVx1_ASAP7_75t_SL g1967 ( 
.A(n_32),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_26),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_930),
.Y(n_1969)
);

BUFx10_ASAP7_75t_L g1970 ( 
.A(n_945),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_551),
.Y(n_1971)
);

BUFx3_ASAP7_75t_L g1972 ( 
.A(n_587),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1116),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1112),
.Y(n_1974)
);

BUFx5_ASAP7_75t_L g1975 ( 
.A(n_847),
.Y(n_1975)
);

CKINVDCx20_ASAP7_75t_R g1976 ( 
.A(n_1172),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_303),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_928),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_636),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_828),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_324),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_948),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_526),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_764),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_959),
.Y(n_1985)
);

CKINVDCx20_ASAP7_75t_R g1986 ( 
.A(n_134),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_368),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_511),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_99),
.Y(n_1989)
);

CKINVDCx16_ASAP7_75t_R g1990 ( 
.A(n_939),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_401),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1147),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_918),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1252),
.Y(n_1994)
);

CKINVDCx20_ASAP7_75t_R g1995 ( 
.A(n_104),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_896),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_902),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1106),
.Y(n_1998)
);

INVx2_ASAP7_75t_SL g1999 ( 
.A(n_998),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_487),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_437),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_356),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1246),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_989),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_513),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_589),
.Y(n_2006)
);

INVx2_ASAP7_75t_SL g2007 ( 
.A(n_882),
.Y(n_2007)
);

BUFx6f_ASAP7_75t_L g2008 ( 
.A(n_1188),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_782),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_669),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_109),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_880),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_221),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_13),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_982),
.Y(n_2015)
);

BUFx10_ASAP7_75t_L g2016 ( 
.A(n_1204),
.Y(n_2016)
);

CKINVDCx20_ASAP7_75t_R g2017 ( 
.A(n_316),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_662),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_368),
.Y(n_2019)
);

INVx2_ASAP7_75t_SL g2020 ( 
.A(n_58),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_196),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_748),
.Y(n_2022)
);

CKINVDCx20_ASAP7_75t_R g2023 ( 
.A(n_1063),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_223),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_955),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_782),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_242),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_374),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_969),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_772),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_883),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_728),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_467),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_852),
.Y(n_2034)
);

CKINVDCx20_ASAP7_75t_R g2035 ( 
.A(n_1115),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_432),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1123),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_371),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1192),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_627),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_910),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_290),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_472),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_870),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_310),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1008),
.Y(n_2046)
);

INVx2_ASAP7_75t_SL g2047 ( 
.A(n_884),
.Y(n_2047)
);

CKINVDCx20_ASAP7_75t_R g2048 ( 
.A(n_922),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_1178),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_217),
.Y(n_2050)
);

INVx1_ASAP7_75t_SL g2051 ( 
.A(n_379),
.Y(n_2051)
);

BUFx10_ASAP7_75t_L g2052 ( 
.A(n_853),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1044),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_192),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_807),
.Y(n_2055)
);

BUFx10_ASAP7_75t_L g2056 ( 
.A(n_863),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_1216),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_779),
.Y(n_2058)
);

BUFx3_ASAP7_75t_L g2059 ( 
.A(n_766),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1064),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1104),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_427),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1133),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1223),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_858),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_69),
.Y(n_2066)
);

INVxp67_ASAP7_75t_L g2067 ( 
.A(n_164),
.Y(n_2067)
);

BUFx5_ASAP7_75t_L g2068 ( 
.A(n_1144),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_941),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_138),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_136),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_947),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_80),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_724),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_1145),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_920),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_395),
.Y(n_2077)
);

BUFx10_ASAP7_75t_L g2078 ( 
.A(n_911),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1648),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1648),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1315),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1288),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1288),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1288),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1288),
.Y(n_2085)
);

CKINVDCx16_ASAP7_75t_R g2086 ( 
.A(n_1323),
.Y(n_2086)
);

BUFx6f_ASAP7_75t_L g2087 ( 
.A(n_1338),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_1506),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1288),
.Y(n_2089)
);

INVxp67_ASAP7_75t_SL g2090 ( 
.A(n_1330),
.Y(n_2090)
);

INVxp67_ASAP7_75t_SL g2091 ( 
.A(n_1330),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1621),
.Y(n_2092)
);

BUFx3_ASAP7_75t_L g2093 ( 
.A(n_1469),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1621),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1621),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1621),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1665),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1621),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1646),
.Y(n_2099)
);

CKINVDCx16_ASAP7_75t_R g2100 ( 
.A(n_1726),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1646),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1646),
.Y(n_2102)
);

CKINVDCx16_ASAP7_75t_R g2103 ( 
.A(n_1732),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1646),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1646),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1782),
.Y(n_2106)
);

INVxp67_ASAP7_75t_SL g2107 ( 
.A(n_1330),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1782),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1782),
.Y(n_2109)
);

HB1xp67_ASAP7_75t_L g2110 ( 
.A(n_1475),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1782),
.Y(n_2111)
);

INVxp67_ASAP7_75t_SL g2112 ( 
.A(n_1344),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1782),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1975),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1975),
.Y(n_2115)
);

INVx3_ASAP7_75t_L g2116 ( 
.A(n_1278),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1975),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1975),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1975),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1282),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1283),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1958),
.B(n_0),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1287),
.Y(n_2123)
);

CKINVDCx20_ASAP7_75t_R g2124 ( 
.A(n_1270),
.Y(n_2124)
);

INVxp67_ASAP7_75t_SL g2125 ( 
.A(n_1344),
.Y(n_2125)
);

XOR2xp5_ASAP7_75t_L g2126 ( 
.A(n_1337),
.B(n_0),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1295),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1311),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_1343),
.Y(n_2129)
);

BUFx2_ASAP7_75t_L g2130 ( 
.A(n_1271),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1344),
.Y(n_2131)
);

INVxp67_ASAP7_75t_L g2132 ( 
.A(n_1375),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1314),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1321),
.Y(n_2134)
);

INVx2_ASAP7_75t_SL g2135 ( 
.A(n_2078),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1327),
.Y(n_2136)
);

CKINVDCx14_ASAP7_75t_R g2137 ( 
.A(n_1419),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1328),
.Y(n_2138)
);

INVx4_ASAP7_75t_R g2139 ( 
.A(n_1448),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1340),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1436),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1356),
.Y(n_2142)
);

INVxp33_ASAP7_75t_L g2143 ( 
.A(n_1960),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1357),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1359),
.Y(n_2145)
);

INVxp67_ASAP7_75t_SL g2146 ( 
.A(n_1436),
.Y(n_2146)
);

CKINVDCx14_ASAP7_75t_R g2147 ( 
.A(n_1596),
.Y(n_2147)
);

CKINVDCx16_ASAP7_75t_R g2148 ( 
.A(n_1876),
.Y(n_2148)
);

INVxp33_ASAP7_75t_L g2149 ( 
.A(n_1523),
.Y(n_2149)
);

INVxp67_ASAP7_75t_L g2150 ( 
.A(n_1676),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1367),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1374),
.Y(n_2152)
);

CKINVDCx16_ASAP7_75t_R g2153 ( 
.A(n_1939),
.Y(n_2153)
);

INVx2_ASAP7_75t_SL g2154 ( 
.A(n_2078),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1381),
.Y(n_2155)
);

CKINVDCx20_ASAP7_75t_R g2156 ( 
.A(n_1289),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1436),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1384),
.Y(n_2158)
);

BUFx3_ASAP7_75t_L g2159 ( 
.A(n_1518),
.Y(n_2159)
);

INVxp67_ASAP7_75t_L g2160 ( 
.A(n_1825),
.Y(n_2160)
);

CKINVDCx20_ASAP7_75t_R g2161 ( 
.A(n_1305),
.Y(n_2161)
);

INVxp33_ASAP7_75t_L g2162 ( 
.A(n_1833),
.Y(n_2162)
);

BUFx3_ASAP7_75t_L g2163 ( 
.A(n_1746),
.Y(n_2163)
);

BUFx3_ASAP7_75t_L g2164 ( 
.A(n_1845),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1386),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1387),
.Y(n_2166)
);

CKINVDCx20_ASAP7_75t_R g2167 ( 
.A(n_1332),
.Y(n_2167)
);

CKINVDCx20_ASAP7_75t_R g2168 ( 
.A(n_1342),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1393),
.Y(n_2169)
);

INVxp67_ASAP7_75t_L g2170 ( 
.A(n_1841),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1397),
.Y(n_2171)
);

INVxp67_ASAP7_75t_SL g2172 ( 
.A(n_1450),
.Y(n_2172)
);

INVxp67_ASAP7_75t_SL g2173 ( 
.A(n_1450),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1404),
.Y(n_2174)
);

BUFx2_ASAP7_75t_L g2175 ( 
.A(n_1990),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1405),
.Y(n_2176)
);

INVxp33_ASAP7_75t_SL g2177 ( 
.A(n_1346),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1450),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1428),
.Y(n_2179)
);

INVxp33_ASAP7_75t_SL g2180 ( 
.A(n_1272),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1432),
.Y(n_2181)
);

BUFx2_ASAP7_75t_SL g2182 ( 
.A(n_1269),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1443),
.Y(n_2183)
);

INVxp67_ASAP7_75t_L g2184 ( 
.A(n_1422),
.Y(n_2184)
);

INVxp67_ASAP7_75t_SL g2185 ( 
.A(n_1461),
.Y(n_2185)
);

INVxp67_ASAP7_75t_SL g2186 ( 
.A(n_1461),
.Y(n_2186)
);

INVxp67_ASAP7_75t_SL g2187 ( 
.A(n_1461),
.Y(n_2187)
);

CKINVDCx16_ASAP7_75t_R g2188 ( 
.A(n_1635),
.Y(n_2188)
);

INVxp33_ASAP7_75t_SL g2189 ( 
.A(n_1275),
.Y(n_2189)
);

CKINVDCx14_ASAP7_75t_R g2190 ( 
.A(n_1269),
.Y(n_2190)
);

INVxp67_ASAP7_75t_SL g2191 ( 
.A(n_1542),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1445),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1446),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1449),
.Y(n_2194)
);

CKINVDCx14_ASAP7_75t_R g2195 ( 
.A(n_1335),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1455),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1542),
.Y(n_2197)
);

CKINVDCx20_ASAP7_75t_R g2198 ( 
.A(n_1379),
.Y(n_2198)
);

CKINVDCx16_ASAP7_75t_R g2199 ( 
.A(n_1385),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1457),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1460),
.Y(n_2201)
);

INVxp33_ASAP7_75t_L g2202 ( 
.A(n_1519),
.Y(n_2202)
);

INVxp33_ASAP7_75t_SL g2203 ( 
.A(n_1279),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1464),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1467),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1542),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1470),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1473),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1474),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1481),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1487),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1493),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1503),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1532),
.Y(n_2214)
);

BUFx3_ASAP7_75t_L g2215 ( 
.A(n_1933),
.Y(n_2215)
);

INVxp67_ASAP7_75t_L g2216 ( 
.A(n_1814),
.Y(n_2216)
);

INVxp67_ASAP7_75t_SL g2217 ( 
.A(n_1589),
.Y(n_2217)
);

INVxp33_ASAP7_75t_SL g2218 ( 
.A(n_1284),
.Y(n_2218)
);

CKINVDCx16_ASAP7_75t_R g2219 ( 
.A(n_1385),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1533),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1538),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1543),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_1505),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1549),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1551),
.Y(n_2225)
);

CKINVDCx5p33_ASAP7_75t_R g2226 ( 
.A(n_1628),
.Y(n_2226)
);

INVxp33_ASAP7_75t_SL g2227 ( 
.A(n_1286),
.Y(n_2227)
);

CKINVDCx20_ASAP7_75t_R g2228 ( 
.A(n_1649),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1556),
.Y(n_2229)
);

INVxp33_ASAP7_75t_SL g2230 ( 
.A(n_1290),
.Y(n_2230)
);

CKINVDCx5p33_ASAP7_75t_R g2231 ( 
.A(n_1776),
.Y(n_2231)
);

INVxp67_ASAP7_75t_SL g2232 ( 
.A(n_1589),
.Y(n_2232)
);

INVxp67_ASAP7_75t_SL g2233 ( 
.A(n_1589),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1580),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1582),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_1963),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1583),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1601),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1602),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1612),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1623),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1720),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1624),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1625),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1627),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_2223),
.Y(n_2246)
);

HB1xp67_ASAP7_75t_L g2247 ( 
.A(n_2202),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2190),
.B(n_1335),
.Y(n_2248)
);

HB1xp67_ASAP7_75t_L g2249 ( 
.A(n_2175),
.Y(n_2249)
);

INVx5_ASAP7_75t_L g2250 ( 
.A(n_2199),
.Y(n_2250)
);

OAI22x1_ASAP7_75t_R g2251 ( 
.A1(n_2081),
.A2(n_1395),
.B1(n_1424),
.B2(n_1349),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2195),
.B(n_1514),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2087),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2090),
.Y(n_2254)
);

AOI22x1_ASAP7_75t_SL g2255 ( 
.A1(n_2124),
.A2(n_1444),
.B1(n_1494),
.B2(n_1437),
.Y(n_2255)
);

HB1xp67_ASAP7_75t_L g2256 ( 
.A(n_2088),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_2087),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2087),
.Y(n_2258)
);

AOI22x1_ASAP7_75t_SL g2259 ( 
.A1(n_2156),
.A2(n_1552),
.B1(n_1569),
.B2(n_1546),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2104),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2105),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_L g2262 ( 
.A(n_2180),
.B(n_2189),
.Y(n_2262)
);

BUFx2_ASAP7_75t_L g2263 ( 
.A(n_2097),
.Y(n_2263)
);

OAI22xp5_ASAP7_75t_SL g2264 ( 
.A1(n_2126),
.A2(n_1637),
.B1(n_1659),
.B2(n_1617),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2091),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_L g2266 ( 
.A1(n_2119),
.A2(n_2083),
.B(n_2082),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2131),
.Y(n_2267)
);

BUFx6f_ASAP7_75t_L g2268 ( 
.A(n_2141),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2107),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2112),
.Y(n_2270)
);

BUFx6f_ASAP7_75t_L g2271 ( 
.A(n_2157),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_2178),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_2226),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2197),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2125),
.Y(n_2275)
);

BUFx6f_ASAP7_75t_L g2276 ( 
.A(n_2206),
.Y(n_2276)
);

INVx4_ASAP7_75t_L g2277 ( 
.A(n_2086),
.Y(n_2277)
);

AOI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2122),
.A2(n_2150),
.B1(n_2160),
.B2(n_2132),
.Y(n_2278)
);

HB1xp67_ASAP7_75t_L g2279 ( 
.A(n_2148),
.Y(n_2279)
);

INVx3_ASAP7_75t_L g2280 ( 
.A(n_2116),
.Y(n_2280)
);

INVx4_ASAP7_75t_L g2281 ( 
.A(n_2100),
.Y(n_2281)
);

INVx5_ASAP7_75t_L g2282 ( 
.A(n_2219),
.Y(n_2282)
);

HB1xp67_ASAP7_75t_L g2283 ( 
.A(n_2153),
.Y(n_2283)
);

INVxp67_ASAP7_75t_L g2284 ( 
.A(n_2182),
.Y(n_2284)
);

BUFx6f_ASAP7_75t_L g2285 ( 
.A(n_2242),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2146),
.Y(n_2286)
);

BUFx6f_ASAP7_75t_L g2287 ( 
.A(n_2116),
.Y(n_2287)
);

BUFx6f_ASAP7_75t_L g2288 ( 
.A(n_2129),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_2103),
.B(n_1514),
.Y(n_2289)
);

BUFx6f_ASAP7_75t_L g2290 ( 
.A(n_2129),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_L g2291 ( 
.A(n_2120),
.Y(n_2291)
);

BUFx6f_ASAP7_75t_L g2292 ( 
.A(n_2121),
.Y(n_2292)
);

INVx5_ASAP7_75t_L g2293 ( 
.A(n_2130),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2172),
.Y(n_2294)
);

HB1xp67_ASAP7_75t_L g2295 ( 
.A(n_2184),
.Y(n_2295)
);

CKINVDCx20_ASAP7_75t_R g2296 ( 
.A(n_2161),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2173),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2084),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2085),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_2123),
.Y(n_2300)
);

INVx5_ASAP7_75t_L g2301 ( 
.A(n_2135),
.Y(n_2301)
);

INVx6_ASAP7_75t_L g2302 ( 
.A(n_2093),
.Y(n_2302)
);

BUFx8_ASAP7_75t_SL g2303 ( 
.A(n_2167),
.Y(n_2303)
);

INVxp33_ASAP7_75t_SL g2304 ( 
.A(n_2231),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2185),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_2236),
.Y(n_2306)
);

INVx6_ASAP7_75t_L g2307 ( 
.A(n_2159),
.Y(n_2307)
);

BUFx8_ASAP7_75t_SL g2308 ( 
.A(n_2168),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2186),
.Y(n_2309)
);

AND2x6_ASAP7_75t_L g2310 ( 
.A(n_2163),
.B(n_1832),
.Y(n_2310)
);

CKINVDCx20_ASAP7_75t_R g2311 ( 
.A(n_2198),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2187),
.Y(n_2312)
);

BUFx6f_ASAP7_75t_L g2313 ( 
.A(n_2127),
.Y(n_2313)
);

AND2x4_ASAP7_75t_L g2314 ( 
.A(n_2164),
.B(n_1910),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2191),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2137),
.B(n_1715),
.Y(n_2316)
);

HB1xp67_ASAP7_75t_L g2317 ( 
.A(n_2216),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2217),
.Y(n_2318)
);

AND2x4_ASAP7_75t_L g2319 ( 
.A(n_2215),
.B(n_1972),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2089),
.Y(n_2320)
);

HB1xp67_ASAP7_75t_L g2321 ( 
.A(n_2170),
.Y(n_2321)
);

BUFx6f_ASAP7_75t_L g2322 ( 
.A(n_2128),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_2188),
.B(n_1715),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2232),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2233),
.Y(n_2325)
);

BUFx6f_ASAP7_75t_L g2326 ( 
.A(n_2133),
.Y(n_2326)
);

OAI22x1_ASAP7_75t_SL g2327 ( 
.A1(n_2228),
.A2(n_1688),
.B1(n_1696),
.B2(n_1666),
.Y(n_2327)
);

BUFx6f_ASAP7_75t_L g2328 ( 
.A(n_2134),
.Y(n_2328)
);

INVx3_ASAP7_75t_L g2329 ( 
.A(n_2136),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2079),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2092),
.Y(n_2331)
);

INVx3_ASAP7_75t_L g2332 ( 
.A(n_2138),
.Y(n_2332)
);

INVx6_ASAP7_75t_L g2333 ( 
.A(n_2177),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2080),
.Y(n_2334)
);

INVx5_ASAP7_75t_L g2335 ( 
.A(n_2154),
.Y(n_2335)
);

BUFx6f_ASAP7_75t_L g2336 ( 
.A(n_2140),
.Y(n_2336)
);

CKINVDCx5p33_ASAP7_75t_R g2337 ( 
.A(n_2203),
.Y(n_2337)
);

BUFx2_ASAP7_75t_L g2338 ( 
.A(n_2110),
.Y(n_2338)
);

INVx4_ASAP7_75t_L g2339 ( 
.A(n_2094),
.Y(n_2339)
);

OAI22x1_ASAP7_75t_R g2340 ( 
.A1(n_2142),
.A2(n_1721),
.B1(n_1733),
.B2(n_1699),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2147),
.B(n_1409),
.Y(n_2341)
);

INVx6_ASAP7_75t_L g2342 ( 
.A(n_2149),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2162),
.B(n_1865),
.Y(n_2343)
);

INVx3_ASAP7_75t_L g2344 ( 
.A(n_2144),
.Y(n_2344)
);

HB1xp67_ASAP7_75t_L g2345 ( 
.A(n_2143),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2095),
.Y(n_2346)
);

OA21x2_ASAP7_75t_L g2347 ( 
.A1(n_2096),
.A2(n_1285),
.B(n_1267),
.Y(n_2347)
);

OAI21x1_ASAP7_75t_L g2348 ( 
.A1(n_2098),
.A2(n_1353),
.B(n_1316),
.Y(n_2348)
);

BUFx2_ASAP7_75t_L g2349 ( 
.A(n_2145),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2151),
.B(n_2152),
.Y(n_2350)
);

OA21x2_ASAP7_75t_L g2351 ( 
.A1(n_2099),
.A2(n_1390),
.B(n_1355),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2155),
.B(n_2158),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2165),
.B(n_1865),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2101),
.Y(n_2354)
);

HB1xp67_ASAP7_75t_L g2355 ( 
.A(n_2218),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2227),
.B(n_1685),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2102),
.B(n_1411),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2166),
.B(n_1883),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2106),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2169),
.B(n_1883),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2108),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2109),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2111),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2113),
.B(n_1413),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2114),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_L g2366 ( 
.A(n_2230),
.B(n_1276),
.Y(n_2366)
);

BUFx12f_ASAP7_75t_L g2367 ( 
.A(n_2139),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_2171),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2115),
.Y(n_2369)
);

BUFx12f_ASAP7_75t_L g2370 ( 
.A(n_2174),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2117),
.Y(n_2371)
);

HB1xp67_ASAP7_75t_L g2372 ( 
.A(n_2176),
.Y(n_2372)
);

INVx4_ASAP7_75t_L g2373 ( 
.A(n_2118),
.Y(n_2373)
);

INVxp67_ASAP7_75t_L g2374 ( 
.A(n_2179),
.Y(n_2374)
);

OA21x2_ASAP7_75t_L g2375 ( 
.A1(n_2181),
.A2(n_1454),
.B(n_1418),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_2183),
.B(n_2059),
.Y(n_2376)
);

BUFx6f_ASAP7_75t_L g2377 ( 
.A(n_2192),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2193),
.B(n_1459),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2194),
.Y(n_2379)
);

INVx5_ASAP7_75t_L g2380 ( 
.A(n_2196),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2200),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2201),
.Y(n_2382)
);

BUFx3_ASAP7_75t_L g2383 ( 
.A(n_2204),
.Y(n_2383)
);

AND2x4_ASAP7_75t_L g2384 ( 
.A(n_2205),
.B(n_2077),
.Y(n_2384)
);

BUFx2_ASAP7_75t_L g2385 ( 
.A(n_2207),
.Y(n_2385)
);

BUFx12f_ASAP7_75t_L g2386 ( 
.A(n_2208),
.Y(n_2386)
);

BUFx3_ASAP7_75t_L g2387 ( 
.A(n_2209),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2210),
.B(n_2211),
.Y(n_2388)
);

BUFx6f_ASAP7_75t_L g2389 ( 
.A(n_2212),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2213),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2214),
.Y(n_2391)
);

INVx5_ASAP7_75t_L g2392 ( 
.A(n_2220),
.Y(n_2392)
);

BUFx12f_ASAP7_75t_L g2393 ( 
.A(n_2221),
.Y(n_2393)
);

INVx5_ASAP7_75t_L g2394 ( 
.A(n_2222),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2224),
.Y(n_2395)
);

BUFx3_ASAP7_75t_L g2396 ( 
.A(n_2225),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_L g2397 ( 
.A(n_2229),
.Y(n_2397)
);

BUFx3_ASAP7_75t_L g2398 ( 
.A(n_2234),
.Y(n_2398)
);

AOI22x1_ASAP7_75t_SL g2399 ( 
.A1(n_2235),
.A2(n_1789),
.B1(n_1800),
.B2(n_1750),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2237),
.Y(n_2400)
);

BUFx12f_ASAP7_75t_L g2401 ( 
.A(n_2238),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_2239),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2240),
.B(n_2016),
.Y(n_2403)
);

INVx3_ASAP7_75t_L g2404 ( 
.A(n_2241),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_2243),
.B(n_1399),
.Y(n_2405)
);

BUFx6f_ASAP7_75t_L g2406 ( 
.A(n_2244),
.Y(n_2406)
);

BUFx8_ASAP7_75t_SL g2407 ( 
.A(n_2245),
.Y(n_2407)
);

INVx4_ASAP7_75t_L g2408 ( 
.A(n_2087),
.Y(n_2408)
);

BUFx6f_ASAP7_75t_L g2409 ( 
.A(n_2087),
.Y(n_2409)
);

BUFx6f_ASAP7_75t_L g2410 ( 
.A(n_2087),
.Y(n_2410)
);

INVx5_ASAP7_75t_L g2411 ( 
.A(n_2199),
.Y(n_2411)
);

BUFx6f_ASAP7_75t_L g2412 ( 
.A(n_2087),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2090),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2090),
.Y(n_2414)
);

BUFx6f_ASAP7_75t_L g2415 ( 
.A(n_2087),
.Y(n_2415)
);

OAI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2202),
.A2(n_1821),
.B1(n_1830),
.B2(n_1813),
.Y(n_2416)
);

OA21x2_ASAP7_75t_L g2417 ( 
.A1(n_2082),
.A2(n_1476),
.B(n_1466),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2090),
.Y(n_2418)
);

AOI22x1_ASAP7_75t_SL g2419 ( 
.A1(n_2124),
.A2(n_1864),
.B1(n_1882),
.B2(n_1847),
.Y(n_2419)
);

BUFx6f_ASAP7_75t_L g2420 ( 
.A(n_2087),
.Y(n_2420)
);

BUFx12f_ASAP7_75t_L g2421 ( 
.A(n_2081),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2090),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2093),
.B(n_1495),
.Y(n_2423)
);

BUFx6f_ASAP7_75t_L g2424 ( 
.A(n_2087),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2202),
.B(n_2016),
.Y(n_2425)
);

NOR2x1_ASAP7_75t_L g2426 ( 
.A(n_2182),
.B(n_1690),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2090),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2087),
.Y(n_2428)
);

HB1xp67_ASAP7_75t_L g2429 ( 
.A(n_2202),
.Y(n_2429)
);

CKINVDCx5p33_ASAP7_75t_R g2430 ( 
.A(n_2223),
.Y(n_2430)
);

AND2x4_ASAP7_75t_L g2431 ( 
.A(n_2093),
.B(n_1787),
.Y(n_2431)
);

BUFx8_ASAP7_75t_SL g2432 ( 
.A(n_2124),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_2093),
.B(n_1797),
.Y(n_2433)
);

INVxp67_ASAP7_75t_L g2434 ( 
.A(n_2182),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_2087),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2090),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2087),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2087),
.Y(n_2438)
);

INVx5_ASAP7_75t_L g2439 ( 
.A(n_2199),
.Y(n_2439)
);

BUFx6f_ASAP7_75t_L g2440 ( 
.A(n_2087),
.Y(n_2440)
);

INVx3_ASAP7_75t_L g2441 ( 
.A(n_2116),
.Y(n_2441)
);

OA21x2_ASAP7_75t_L g2442 ( 
.A1(n_2082),
.A2(n_1485),
.B(n_1477),
.Y(n_2442)
);

AOI22x1_ASAP7_75t_SL g2443 ( 
.A1(n_2124),
.A2(n_1899),
.B1(n_1903),
.B2(n_1898),
.Y(n_2443)
);

BUFx3_ASAP7_75t_L g2444 ( 
.A(n_2116),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2093),
.B(n_1804),
.Y(n_2445)
);

BUFx6f_ASAP7_75t_L g2446 ( 
.A(n_2087),
.Y(n_2446)
);

AOI22xp5_ASAP7_75t_L g2447 ( 
.A1(n_2202),
.A2(n_1920),
.B1(n_1925),
.B2(n_1911),
.Y(n_2447)
);

INVxp67_ASAP7_75t_SL g2448 ( 
.A(n_2184),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2087),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2087),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2090),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_2086),
.B(n_1513),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2087),
.Y(n_2453)
);

BUFx8_ASAP7_75t_L g2454 ( 
.A(n_2175),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2087),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2087),
.Y(n_2456)
);

BUFx8_ASAP7_75t_L g2457 ( 
.A(n_2175),
.Y(n_2457)
);

BUFx6f_ASAP7_75t_L g2458 ( 
.A(n_2087),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2202),
.B(n_1442),
.Y(n_2459)
);

HB1xp67_ASAP7_75t_L g2460 ( 
.A(n_2202),
.Y(n_2460)
);

BUFx6f_ASAP7_75t_L g2461 ( 
.A(n_2087),
.Y(n_2461)
);

INVx3_ASAP7_75t_L g2462 ( 
.A(n_2116),
.Y(n_2462)
);

INVx5_ASAP7_75t_L g2463 ( 
.A(n_2086),
.Y(n_2463)
);

OAI21x1_ASAP7_75t_L g2464 ( 
.A1(n_2104),
.A2(n_1535),
.B(n_1509),
.Y(n_2464)
);

BUFx2_ASAP7_75t_L g2465 ( 
.A(n_2088),
.Y(n_2465)
);

BUFx2_ASAP7_75t_L g2466 ( 
.A(n_2088),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2090),
.Y(n_2467)
);

BUFx2_ASAP7_75t_L g2468 ( 
.A(n_2088),
.Y(n_2468)
);

HB1xp67_ASAP7_75t_L g2469 ( 
.A(n_2202),
.Y(n_2469)
);

BUFx12f_ASAP7_75t_L g2470 ( 
.A(n_2081),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2090),
.Y(n_2471)
);

BUFx6f_ASAP7_75t_L g2472 ( 
.A(n_2087),
.Y(n_2472)
);

BUFx12f_ASAP7_75t_L g2473 ( 
.A(n_2081),
.Y(n_2473)
);

BUFx6f_ASAP7_75t_L g2474 ( 
.A(n_2087),
.Y(n_2474)
);

BUFx12f_ASAP7_75t_L g2475 ( 
.A(n_2081),
.Y(n_2475)
);

BUFx8_ASAP7_75t_SL g2476 ( 
.A(n_2124),
.Y(n_2476)
);

INVx5_ASAP7_75t_L g2477 ( 
.A(n_2199),
.Y(n_2477)
);

BUFx8_ASAP7_75t_SL g2478 ( 
.A(n_2124),
.Y(n_2478)
);

BUFx2_ASAP7_75t_L g2479 ( 
.A(n_2088),
.Y(n_2479)
);

INVx3_ASAP7_75t_L g2480 ( 
.A(n_2116),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2090),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_2202),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2137),
.B(n_1536),
.Y(n_2483)
);

OAI21x1_ASAP7_75t_L g2484 ( 
.A1(n_2104),
.A2(n_1560),
.B(n_1547),
.Y(n_2484)
);

BUFx6f_ASAP7_75t_L g2485 ( 
.A(n_2087),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2090),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_2087),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2137),
.B(n_1566),
.Y(n_2488)
);

AND2x4_ASAP7_75t_L g2489 ( 
.A(n_2093),
.B(n_1834),
.Y(n_2489)
);

BUFx12f_ASAP7_75t_L g2490 ( 
.A(n_2081),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2137),
.B(n_1605),
.Y(n_2491)
);

HB1xp67_ASAP7_75t_L g2492 ( 
.A(n_2202),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2090),
.Y(n_2493)
);

INVx5_ASAP7_75t_L g2494 ( 
.A(n_2199),
.Y(n_2494)
);

BUFx2_ASAP7_75t_L g2495 ( 
.A(n_2088),
.Y(n_2495)
);

AOI22xp5_ASAP7_75t_L g2496 ( 
.A1(n_2202),
.A2(n_1986),
.B1(n_2017),
.B2(n_1995),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2087),
.Y(n_2497)
);

BUFx12f_ASAP7_75t_L g2498 ( 
.A(n_2081),
.Y(n_2498)
);

AND2x4_ASAP7_75t_L g2499 ( 
.A(n_2093),
.B(n_1965),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2090),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2137),
.B(n_1609),
.Y(n_2501)
);

OA21x2_ASAP7_75t_L g2502 ( 
.A1(n_2082),
.A2(n_1622),
.B(n_1613),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2087),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2087),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2087),
.Y(n_2505)
);

HB1xp67_ASAP7_75t_L g2506 ( 
.A(n_2202),
.Y(n_2506)
);

BUFx8_ASAP7_75t_SL g2507 ( 
.A(n_2124),
.Y(n_2507)
);

BUFx6f_ASAP7_75t_L g2508 ( 
.A(n_2087),
.Y(n_2508)
);

BUFx6f_ASAP7_75t_L g2509 ( 
.A(n_2087),
.Y(n_2509)
);

AND2x6_ASAP7_75t_L g2510 ( 
.A(n_2122),
.B(n_1720),
.Y(n_2510)
);

BUFx6f_ASAP7_75t_L g2511 ( 
.A(n_2087),
.Y(n_2511)
);

INVx2_ASAP7_75t_SL g2512 ( 
.A(n_2093),
.Y(n_2512)
);

AOI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_2202),
.A2(n_2048),
.B1(n_2023),
.B2(n_2035),
.Y(n_2513)
);

CKINVDCx5p33_ASAP7_75t_R g2514 ( 
.A(n_2223),
.Y(n_2514)
);

AND2x4_ASAP7_75t_L g2515 ( 
.A(n_2093),
.B(n_2007),
.Y(n_2515)
);

CKINVDCx5p33_ASAP7_75t_R g2516 ( 
.A(n_2223),
.Y(n_2516)
);

BUFx3_ASAP7_75t_L g2517 ( 
.A(n_2116),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_L g2518 ( 
.A(n_2180),
.B(n_1844),
.Y(n_2518)
);

AND2x4_ASAP7_75t_L g2519 ( 
.A(n_2093),
.B(n_2020),
.Y(n_2519)
);

BUFx12f_ASAP7_75t_L g2520 ( 
.A(n_2081),
.Y(n_2520)
);

BUFx3_ASAP7_75t_L g2521 ( 
.A(n_2116),
.Y(n_2521)
);

BUFx8_ASAP7_75t_SL g2522 ( 
.A(n_2124),
.Y(n_2522)
);

BUFx6f_ASAP7_75t_L g2523 ( 
.A(n_2087),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2087),
.Y(n_2524)
);

BUFx3_ASAP7_75t_L g2525 ( 
.A(n_2116),
.Y(n_2525)
);

NOR2xp33_ASAP7_75t_L g2526 ( 
.A(n_2180),
.B(n_1955),
.Y(n_2526)
);

HB1xp67_ASAP7_75t_L g2527 ( 
.A(n_2202),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2137),
.B(n_1626),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_L g2529 ( 
.A(n_2180),
.B(n_1647),
.Y(n_2529)
);

INVx3_ASAP7_75t_L g2530 ( 
.A(n_2116),
.Y(n_2530)
);

AND2x4_ASAP7_75t_L g2531 ( 
.A(n_2093),
.B(n_2047),
.Y(n_2531)
);

BUFx12f_ASAP7_75t_L g2532 ( 
.A(n_2081),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2090),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2087),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2137),
.B(n_1704),
.Y(n_2535)
);

OAI21x1_ASAP7_75t_L g2536 ( 
.A1(n_2104),
.A2(n_1728),
.B(n_1716),
.Y(n_2536)
);

BUFx3_ASAP7_75t_L g2537 ( 
.A(n_2116),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2090),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2090),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2090),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2087),
.Y(n_2541)
);

BUFx6f_ASAP7_75t_L g2542 ( 
.A(n_2087),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2090),
.Y(n_2543)
);

BUFx6f_ASAP7_75t_L g2544 ( 
.A(n_2087),
.Y(n_2544)
);

BUFx3_ASAP7_75t_L g2545 ( 
.A(n_2116),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2090),
.Y(n_2546)
);

BUFx6f_ASAP7_75t_L g2547 ( 
.A(n_2087),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2087),
.Y(n_2548)
);

INVxp33_ASAP7_75t_SL g2549 ( 
.A(n_2223),
.Y(n_2549)
);

NOR2xp67_ASAP7_75t_L g2550 ( 
.A(n_2184),
.B(n_1579),
.Y(n_2550)
);

AOI22x1_ASAP7_75t_SL g2551 ( 
.A1(n_2124),
.A2(n_1292),
.B1(n_1296),
.B2(n_1291),
.Y(n_2551)
);

XOR2xp5_ASAP7_75t_L g2552 ( 
.A(n_2124),
.B(n_1976),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2087),
.Y(n_2553)
);

BUFx6f_ASAP7_75t_L g2554 ( 
.A(n_2087),
.Y(n_2554)
);

AND2x4_ASAP7_75t_L g2555 ( 
.A(n_2093),
.B(n_1755),
.Y(n_2555)
);

INVx6_ASAP7_75t_L g2556 ( 
.A(n_2199),
.Y(n_2556)
);

BUFx8_ASAP7_75t_SL g2557 ( 
.A(n_2124),
.Y(n_2557)
);

AND2x4_ASAP7_75t_L g2558 ( 
.A(n_2093),
.B(n_1769),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2090),
.Y(n_2559)
);

AND2x4_ASAP7_75t_L g2560 ( 
.A(n_2093),
.B(n_2067),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2087),
.Y(n_2561)
);

INVx3_ASAP7_75t_L g2562 ( 
.A(n_2116),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2090),
.Y(n_2563)
);

BUFx2_ASAP7_75t_L g2564 ( 
.A(n_2088),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_2223),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_SL g2566 ( 
.A(n_2188),
.B(n_1298),
.Y(n_2566)
);

NOR2xp33_ASAP7_75t_L g2567 ( 
.A(n_2180),
.B(n_1738),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2090),
.Y(n_2568)
);

BUFx3_ASAP7_75t_L g2569 ( 
.A(n_2116),
.Y(n_2569)
);

INVxp67_ASAP7_75t_L g2570 ( 
.A(n_2182),
.Y(n_2570)
);

INVx4_ASAP7_75t_L g2571 ( 
.A(n_2087),
.Y(n_2571)
);

BUFx12f_ASAP7_75t_L g2572 ( 
.A(n_2081),
.Y(n_2572)
);

BUFx8_ASAP7_75t_SL g2573 ( 
.A(n_2124),
.Y(n_2573)
);

CKINVDCx5p33_ASAP7_75t_R g2574 ( 
.A(n_2303),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_2573),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2330),
.Y(n_2576)
);

INVx1_ASAP7_75t_SL g2577 ( 
.A(n_2342),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_2308),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2334),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2381),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2247),
.B(n_1442),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2260),
.Y(n_2582)
);

OA21x2_ASAP7_75t_L g2583 ( 
.A1(n_2348),
.A2(n_1748),
.B(n_1747),
.Y(n_2583)
);

INVx3_ASAP7_75t_L g2584 ( 
.A(n_2287),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2382),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2400),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2353),
.B(n_1273),
.Y(n_2587)
);

BUFx2_ASAP7_75t_L g2588 ( 
.A(n_2429),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2291),
.Y(n_2589)
);

CKINVDCx5p33_ASAP7_75t_R g2590 ( 
.A(n_2432),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2261),
.Y(n_2591)
);

CKINVDCx5p33_ASAP7_75t_R g2592 ( 
.A(n_2476),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_2478),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2268),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_2507),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2358),
.B(n_1319),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2292),
.Y(n_2597)
);

CKINVDCx5p33_ASAP7_75t_R g2598 ( 
.A(n_2522),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2360),
.B(n_2403),
.Y(n_2599)
);

CKINVDCx5p33_ASAP7_75t_R g2600 ( 
.A(n_2557),
.Y(n_2600)
);

CKINVDCx6p67_ASAP7_75t_R g2601 ( 
.A(n_2421),
.Y(n_2601)
);

NOR2xp33_ASAP7_75t_L g2602 ( 
.A(n_2339),
.B(n_1749),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2300),
.Y(n_2603)
);

CKINVDCx20_ASAP7_75t_R g2604 ( 
.A(n_2296),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2313),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2322),
.Y(n_2606)
);

OA21x2_ASAP7_75t_L g2607 ( 
.A1(n_2464),
.A2(n_1796),
.B(n_1751),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2326),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_2246),
.Y(n_2609)
);

BUFx3_ASAP7_75t_L g2610 ( 
.A(n_2367),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_2273),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2271),
.Y(n_2612)
);

NAND2xp33_ASAP7_75t_SL g2613 ( 
.A(n_2337),
.B(n_1299),
.Y(n_2613)
);

CKINVDCx5p33_ASAP7_75t_R g2614 ( 
.A(n_2306),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2460),
.B(n_1479),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2328),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2336),
.Y(n_2617)
);

CKINVDCx5p33_ASAP7_75t_R g2618 ( 
.A(n_2430),
.Y(n_2618)
);

CKINVDCx16_ASAP7_75t_R g2619 ( 
.A(n_2469),
.Y(n_2619)
);

BUFx6f_ASAP7_75t_L g2620 ( 
.A(n_2288),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2272),
.Y(n_2621)
);

AND2x4_ASAP7_75t_L g2622 ( 
.A(n_2482),
.B(n_1303),
.Y(n_2622)
);

CKINVDCx5p33_ASAP7_75t_R g2623 ( 
.A(n_2514),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2492),
.B(n_1479),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2276),
.Y(n_2625)
);

CKINVDCx20_ASAP7_75t_R g2626 ( 
.A(n_2311),
.Y(n_2626)
);

INVx3_ASAP7_75t_L g2627 ( 
.A(n_2290),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2285),
.Y(n_2628)
);

CKINVDCx6p67_ASAP7_75t_R g2629 ( 
.A(n_2470),
.Y(n_2629)
);

CKINVDCx5p33_ASAP7_75t_R g2630 ( 
.A(n_2516),
.Y(n_2630)
);

CKINVDCx5p33_ASAP7_75t_R g2631 ( 
.A(n_2565),
.Y(n_2631)
);

CKINVDCx20_ASAP7_75t_R g2632 ( 
.A(n_2552),
.Y(n_2632)
);

AND3x1_ASAP7_75t_L g2633 ( 
.A(n_2356),
.B(n_1645),
.C(n_1638),
.Y(n_2633)
);

CKINVDCx20_ASAP7_75t_R g2634 ( 
.A(n_2506),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_R g2635 ( 
.A(n_2473),
.B(n_2475),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2368),
.Y(n_2636)
);

AND2x6_ASAP7_75t_L g2637 ( 
.A(n_2248),
.B(n_1799),
.Y(n_2637)
);

NOR2xp33_ASAP7_75t_L g2638 ( 
.A(n_2373),
.B(n_1802),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_2304),
.Y(n_2639)
);

BUFx6f_ASAP7_75t_L g2640 ( 
.A(n_2257),
.Y(n_2640)
);

BUFx2_ASAP7_75t_L g2641 ( 
.A(n_2527),
.Y(n_2641)
);

CKINVDCx5p33_ASAP7_75t_R g2642 ( 
.A(n_2549),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2377),
.Y(n_2643)
);

CKINVDCx5p33_ASAP7_75t_R g2644 ( 
.A(n_2490),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2389),
.Y(n_2645)
);

BUFx6f_ASAP7_75t_L g2646 ( 
.A(n_2409),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2345),
.B(n_1486),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_2498),
.Y(n_2648)
);

INVxp67_ASAP7_75t_L g2649 ( 
.A(n_2425),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2397),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2266),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2402),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2529),
.B(n_2567),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_2267),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2406),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2379),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2390),
.Y(n_2657)
);

CKINVDCx20_ASAP7_75t_R g2658 ( 
.A(n_2454),
.Y(n_2658)
);

HB1xp67_ASAP7_75t_L g2659 ( 
.A(n_2249),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2391),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_2520),
.Y(n_2661)
);

CKINVDCx5p33_ASAP7_75t_R g2662 ( 
.A(n_2532),
.Y(n_2662)
);

INVx5_ASAP7_75t_L g2663 ( 
.A(n_2556),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2366),
.B(n_2518),
.Y(n_2664)
);

HB1xp67_ASAP7_75t_L g2665 ( 
.A(n_2459),
.Y(n_2665)
);

BUFx3_ASAP7_75t_L g2666 ( 
.A(n_2444),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2395),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2346),
.Y(n_2668)
);

OAI22xp5_ASAP7_75t_SL g2669 ( 
.A1(n_2264),
.A2(n_1578),
.B1(n_1672),
.B2(n_1308),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_2572),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2274),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2354),
.Y(n_2672)
);

BUFx6f_ASAP7_75t_L g2673 ( 
.A(n_2410),
.Y(n_2673)
);

AND2x4_ASAP7_75t_L g2674 ( 
.A(n_2463),
.B(n_1717),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2343),
.B(n_1486),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2253),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2526),
.B(n_1324),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2361),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2258),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2263),
.Y(n_2680)
);

CKINVDCx5p33_ASAP7_75t_R g2681 ( 
.A(n_2465),
.Y(n_2681)
);

CKINVDCx20_ASAP7_75t_R g2682 ( 
.A(n_2457),
.Y(n_2682)
);

BUFx2_ASAP7_75t_L g2683 ( 
.A(n_2279),
.Y(n_2683)
);

CKINVDCx5p33_ASAP7_75t_R g2684 ( 
.A(n_2466),
.Y(n_2684)
);

BUFx3_ASAP7_75t_L g2685 ( 
.A(n_2517),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_2468),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2362),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2428),
.Y(n_2688)
);

CKINVDCx5p33_ASAP7_75t_R g2689 ( 
.A(n_2479),
.Y(n_2689)
);

CKINVDCx5p33_ASAP7_75t_R g2690 ( 
.A(n_2495),
.Y(n_2690)
);

CKINVDCx5p33_ASAP7_75t_R g2691 ( 
.A(n_2564),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2437),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_2355),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2365),
.Y(n_2694)
);

AND2x4_ASAP7_75t_L g2695 ( 
.A(n_2463),
.B(n_1768),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2254),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2265),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2298),
.B(n_1348),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2269),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2321),
.B(n_1499),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2438),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_2333),
.Y(n_2702)
);

CKINVDCx5p33_ASAP7_75t_R g2703 ( 
.A(n_2416),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2270),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2275),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2286),
.Y(n_2706)
);

OA21x2_ASAP7_75t_L g2707 ( 
.A1(n_2484),
.A2(n_1827),
.B(n_1820),
.Y(n_2707)
);

BUFx6f_ASAP7_75t_L g2708 ( 
.A(n_2412),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2294),
.Y(n_2709)
);

CKINVDCx5p33_ASAP7_75t_R g2710 ( 
.A(n_2250),
.Y(n_2710)
);

HB1xp67_ASAP7_75t_L g2711 ( 
.A(n_2283),
.Y(n_2711)
);

CKINVDCx5p33_ASAP7_75t_R g2712 ( 
.A(n_2282),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2297),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2305),
.Y(n_2714)
);

BUFx3_ASAP7_75t_L g2715 ( 
.A(n_2521),
.Y(n_2715)
);

INVx3_ASAP7_75t_L g2716 ( 
.A(n_2302),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2295),
.B(n_1499),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2449),
.Y(n_2718)
);

CKINVDCx20_ASAP7_75t_R g2719 ( 
.A(n_2256),
.Y(n_2719)
);

AND2x4_ASAP7_75t_L g2720 ( 
.A(n_2512),
.B(n_1829),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2450),
.Y(n_2721)
);

BUFx10_ASAP7_75t_L g2722 ( 
.A(n_2262),
.Y(n_2722)
);

BUFx6f_ASAP7_75t_L g2723 ( 
.A(n_2415),
.Y(n_2723)
);

CKINVDCx5p33_ASAP7_75t_R g2724 ( 
.A(n_2411),
.Y(n_2724)
);

CKINVDCx5p33_ASAP7_75t_R g2725 ( 
.A(n_2439),
.Y(n_2725)
);

BUFx6f_ASAP7_75t_L g2726 ( 
.A(n_2420),
.Y(n_2726)
);

BUFx6f_ASAP7_75t_L g2727 ( 
.A(n_2424),
.Y(n_2727)
);

AND2x4_ASAP7_75t_L g2728 ( 
.A(n_2477),
.B(n_1862),
.Y(n_2728)
);

NOR2xp33_ASAP7_75t_R g2729 ( 
.A(n_2494),
.B(n_1268),
.Y(n_2729)
);

BUFx2_ASAP7_75t_L g2730 ( 
.A(n_2338),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2309),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2453),
.Y(n_2732)
);

CKINVDCx5p33_ASAP7_75t_R g2733 ( 
.A(n_2307),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2312),
.Y(n_2734)
);

NOR2xp33_ASAP7_75t_SL g2735 ( 
.A(n_2566),
.B(n_1884),
.Y(n_2735)
);

HB1xp67_ASAP7_75t_L g2736 ( 
.A(n_2317),
.Y(n_2736)
);

CKINVDCx20_ASAP7_75t_R g2737 ( 
.A(n_2277),
.Y(n_2737)
);

NAND2xp33_ASAP7_75t_SL g2738 ( 
.A(n_2281),
.B(n_1300),
.Y(n_2738)
);

BUFx3_ASAP7_75t_L g2739 ( 
.A(n_2525),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_2407),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2455),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2315),
.Y(n_2742)
);

HB1xp67_ASAP7_75t_L g2743 ( 
.A(n_2293),
.Y(n_2743)
);

INVx3_ASAP7_75t_L g2744 ( 
.A(n_2537),
.Y(n_2744)
);

HB1xp67_ASAP7_75t_L g2745 ( 
.A(n_2314),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2370),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2318),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2324),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2325),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2413),
.Y(n_2750)
);

CKINVDCx20_ASAP7_75t_R g2751 ( 
.A(n_2513),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2456),
.Y(n_2752)
);

CKINVDCx5p33_ASAP7_75t_R g2753 ( 
.A(n_2386),
.Y(n_2753)
);

BUFx6f_ASAP7_75t_L g2754 ( 
.A(n_2435),
.Y(n_2754)
);

BUFx10_ASAP7_75t_L g2755 ( 
.A(n_2555),
.Y(n_2755)
);

INVx1_ASAP7_75t_SL g2756 ( 
.A(n_2252),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2414),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2497),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2299),
.B(n_1515),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2418),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2503),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2320),
.B(n_1571),
.Y(n_2762)
);

CKINVDCx5p33_ASAP7_75t_R g2763 ( 
.A(n_2393),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2349),
.B(n_1530),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2504),
.Y(n_2765)
);

CKINVDCx5p33_ASAP7_75t_R g2766 ( 
.A(n_2401),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_2310),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2505),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2331),
.B(n_2359),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2422),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2427),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2436),
.Y(n_2772)
);

CKINVDCx20_ASAP7_75t_R g2773 ( 
.A(n_2447),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2451),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2524),
.Y(n_2775)
);

HB1xp67_ASAP7_75t_L g2776 ( 
.A(n_2319),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2467),
.Y(n_2777)
);

BUFx6f_ASAP7_75t_L g2778 ( 
.A(n_2440),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2534),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2541),
.Y(n_2780)
);

CKINVDCx5p33_ASAP7_75t_R g2781 ( 
.A(n_2310),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2471),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2385),
.B(n_1530),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_SL g2784 ( 
.A(n_2284),
.B(n_2434),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2316),
.B(n_1577),
.Y(n_2785)
);

BUFx2_ASAP7_75t_L g2786 ( 
.A(n_2448),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2481),
.Y(n_2787)
);

BUFx6f_ASAP7_75t_L g2788 ( 
.A(n_2446),
.Y(n_2788)
);

CKINVDCx5p33_ASAP7_75t_R g2789 ( 
.A(n_2545),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2278),
.B(n_1577),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2548),
.Y(n_2791)
);

HB1xp67_ASAP7_75t_L g2792 ( 
.A(n_2569),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2553),
.Y(n_2793)
);

CKINVDCx5p33_ASAP7_75t_R g2794 ( 
.A(n_2327),
.Y(n_2794)
);

INVxp33_ASAP7_75t_L g2795 ( 
.A(n_2251),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2561),
.Y(n_2796)
);

HB1xp67_ASAP7_75t_L g2797 ( 
.A(n_2558),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2363),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2369),
.B(n_1722),
.Y(n_2799)
);

HB1xp67_ASAP7_75t_L g2800 ( 
.A(n_2560),
.Y(n_2800)
);

HB1xp67_ASAP7_75t_L g2801 ( 
.A(n_2280),
.Y(n_2801)
);

CKINVDCx5p33_ASAP7_75t_R g2802 ( 
.A(n_2551),
.Y(n_2802)
);

AND2x6_ASAP7_75t_L g2803 ( 
.A(n_2426),
.B(n_1868),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2486),
.Y(n_2804)
);

HB1xp67_ASAP7_75t_L g2805 ( 
.A(n_2441),
.Y(n_2805)
);

AND2x2_ASAP7_75t_L g2806 ( 
.A(n_2374),
.B(n_1632),
.Y(n_2806)
);

BUFx3_ASAP7_75t_L g2807 ( 
.A(n_2462),
.Y(n_2807)
);

CKINVDCx20_ASAP7_75t_R g2808 ( 
.A(n_2496),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2493),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2500),
.Y(n_2810)
);

BUFx6f_ASAP7_75t_L g2811 ( 
.A(n_2458),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2383),
.B(n_1632),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2371),
.Y(n_2813)
);

CKINVDCx5p33_ASAP7_75t_R g2814 ( 
.A(n_2570),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2510),
.B(n_1818),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2533),
.Y(n_2816)
);

INVx3_ASAP7_75t_L g2817 ( 
.A(n_2480),
.Y(n_2817)
);

NOR2xp33_ASAP7_75t_L g2818 ( 
.A(n_2483),
.B(n_1887),
.Y(n_2818)
);

BUFx2_ASAP7_75t_L g2819 ( 
.A(n_2510),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_SL g2820 ( 
.A(n_2301),
.B(n_1302),
.Y(n_2820)
);

CKINVDCx5p33_ASAP7_75t_R g2821 ( 
.A(n_2255),
.Y(n_2821)
);

INVx3_ASAP7_75t_L g2822 ( 
.A(n_2530),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2538),
.Y(n_2823)
);

BUFx6f_ASAP7_75t_L g2824 ( 
.A(n_2461),
.Y(n_2824)
);

CKINVDCx5p33_ASAP7_75t_R g2825 ( 
.A(n_2259),
.Y(n_2825)
);

CKINVDCx5p33_ASAP7_75t_R g2826 ( 
.A(n_2419),
.Y(n_2826)
);

AND2x4_ASAP7_75t_L g2827 ( 
.A(n_2335),
.B(n_1942),
.Y(n_2827)
);

HB1xp67_ASAP7_75t_L g2828 ( 
.A(n_2562),
.Y(n_2828)
);

NAND2xp33_ASAP7_75t_SL g2829 ( 
.A(n_2372),
.B(n_1304),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2539),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2540),
.Y(n_2831)
);

BUFx6f_ASAP7_75t_L g2832 ( 
.A(n_2472),
.Y(n_2832)
);

HB1xp67_ASAP7_75t_L g2833 ( 
.A(n_2387),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2474),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2485),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2487),
.Y(n_2836)
);

BUFx2_ASAP7_75t_L g2837 ( 
.A(n_2423),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2543),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2546),
.Y(n_2839)
);

CKINVDCx5p33_ASAP7_75t_R g2840 ( 
.A(n_2443),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2559),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2563),
.B(n_1611),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2568),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2396),
.Y(n_2844)
);

CKINVDCx8_ASAP7_75t_R g2845 ( 
.A(n_2301),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2398),
.Y(n_2846)
);

CKINVDCx5p33_ASAP7_75t_R g2847 ( 
.A(n_2399),
.Y(n_2847)
);

NOR2xp67_ASAP7_75t_L g2848 ( 
.A(n_2380),
.B(n_1890),
.Y(n_2848)
);

INVx3_ASAP7_75t_L g2849 ( 
.A(n_2329),
.Y(n_2849)
);

CKINVDCx5p33_ASAP7_75t_R g2850 ( 
.A(n_2341),
.Y(n_2850)
);

AND2x6_ASAP7_75t_L g2851 ( 
.A(n_2350),
.B(n_1895),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2352),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2508),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2509),
.Y(n_2854)
);

AND2x4_ASAP7_75t_L g2855 ( 
.A(n_2431),
.B(n_1967),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2357),
.B(n_1999),
.Y(n_2856)
);

CKINVDCx5p33_ASAP7_75t_R g2857 ( 
.A(n_2488),
.Y(n_2857)
);

BUFx6f_ASAP7_75t_L g2858 ( 
.A(n_2511),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2364),
.B(n_1274),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2491),
.B(n_1277),
.Y(n_2860)
);

OAI21x1_ASAP7_75t_L g2861 ( 
.A1(n_2536),
.A2(n_1923),
.B(n_1908),
.Y(n_2861)
);

BUFx6f_ASAP7_75t_L g2862 ( 
.A(n_2523),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2388),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2332),
.B(n_1655),
.Y(n_2864)
);

INVx3_ASAP7_75t_L g2865 ( 
.A(n_2344),
.Y(n_2865)
);

CKINVDCx5p33_ASAP7_75t_R g2866 ( 
.A(n_2501),
.Y(n_2866)
);

AND2x6_ASAP7_75t_L g2867 ( 
.A(n_2528),
.B(n_1935),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2404),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2375),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2378),
.Y(n_2870)
);

CKINVDCx20_ASAP7_75t_R g2871 ( 
.A(n_2340),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2347),
.Y(n_2872)
);

INVx3_ASAP7_75t_L g2873 ( 
.A(n_2408),
.Y(n_2873)
);

CKINVDCx5p33_ASAP7_75t_R g2874 ( 
.A(n_2535),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2351),
.Y(n_2875)
);

CKINVDCx5p33_ASAP7_75t_R g2876 ( 
.A(n_2289),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2542),
.Y(n_2877)
);

INVx3_ASAP7_75t_L g2878 ( 
.A(n_2571),
.Y(n_2878)
);

BUFx3_ASAP7_75t_L g2879 ( 
.A(n_2544),
.Y(n_2879)
);

CKINVDCx5p33_ASAP7_75t_R g2880 ( 
.A(n_2323),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2550),
.B(n_2405),
.Y(n_2881)
);

BUFx2_ASAP7_75t_L g2882 ( 
.A(n_2433),
.Y(n_2882)
);

OAI21x1_ASAP7_75t_L g2883 ( 
.A1(n_2417),
.A2(n_1952),
.B(n_1940),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2442),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2502),
.Y(n_2885)
);

CKINVDCx5p33_ASAP7_75t_R g2886 ( 
.A(n_2452),
.Y(n_2886)
);

INVx2_ASAP7_75t_SL g2887 ( 
.A(n_2577),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2582),
.Y(n_2888)
);

AOI22xp33_ASAP7_75t_L g2889 ( 
.A1(n_2851),
.A2(n_2489),
.B1(n_2499),
.B2(n_2445),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2653),
.B(n_2515),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2696),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2697),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2664),
.B(n_2519),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2699),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2870),
.B(n_2531),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2591),
.Y(n_2896)
);

BUFx2_ASAP7_75t_L g2897 ( 
.A(n_2730),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2654),
.Y(n_2898)
);

INVx3_ASAP7_75t_L g2899 ( 
.A(n_2733),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2671),
.Y(n_2900)
);

BUFx10_ASAP7_75t_L g2901 ( 
.A(n_2574),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2798),
.Y(n_2902)
);

AOI22xp33_ASAP7_75t_L g2903 ( 
.A1(n_2851),
.A2(n_2384),
.B1(n_2376),
.B2(n_2051),
.Y(n_2903)
);

AND2x2_ASAP7_75t_L g2904 ( 
.A(n_2588),
.B(n_2392),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2677),
.B(n_2818),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2813),
.Y(n_2906)
);

AO21x2_ASAP7_75t_L g2907 ( 
.A1(n_2869),
.A2(n_1973),
.B(n_1962),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2580),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_SL g2909 ( 
.A(n_2814),
.B(n_2394),
.Y(n_2909)
);

AND2x6_ASAP7_75t_L g2910 ( 
.A(n_2864),
.B(n_2806),
.Y(n_2910)
);

OR2x6_ASAP7_75t_L g2911 ( 
.A(n_2610),
.B(n_1891),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2857),
.B(n_1720),
.Y(n_2912)
);

INVx2_ASAP7_75t_SL g2913 ( 
.A(n_2619),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2866),
.B(n_1859),
.Y(n_2914)
);

INVx4_ASAP7_75t_L g2915 ( 
.A(n_2702),
.Y(n_2915)
);

OR2x6_ASAP7_75t_L g2916 ( 
.A(n_2683),
.B(n_1320),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2585),
.Y(n_2917)
);

INVx5_ASAP7_75t_L g2918 ( 
.A(n_2663),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2874),
.B(n_1859),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2586),
.Y(n_2920)
);

NOR2xp33_ASAP7_75t_L g2921 ( 
.A(n_2850),
.B(n_2028),
.Y(n_2921)
);

BUFx6f_ASAP7_75t_SL g2922 ( 
.A(n_2728),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2676),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2704),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2679),
.Y(n_2925)
);

HB1xp67_ASAP7_75t_L g2926 ( 
.A(n_2641),
.Y(n_2926)
);

INVx2_ASAP7_75t_SL g2927 ( 
.A(n_2663),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2705),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2622),
.B(n_1655),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2706),
.Y(n_2930)
);

INVxp33_ASAP7_75t_L g2931 ( 
.A(n_2659),
.Y(n_2931)
);

BUFx3_ASAP7_75t_L g2932 ( 
.A(n_2604),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2709),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2713),
.Y(n_2934)
);

BUFx6f_ASAP7_75t_SL g2935 ( 
.A(n_2674),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2714),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2688),
.Y(n_2937)
);

INVx3_ASAP7_75t_L g2938 ( 
.A(n_2716),
.Y(n_2938)
);

NOR2xp33_ASAP7_75t_SL g2939 ( 
.A(n_2609),
.B(n_1661),
.Y(n_2939)
);

AND2x4_ASAP7_75t_L g2940 ( 
.A(n_2634),
.B(n_2626),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2599),
.B(n_1859),
.Y(n_2941)
);

INVx3_ASAP7_75t_L g2942 ( 
.A(n_2620),
.Y(n_2942)
);

NAND2xp33_ASAP7_75t_L g2943 ( 
.A(n_2611),
.B(n_1309),
.Y(n_2943)
);

CKINVDCx5p33_ASAP7_75t_R g2944 ( 
.A(n_2614),
.Y(n_2944)
);

AOI21x1_ASAP7_75t_L g2945 ( 
.A1(n_2651),
.A2(n_2039),
.B(n_2037),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2692),
.Y(n_2946)
);

OR2x2_ASAP7_75t_L g2947 ( 
.A(n_2693),
.B(n_1656),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2701),
.Y(n_2948)
);

INVx4_ASAP7_75t_L g2949 ( 
.A(n_2644),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2731),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2718),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2721),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2732),
.Y(n_2953)
);

INVx3_ASAP7_75t_L g2954 ( 
.A(n_2620),
.Y(n_2954)
);

NAND3xp33_ASAP7_75t_L g2955 ( 
.A(n_2649),
.B(n_1313),
.C(n_1312),
.Y(n_2955)
);

NOR2xp33_ASAP7_75t_L g2956 ( 
.A(n_2665),
.B(n_1317),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2741),
.Y(n_2957)
);

AND2x6_ASAP7_75t_L g2958 ( 
.A(n_2675),
.B(n_2053),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2867),
.B(n_1930),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2752),
.Y(n_2960)
);

AND3x2_ASAP7_75t_L g2961 ( 
.A(n_2735),
.B(n_1378),
.C(n_1364),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2758),
.Y(n_2962)
);

INVx1_ASAP7_75t_SL g2963 ( 
.A(n_2680),
.Y(n_2963)
);

INVx4_ASAP7_75t_L g2964 ( 
.A(n_2648),
.Y(n_2964)
);

BUFx6f_ASAP7_75t_L g2965 ( 
.A(n_2640),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2867),
.B(n_1930),
.Y(n_2966)
);

INVx3_ASAP7_75t_L g2967 ( 
.A(n_2666),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2722),
.B(n_1325),
.Y(n_2968)
);

AOI21x1_ASAP7_75t_L g2969 ( 
.A1(n_2872),
.A2(n_2884),
.B(n_2875),
.Y(n_2969)
);

INVxp33_ASAP7_75t_L g2970 ( 
.A(n_2711),
.Y(n_2970)
);

CKINVDCx5p33_ASAP7_75t_R g2971 ( 
.A(n_2618),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2761),
.Y(n_2972)
);

INVx2_ASAP7_75t_SL g2973 ( 
.A(n_2755),
.Y(n_2973)
);

INVx1_ASAP7_75t_SL g2974 ( 
.A(n_2681),
.Y(n_2974)
);

INVx4_ASAP7_75t_L g2975 ( 
.A(n_2661),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_SL g2976 ( 
.A(n_2789),
.B(n_1326),
.Y(n_2976)
);

INVx3_ASAP7_75t_L g2977 ( 
.A(n_2685),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2734),
.Y(n_2978)
);

NAND2xp33_ASAP7_75t_L g2979 ( 
.A(n_2623),
.B(n_1329),
.Y(n_2979)
);

CKINVDCx20_ASAP7_75t_R g2980 ( 
.A(n_2632),
.Y(n_2980)
);

OR2x2_ASAP7_75t_L g2981 ( 
.A(n_2684),
.B(n_1657),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2765),
.Y(n_2982)
);

NAND3xp33_ASAP7_75t_L g2983 ( 
.A(n_2633),
.B(n_1350),
.C(n_1336),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2867),
.B(n_1930),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_SL g2985 ( 
.A(n_2786),
.B(n_1351),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2742),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_SL g2987 ( 
.A(n_2827),
.B(n_1352),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_SL g2988 ( 
.A(n_2630),
.B(n_1354),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2860),
.B(n_2032),
.Y(n_2989)
);

CKINVDCx5p33_ASAP7_75t_R g2990 ( 
.A(n_2631),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2647),
.B(n_2581),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2747),
.Y(n_2992)
);

INVxp67_ASAP7_75t_R g2993 ( 
.A(n_2743),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2748),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2749),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2768),
.Y(n_2996)
);

INVx5_ASAP7_75t_L g2997 ( 
.A(n_2803),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2775),
.Y(n_2998)
);

AOI22xp33_ASAP7_75t_SL g2999 ( 
.A1(n_2703),
.A2(n_1806),
.B1(n_1929),
.B2(n_1661),
.Y(n_2999)
);

INVx8_ASAP7_75t_L g3000 ( 
.A(n_2737),
.Y(n_3000)
);

NAND2xp33_ASAP7_75t_L g3001 ( 
.A(n_2639),
.B(n_1360),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2779),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2668),
.B(n_2672),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2750),
.Y(n_3004)
);

INVx3_ASAP7_75t_L g3005 ( 
.A(n_2715),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2678),
.B(n_2032),
.Y(n_3006)
);

OAI21xp33_ASAP7_75t_SL g3007 ( 
.A1(n_2687),
.A2(n_2694),
.B(n_2657),
.Y(n_3007)
);

AOI22xp33_ASAP7_75t_L g3008 ( 
.A1(n_2851),
.A2(n_1429),
.B1(n_1484),
.B2(n_1394),
.Y(n_3008)
);

INVx3_ASAP7_75t_L g3009 ( 
.A(n_2739),
.Y(n_3009)
);

NOR2x1p5_ASAP7_75t_L g3010 ( 
.A(n_2601),
.B(n_1363),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2757),
.B(n_2760),
.Y(n_3011)
);

AOI22xp33_ASAP7_75t_L g3012 ( 
.A1(n_2790),
.A2(n_1553),
.B1(n_1588),
.B2(n_1510),
.Y(n_3012)
);

BUFx6f_ASAP7_75t_L g3013 ( 
.A(n_2640),
.Y(n_3013)
);

BUFx3_ASAP7_75t_L g3014 ( 
.A(n_2662),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2780),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2770),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2771),
.B(n_2032),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2772),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2774),
.B(n_2777),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2782),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2791),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2793),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2796),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2576),
.Y(n_3024)
);

INVx3_ASAP7_75t_L g3025 ( 
.A(n_2646),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2787),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2804),
.B(n_2809),
.Y(n_3027)
);

INVx3_ASAP7_75t_L g3028 ( 
.A(n_2646),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2579),
.Y(n_3029)
);

INVx3_ASAP7_75t_L g3030 ( 
.A(n_2673),
.Y(n_3030)
);

BUFx6f_ASAP7_75t_SL g3031 ( 
.A(n_2695),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2810),
.Y(n_3032)
);

INVx3_ASAP7_75t_L g3033 ( 
.A(n_2673),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2656),
.Y(n_3034)
);

INVx2_ASAP7_75t_SL g3035 ( 
.A(n_2720),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2660),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2667),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2816),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2823),
.B(n_2830),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2831),
.B(n_1366),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2838),
.B(n_1369),
.Y(n_3041)
);

BUFx10_ASAP7_75t_L g3042 ( 
.A(n_2575),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2839),
.B(n_1370),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2868),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_L g3045 ( 
.A(n_2756),
.B(n_1371),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_L g3046 ( 
.A(n_2587),
.B(n_1372),
.Y(n_3046)
);

NOR2xp33_ASAP7_75t_L g3047 ( 
.A(n_2596),
.B(n_2886),
.Y(n_3047)
);

AOI22xp33_ASAP7_75t_SL g3048 ( 
.A1(n_2669),
.A2(n_1929),
.B1(n_1945),
.B2(n_1806),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2841),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2736),
.B(n_1373),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2843),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_SL g3052 ( 
.A(n_2686),
.B(n_1376),
.Y(n_3052)
);

BUFx6f_ASAP7_75t_L g3053 ( 
.A(n_2708),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_2876),
.B(n_1377),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2769),
.Y(n_3055)
);

BUFx2_ASAP7_75t_L g3056 ( 
.A(n_2719),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2885),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_SL g3058 ( 
.A(n_2689),
.B(n_2690),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2852),
.Y(n_3059)
);

INVx2_ASAP7_75t_L g3060 ( 
.A(n_2607),
.Y(n_3060)
);

NOR2xp33_ASAP7_75t_L g3061 ( 
.A(n_2880),
.B(n_1380),
.Y(n_3061)
);

OAI22xp5_ASAP7_75t_L g3062 ( 
.A1(n_2863),
.A2(n_1383),
.B1(n_1391),
.B2(n_1382),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2707),
.Y(n_3063)
);

INVxp67_ASAP7_75t_SL g3064 ( 
.A(n_2833),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2844),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2846),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2849),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2859),
.B(n_1392),
.Y(n_3068)
);

CKINVDCx20_ASAP7_75t_R g3069 ( 
.A(n_2642),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2865),
.Y(n_3070)
);

INVx1_ASAP7_75t_SL g3071 ( 
.A(n_2691),
.Y(n_3071)
);

INVx1_ASAP7_75t_SL g3072 ( 
.A(n_2615),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2817),
.Y(n_3073)
);

NAND2xp33_ASAP7_75t_SL g3074 ( 
.A(n_2767),
.B(n_1396),
.Y(n_3074)
);

AND2x2_ASAP7_75t_L g3075 ( 
.A(n_2624),
.B(n_1945),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_SL g3076 ( 
.A(n_2781),
.B(n_1398),
.Y(n_3076)
);

NOR2xp33_ASAP7_75t_R g3077 ( 
.A(n_2670),
.B(n_1280),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2822),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2883),
.Y(n_3079)
);

INVx2_ASAP7_75t_SL g3080 ( 
.A(n_2812),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2594),
.Y(n_3081)
);

INVx3_ASAP7_75t_L g3082 ( 
.A(n_2708),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2801),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2612),
.Y(n_3084)
);

BUFx3_ASAP7_75t_L g3085 ( 
.A(n_2578),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2621),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2805),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2602),
.B(n_1400),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2828),
.Y(n_3089)
);

BUFx2_ASAP7_75t_L g3090 ( 
.A(n_2797),
.Y(n_3090)
);

AOI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_2638),
.A2(n_2061),
.B1(n_2064),
.B2(n_2060),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_2625),
.Y(n_3092)
);

NAND2xp33_ASAP7_75t_SL g3093 ( 
.A(n_2729),
.B(n_2635),
.Y(n_3093)
);

AND2x2_ASAP7_75t_L g3094 ( 
.A(n_2764),
.B(n_1970),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2698),
.B(n_1401),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_SL g3096 ( 
.A(n_2819),
.B(n_1403),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2842),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2807),
.Y(n_3098)
);

OR2x6_ASAP7_75t_L g3099 ( 
.A(n_2800),
.B(n_1629),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2759),
.Y(n_3100)
);

NAND2xp33_ASAP7_75t_L g3101 ( 
.A(n_2637),
.B(n_1406),
.Y(n_3101)
);

AO22x2_ASAP7_75t_L g3102 ( 
.A1(n_2773),
.A2(n_1658),
.B1(n_1668),
.B2(n_1662),
.Y(n_3102)
);

NAND3xp33_ASAP7_75t_L g3103 ( 
.A(n_2613),
.B(n_2783),
.C(n_2700),
.Y(n_3103)
);

NAND2xp33_ASAP7_75t_R g3104 ( 
.A(n_2746),
.B(n_1408),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2628),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2762),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2834),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2799),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2835),
.Y(n_3109)
);

NOR2xp33_ASAP7_75t_L g3110 ( 
.A(n_2784),
.B(n_1410),
.Y(n_3110)
);

INVx5_ASAP7_75t_L g3111 ( 
.A(n_2803),
.Y(n_3111)
);

AOI22xp33_ASAP7_75t_L g3112 ( 
.A1(n_2637),
.A2(n_1671),
.B1(n_1703),
.B2(n_1654),
.Y(n_3112)
);

INVx2_ASAP7_75t_SL g3113 ( 
.A(n_2785),
.Y(n_3113)
);

NAND3xp33_ASAP7_75t_L g3114 ( 
.A(n_2829),
.B(n_1415),
.C(n_1414),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2589),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2836),
.Y(n_3116)
);

CKINVDCx6p67_ASAP7_75t_R g3117 ( 
.A(n_2629),
.Y(n_3117)
);

INVx1_ASAP7_75t_SL g3118 ( 
.A(n_2837),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2597),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2853),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2854),
.Y(n_3121)
);

OR2x2_ASAP7_75t_L g3122 ( 
.A(n_2882),
.B(n_1675),
.Y(n_3122)
);

NAND3xp33_ASAP7_75t_L g3123 ( 
.A(n_2717),
.B(n_1420),
.C(n_1417),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_2877),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2603),
.Y(n_3125)
);

INVx3_ASAP7_75t_L g3126 ( 
.A(n_2723),
.Y(n_3126)
);

NOR2xp33_ASAP7_75t_L g3127 ( 
.A(n_2745),
.B(n_1421),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_2583),
.Y(n_3128)
);

NOR2xp33_ASAP7_75t_L g3129 ( 
.A(n_2921),
.B(n_2751),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2905),
.B(n_2637),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_SL g3131 ( 
.A(n_2963),
.B(n_2744),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2888),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_2893),
.B(n_2815),
.Y(n_3133)
);

OR2x6_ASAP7_75t_L g3134 ( 
.A(n_3000),
.B(n_2776),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2891),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_3100),
.B(n_2856),
.Y(n_3136)
);

NOR2xp33_ASAP7_75t_L g3137 ( 
.A(n_3047),
.B(n_2808),
.Y(n_3137)
);

INVx3_ASAP7_75t_L g3138 ( 
.A(n_2915),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_3106),
.B(n_2803),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_3108),
.B(n_2855),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_2974),
.B(n_2845),
.Y(n_3141)
);

NOR2xp33_ASAP7_75t_L g3142 ( 
.A(n_3071),
.B(n_2753),
.Y(n_3142)
);

INVx2_ASAP7_75t_SL g3143 ( 
.A(n_2887),
.Y(n_3143)
);

INVxp67_ASAP7_75t_L g3144 ( 
.A(n_2897),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_SL g3145 ( 
.A(n_2944),
.B(n_2710),
.Y(n_3145)
);

NOR3xp33_ASAP7_75t_L g3146 ( 
.A(n_3058),
.B(n_2738),
.C(n_2820),
.Y(n_3146)
);

NOR2xp33_ASAP7_75t_L g3147 ( 
.A(n_2970),
.B(n_2763),
.Y(n_3147)
);

CKINVDCx20_ASAP7_75t_R g3148 ( 
.A(n_3069),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_2896),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2898),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_3097),
.B(n_2792),
.Y(n_3151)
);

NAND3xp33_ASAP7_75t_L g3152 ( 
.A(n_2968),
.B(n_2990),
.C(n_2971),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2892),
.Y(n_3153)
);

NOR2xp67_ASAP7_75t_L g3154 ( 
.A(n_2918),
.B(n_2712),
.Y(n_3154)
);

NOR2xp67_ASAP7_75t_L g3155 ( 
.A(n_2918),
.B(n_2724),
.Y(n_3155)
);

NOR2xp67_ASAP7_75t_L g3156 ( 
.A(n_2949),
.B(n_2725),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2894),
.Y(n_3157)
);

NAND3xp33_ASAP7_75t_L g3158 ( 
.A(n_2943),
.B(n_2592),
.C(n_2590),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_3046),
.B(n_2881),
.Y(n_3159)
);

AND2x4_ASAP7_75t_L g3160 ( 
.A(n_2932),
.B(n_2766),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2924),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_3055),
.B(n_3088),
.Y(n_3162)
);

NAND2xp33_ASAP7_75t_L g3163 ( 
.A(n_2910),
.B(n_2593),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2928),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2930),
.B(n_2873),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_SL g3166 ( 
.A(n_2997),
.B(n_2878),
.Y(n_3166)
);

HB1xp67_ASAP7_75t_L g3167 ( 
.A(n_2926),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2900),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_SL g3169 ( 
.A(n_2997),
.B(n_2584),
.Y(n_3169)
);

NOR2xp67_ASAP7_75t_L g3170 ( 
.A(n_2964),
.B(n_2595),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_3111),
.B(n_2627),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2902),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2933),
.B(n_2605),
.Y(n_3173)
);

INVxp33_ASAP7_75t_L g3174 ( 
.A(n_2940),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2934),
.B(n_2606),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2936),
.Y(n_3176)
);

INVx2_ASAP7_75t_SL g3177 ( 
.A(n_2913),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2950),
.Y(n_3178)
);

NOR2xp33_ASAP7_75t_L g3179 ( 
.A(n_2931),
.B(n_2795),
.Y(n_3179)
);

NAND2xp33_ASAP7_75t_L g3180 ( 
.A(n_2910),
.B(n_2598),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_SL g3181 ( 
.A(n_3111),
.B(n_2848),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2906),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_SL g3183 ( 
.A(n_3103),
.B(n_2608),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2978),
.Y(n_3184)
);

BUFx6f_ASAP7_75t_L g3185 ( 
.A(n_2965),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2908),
.Y(n_3186)
);

BUFx2_ASAP7_75t_L g3187 ( 
.A(n_3056),
.Y(n_3187)
);

NOR2xp33_ASAP7_75t_L g3188 ( 
.A(n_3072),
.B(n_2616),
.Y(n_3188)
);

NOR2xp33_ASAP7_75t_L g3189 ( 
.A(n_3118),
.B(n_2617),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2986),
.B(n_2636),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2992),
.Y(n_3191)
);

AO221x1_ASAP7_75t_L g3192 ( 
.A1(n_3102),
.A2(n_2727),
.B1(n_2754),
.B2(n_2726),
.C(n_2723),
.Y(n_3192)
);

INVx2_ASAP7_75t_L g3193 ( 
.A(n_2917),
.Y(n_3193)
);

NAND2xp33_ASAP7_75t_L g3194 ( 
.A(n_2910),
.B(n_2600),
.Y(n_3194)
);

OAI21xp5_ASAP7_75t_L g3195 ( 
.A1(n_3007),
.A2(n_2861),
.B(n_1682),
.Y(n_3195)
);

NAND2xp33_ASAP7_75t_L g3196 ( 
.A(n_3068),
.B(n_1423),
.Y(n_3196)
);

AOI22xp33_ASAP7_75t_L g3197 ( 
.A1(n_2958),
.A2(n_2645),
.B1(n_2650),
.B2(n_2643),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2920),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_SL g3199 ( 
.A(n_3113),
.B(n_2652),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2994),
.B(n_2655),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2995),
.B(n_1680),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2923),
.Y(n_3202)
);

BUFx5_ASAP7_75t_L g3203 ( 
.A(n_3004),
.Y(n_3203)
);

INVx2_ASAP7_75t_SL g3204 ( 
.A(n_3000),
.Y(n_3204)
);

INVxp67_ASAP7_75t_L g3205 ( 
.A(n_3090),
.Y(n_3205)
);

INVx4_ASAP7_75t_L g3206 ( 
.A(n_2899),
.Y(n_3206)
);

INVx3_ASAP7_75t_L g3207 ( 
.A(n_3014),
.Y(n_3207)
);

BUFx6f_ASAP7_75t_SL g3208 ( 
.A(n_3085),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_2925),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_L g3210 ( 
.A(n_3054),
.B(n_2740),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_3016),
.B(n_1683),
.Y(n_3211)
);

INVx1_ASAP7_75t_SL g3212 ( 
.A(n_2980),
.Y(n_3212)
);

AND2x2_ASAP7_75t_L g3213 ( 
.A(n_3094),
.B(n_2879),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3018),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_SL g3215 ( 
.A(n_3080),
.B(n_1430),
.Y(n_3215)
);

OR2x2_ASAP7_75t_L g3216 ( 
.A(n_2947),
.B(n_2726),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_2937),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_3020),
.B(n_1686),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_3026),
.B(n_3032),
.Y(n_3219)
);

NOR2xp33_ASAP7_75t_L g3220 ( 
.A(n_3061),
.B(n_2871),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_SL g3221 ( 
.A(n_2939),
.B(n_1431),
.Y(n_3221)
);

INVx2_ASAP7_75t_SL g3222 ( 
.A(n_2965),
.Y(n_3222)
);

BUFx8_ASAP7_75t_L g3223 ( 
.A(n_2922),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2946),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3038),
.Y(n_3225)
);

AOI22xp33_ASAP7_75t_L g3226 ( 
.A1(n_2958),
.A2(n_2052),
.B1(n_2056),
.B2(n_1970),
.Y(n_3226)
);

NOR3xp33_ASAP7_75t_L g3227 ( 
.A(n_3001),
.B(n_1701),
.C(n_1687),
.Y(n_3227)
);

AND2x6_ASAP7_75t_L g3228 ( 
.A(n_3049),
.B(n_1331),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_SL g3229 ( 
.A(n_2991),
.B(n_1433),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_2948),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3051),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_3011),
.B(n_1714),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_SL g3233 ( 
.A(n_3019),
.B(n_1434),
.Y(n_3233)
);

BUFx3_ASAP7_75t_L g3234 ( 
.A(n_2901),
.Y(n_3234)
);

AND2x2_ASAP7_75t_SL g3235 ( 
.A(n_3101),
.B(n_2658),
.Y(n_3235)
);

NOR3xp33_ASAP7_75t_L g3236 ( 
.A(n_2979),
.B(n_1735),
.C(n_1719),
.Y(n_3236)
);

INVx8_ASAP7_75t_L g3237 ( 
.A(n_2911),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_3027),
.B(n_1736),
.Y(n_3238)
);

NOR2xp33_ASAP7_75t_L g3239 ( 
.A(n_2890),
.B(n_2682),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_3045),
.B(n_2727),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_3075),
.B(n_2895),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3024),
.Y(n_3242)
);

NOR2xp33_ASAP7_75t_L g3243 ( 
.A(n_2981),
.B(n_2754),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3039),
.B(n_1740),
.Y(n_3244)
);

INVx2_ASAP7_75t_SL g3245 ( 
.A(n_3013),
.Y(n_3245)
);

INVx2_ASAP7_75t_L g3246 ( 
.A(n_2951),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_SL g3247 ( 
.A(n_2912),
.B(n_1435),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_3029),
.B(n_1743),
.Y(n_3248)
);

NAND2xp33_ASAP7_75t_L g3249 ( 
.A(n_3003),
.B(n_1438),
.Y(n_3249)
);

NAND3xp33_ASAP7_75t_L g3250 ( 
.A(n_3050),
.B(n_2956),
.C(n_3127),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_SL g3251 ( 
.A(n_2914),
.B(n_2919),
.Y(n_3251)
);

BUFx6f_ASAP7_75t_L g3252 ( 
.A(n_3013),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3034),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_3036),
.B(n_1752),
.Y(n_3254)
);

NAND2xp33_ASAP7_75t_L g3255 ( 
.A(n_3093),
.B(n_1440),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3037),
.Y(n_3256)
);

NOR3xp33_ASAP7_75t_L g3257 ( 
.A(n_3123),
.B(n_1762),
.C(n_1753),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3059),
.B(n_1765),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_2958),
.B(n_1766),
.Y(n_3259)
);

AO221x1_ASAP7_75t_L g3260 ( 
.A1(n_3062),
.A2(n_2811),
.B1(n_2824),
.B2(n_2788),
.C(n_2778),
.Y(n_3260)
);

AO221x1_ASAP7_75t_L g3261 ( 
.A1(n_2999),
.A2(n_2811),
.B1(n_2824),
.B2(n_2788),
.C(n_2778),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_2952),
.Y(n_3262)
);

NAND2xp33_ASAP7_75t_L g3263 ( 
.A(n_2989),
.B(n_1456),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2953),
.Y(n_3264)
);

NOR2xp33_ASAP7_75t_L g3265 ( 
.A(n_3064),
.B(n_3035),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3065),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3066),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_2957),
.Y(n_3268)
);

NOR2xp67_ASAP7_75t_L g3269 ( 
.A(n_2975),
.B(n_2832),
.Y(n_3269)
);

INVxp67_ASAP7_75t_L g3270 ( 
.A(n_2904),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_SL g3271 ( 
.A(n_2967),
.B(n_1458),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_SL g3272 ( 
.A(n_2977),
.B(n_1462),
.Y(n_3272)
);

NOR2xp33_ASAP7_75t_L g3273 ( 
.A(n_3083),
.B(n_2832),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3044),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3095),
.B(n_1767),
.Y(n_3275)
);

OR2x2_ASAP7_75t_L g3276 ( 
.A(n_3122),
.B(n_2858),
.Y(n_3276)
);

NAND3xp33_ASAP7_75t_L g3277 ( 
.A(n_3110),
.B(n_1478),
.C(n_1468),
.Y(n_3277)
);

CKINVDCx5p33_ASAP7_75t_R g3278 ( 
.A(n_3117),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3017),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_2960),
.Y(n_3280)
);

OR2x6_ASAP7_75t_L g3281 ( 
.A(n_2927),
.B(n_2858),
.Y(n_3281)
);

NOR3xp33_ASAP7_75t_L g3282 ( 
.A(n_3114),
.B(n_1771),
.C(n_1770),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_2941),
.B(n_1773),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3091),
.B(n_1775),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3057),
.Y(n_3285)
);

NOR2xp33_ASAP7_75t_L g3286 ( 
.A(n_3087),
.B(n_3089),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2962),
.Y(n_3287)
);

INVxp67_ASAP7_75t_L g3288 ( 
.A(n_2929),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_SL g3289 ( 
.A(n_3005),
.B(n_1482),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3135),
.Y(n_3290)
);

NAND2x1p5_ASAP7_75t_L g3291 ( 
.A(n_3207),
.B(n_3009),
.Y(n_3291)
);

NAND2x1p5_ASAP7_75t_L g3292 ( 
.A(n_3212),
.B(n_2973),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3153),
.Y(n_3293)
);

NAND3xp33_ASAP7_75t_SL g3294 ( 
.A(n_3250),
.B(n_3077),
.C(n_3048),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3157),
.Y(n_3295)
);

AND2x2_ASAP7_75t_L g3296 ( 
.A(n_3137),
.B(n_2916),
.Y(n_3296)
);

INVx2_ASAP7_75t_SL g3297 ( 
.A(n_3237),
.Y(n_3297)
);

AO22x2_ASAP7_75t_L g3298 ( 
.A1(n_3242),
.A2(n_2983),
.B1(n_3119),
.B2(n_3115),
.Y(n_3298)
);

CKINVDCx5p33_ASAP7_75t_R g3299 ( 
.A(n_3148),
.Y(n_3299)
);

NAND2x1p5_ASAP7_75t_L g3300 ( 
.A(n_3185),
.B(n_3053),
.Y(n_3300)
);

AND2x2_ASAP7_75t_L g3301 ( 
.A(n_3129),
.B(n_2916),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3161),
.Y(n_3302)
);

BUFx8_ASAP7_75t_L g3303 ( 
.A(n_3208),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3164),
.Y(n_3304)
);

AO22x2_ASAP7_75t_L g3305 ( 
.A1(n_3253),
.A2(n_3125),
.B1(n_2987),
.B2(n_3084),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3176),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3241),
.B(n_3012),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_SL g3308 ( 
.A(n_3152),
.B(n_2889),
.Y(n_3308)
);

OAI221xp5_ASAP7_75t_L g3309 ( 
.A1(n_3288),
.A2(n_2903),
.B1(n_2985),
.B2(n_3052),
.C(n_3112),
.Y(n_3309)
);

INVxp67_ASAP7_75t_L g3310 ( 
.A(n_3167),
.Y(n_3310)
);

OAI221xp5_ASAP7_75t_L g3311 ( 
.A1(n_3226),
.A2(n_3227),
.B1(n_3236),
.B2(n_3210),
.C(n_3142),
.Y(n_3311)
);

AO22x2_ASAP7_75t_L g3312 ( 
.A1(n_3256),
.A2(n_3086),
.B1(n_3092),
.B2(n_3081),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3178),
.Y(n_3313)
);

BUFx8_ASAP7_75t_L g3314 ( 
.A(n_3187),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3184),
.Y(n_3315)
);

NOR2xp33_ASAP7_75t_L g3316 ( 
.A(n_3144),
.B(n_2988),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3191),
.Y(n_3317)
);

INVx3_ASAP7_75t_L g3318 ( 
.A(n_3185),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_3186),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3214),
.Y(n_3320)
);

NAND2x1p5_ASAP7_75t_L g3321 ( 
.A(n_3252),
.B(n_3053),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3225),
.Y(n_3322)
);

NAND2x1p5_ASAP7_75t_L g3323 ( 
.A(n_3252),
.B(n_2942),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_3133),
.B(n_3008),
.Y(n_3324)
);

AND2x4_ASAP7_75t_L g3325 ( 
.A(n_3134),
.B(n_3160),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3231),
.Y(n_3326)
);

NAND2x1p5_ASAP7_75t_L g3327 ( 
.A(n_3234),
.B(n_2954),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_3193),
.Y(n_3328)
);

NAND2x1p5_ASAP7_75t_L g3329 ( 
.A(n_3143),
.B(n_2938),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_3266),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3267),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3219),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3198),
.Y(n_3333)
);

AO22x2_ASAP7_75t_L g3334 ( 
.A1(n_3274),
.A2(n_3105),
.B1(n_3109),
.B2(n_3107),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3285),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3173),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3175),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_3132),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3190),
.Y(n_3339)
);

AOI22xp5_ASAP7_75t_L g3340 ( 
.A1(n_3220),
.A2(n_3104),
.B1(n_3074),
.B2(n_2935),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3162),
.B(n_3040),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3200),
.Y(n_3342)
);

AND2x4_ASAP7_75t_L g3343 ( 
.A(n_3134),
.B(n_3025),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3287),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3149),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_3150),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3168),
.Y(n_3347)
);

OAI221xp5_ASAP7_75t_L g3348 ( 
.A1(n_3205),
.A2(n_3043),
.B1(n_3041),
.B2(n_2976),
.C(n_2955),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_3172),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3182),
.Y(n_3350)
);

AO22x2_ASAP7_75t_L g3351 ( 
.A1(n_3192),
.A2(n_3120),
.B1(n_3121),
.B2(n_3116),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3202),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3209),
.Y(n_3353)
);

NAND2x1p5_ASAP7_75t_L g3354 ( 
.A(n_3206),
.B(n_3028),
.Y(n_3354)
);

BUFx6f_ASAP7_75t_L g3355 ( 
.A(n_3237),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3217),
.Y(n_3356)
);

AO22x2_ASAP7_75t_L g3357 ( 
.A1(n_3259),
.A2(n_3124),
.B1(n_3096),
.B2(n_3098),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_3224),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3230),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3246),
.Y(n_3360)
);

AND2x2_ASAP7_75t_L g3361 ( 
.A(n_3213),
.B(n_3099),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3262),
.Y(n_3362)
);

AO22x2_ASAP7_75t_L g3363 ( 
.A1(n_3130),
.A2(n_3076),
.B1(n_2961),
.B2(n_3070),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3159),
.B(n_3067),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3264),
.Y(n_3365)
);

BUFx8_ASAP7_75t_L g3366 ( 
.A(n_3204),
.Y(n_3366)
);

NOR2xp33_ASAP7_75t_L g3367 ( 
.A(n_3174),
.B(n_3099),
.Y(n_3367)
);

NAND2x1p5_ASAP7_75t_L g3368 ( 
.A(n_3222),
.B(n_3030),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3136),
.B(n_3073),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3268),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3280),
.Y(n_3371)
);

BUFx6f_ASAP7_75t_SL g3372 ( 
.A(n_3177),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3248),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3243),
.B(n_2993),
.Y(n_3374)
);

OAI221xp5_ASAP7_75t_L g3375 ( 
.A1(n_3221),
.A2(n_2911),
.B1(n_3078),
.B2(n_2909),
.C(n_3033),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3254),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3201),
.Y(n_3377)
);

INVx2_ASAP7_75t_L g3378 ( 
.A(n_3203),
.Y(n_3378)
);

AO22x2_ASAP7_75t_L g3379 ( 
.A1(n_3216),
.A2(n_3183),
.B1(n_3140),
.B2(n_3276),
.Y(n_3379)
);

AO22x2_ASAP7_75t_L g3380 ( 
.A1(n_3139),
.A2(n_2982),
.B1(n_2996),
.B2(n_2972),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3211),
.Y(n_3381)
);

AO22x2_ASAP7_75t_L g3382 ( 
.A1(n_3229),
.A2(n_3002),
.B1(n_3015),
.B2(n_2998),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_3203),
.Y(n_3383)
);

AO22x2_ASAP7_75t_L g3384 ( 
.A1(n_3284),
.A2(n_3022),
.B1(n_3023),
.B2(n_3021),
.Y(n_3384)
);

AND2x2_ASAP7_75t_L g3385 ( 
.A(n_3286),
.B(n_3082),
.Y(n_3385)
);

AND2x6_ASAP7_75t_L g3386 ( 
.A(n_3138),
.B(n_3126),
.Y(n_3386)
);

BUFx3_ASAP7_75t_L g3387 ( 
.A(n_3223),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3218),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3258),
.Y(n_3389)
);

NAND2x1p5_ASAP7_75t_L g3390 ( 
.A(n_3245),
.B(n_3010),
.Y(n_3390)
);

AO22x2_ASAP7_75t_L g3391 ( 
.A1(n_3270),
.A2(n_2959),
.B1(n_2984),
.B2(n_2966),
.Y(n_3391)
);

HB1xp67_ASAP7_75t_L g3392 ( 
.A(n_3281),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3151),
.Y(n_3393)
);

INVx2_ASAP7_75t_SL g3394 ( 
.A(n_3281),
.Y(n_3394)
);

AND2x4_ASAP7_75t_L g3395 ( 
.A(n_3269),
.B(n_2862),
.Y(n_3395)
);

AND2x4_ASAP7_75t_L g3396 ( 
.A(n_3170),
.B(n_2862),
.Y(n_3396)
);

INVxp67_ASAP7_75t_L g3397 ( 
.A(n_3189),
.Y(n_3397)
);

NAND2x1p5_ASAP7_75t_L g3398 ( 
.A(n_3154),
.B(n_3042),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3165),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_3283),
.Y(n_3400)
);

NAND2x1p5_ASAP7_75t_L g3401 ( 
.A(n_3155),
.B(n_3031),
.Y(n_3401)
);

NAND2x1p5_ASAP7_75t_L g3402 ( 
.A(n_3145),
.B(n_2969),
.Y(n_3402)
);

AO22x2_ASAP7_75t_L g3403 ( 
.A1(n_3233),
.A2(n_3060),
.B1(n_3063),
.B2(n_3128),
.Y(n_3403)
);

BUFx6f_ASAP7_75t_L g3404 ( 
.A(n_3278),
.Y(n_3404)
);

BUFx8_ASAP7_75t_L g3405 ( 
.A(n_3228),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3232),
.Y(n_3406)
);

AOI22xp5_ASAP7_75t_L g3407 ( 
.A1(n_3179),
.A2(n_2802),
.B1(n_3006),
.B2(n_1489),
.Y(n_3407)
);

AND2x2_ASAP7_75t_SL g3408 ( 
.A(n_3235),
.B(n_1706),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3240),
.B(n_2907),
.Y(n_3409)
);

NAND2xp33_ASAP7_75t_L g3410 ( 
.A(n_3203),
.B(n_3079),
.Y(n_3410)
);

AND2x6_ASAP7_75t_SL g3411 ( 
.A(n_3147),
.B(n_1790),
.Y(n_3411)
);

AO22x2_ASAP7_75t_L g3412 ( 
.A1(n_3257),
.A2(n_3277),
.B1(n_3215),
.B2(n_3199),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_3265),
.B(n_2052),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_3203),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3238),
.Y(n_3415)
);

NAND2x1p5_ASAP7_75t_L g3416 ( 
.A(n_3156),
.B(n_2547),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3244),
.Y(n_3417)
);

CKINVDCx20_ASAP7_75t_R g3418 ( 
.A(n_3158),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3275),
.B(n_1483),
.Y(n_3419)
);

NAND2x1p5_ASAP7_75t_L g3420 ( 
.A(n_3141),
.B(n_2554),
.Y(n_3420)
);

AO22x2_ASAP7_75t_L g3421 ( 
.A1(n_3279),
.A2(n_2794),
.B1(n_2847),
.B2(n_1803),
.Y(n_3421)
);

NAND2x1p5_ASAP7_75t_L g3422 ( 
.A(n_3169),
.B(n_2945),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3260),
.Y(n_3423)
);

AOI21xp5_ASAP7_75t_L g3424 ( 
.A1(n_3410),
.A2(n_3251),
.B(n_3196),
.Y(n_3424)
);

NOR2xp33_ASAP7_75t_SL g3425 ( 
.A(n_3299),
.B(n_3408),
.Y(n_3425)
);

INVx3_ASAP7_75t_L g3426 ( 
.A(n_3355),
.Y(n_3426)
);

BUFx4f_ASAP7_75t_L g3427 ( 
.A(n_3355),
.Y(n_3427)
);

AOI22xp33_ASAP7_75t_L g3428 ( 
.A1(n_3397),
.A2(n_3261),
.B1(n_3188),
.B2(n_3228),
.Y(n_3428)
);

BUFx2_ASAP7_75t_L g3429 ( 
.A(n_3314),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3290),
.Y(n_3430)
);

AOI21xp5_ASAP7_75t_L g3431 ( 
.A1(n_3341),
.A2(n_3195),
.B(n_3263),
.Y(n_3431)
);

AOI21xp5_ASAP7_75t_L g3432 ( 
.A1(n_3364),
.A2(n_3249),
.B(n_3247),
.Y(n_3432)
);

AOI21xp5_ASAP7_75t_L g3433 ( 
.A1(n_3378),
.A2(n_3272),
.B(n_3271),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3319),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3328),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3293),
.Y(n_3436)
);

AO22x1_ASAP7_75t_L g3437 ( 
.A1(n_3405),
.A2(n_3228),
.B1(n_3303),
.B2(n_3296),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_3383),
.A2(n_3414),
.B(n_3332),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_3393),
.B(n_3239),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3406),
.B(n_3273),
.Y(n_3440)
);

O2A1O1Ixp33_ASAP7_75t_L g3441 ( 
.A1(n_3311),
.A2(n_3255),
.B(n_3282),
.C(n_3131),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_SL g3442 ( 
.A(n_3423),
.B(n_3197),
.Y(n_3442)
);

AOI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_3308),
.A2(n_3289),
.B(n_3146),
.Y(n_3443)
);

OR2x2_ASAP7_75t_L g3444 ( 
.A(n_3310),
.B(n_3171),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3415),
.B(n_3163),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3295),
.Y(n_3446)
);

INVxp67_ASAP7_75t_L g3447 ( 
.A(n_3385),
.Y(n_3447)
);

AOI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_3336),
.A2(n_3194),
.B(n_3180),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3417),
.B(n_3166),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3377),
.B(n_3181),
.Y(n_3450)
);

OAI21xp5_ASAP7_75t_L g3451 ( 
.A1(n_3419),
.A2(n_1837),
.B(n_1812),
.Y(n_3451)
);

BUFx6f_ASAP7_75t_L g3452 ( 
.A(n_3325),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3302),
.Y(n_3453)
);

OAI21xp33_ASAP7_75t_L g3454 ( 
.A1(n_3294),
.A2(n_1497),
.B(n_1490),
.Y(n_3454)
);

AOI21xp5_ASAP7_75t_L g3455 ( 
.A1(n_3337),
.A2(n_1607),
.B(n_1365),
.Y(n_3455)
);

INVx2_ASAP7_75t_SL g3456 ( 
.A(n_3366),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3381),
.B(n_1498),
.Y(n_3457)
);

AOI21x1_ASAP7_75t_L g3458 ( 
.A1(n_3409),
.A2(n_2046),
.B(n_1784),
.Y(n_3458)
);

O2A1O1Ixp5_ASAP7_75t_L g3459 ( 
.A1(n_3399),
.A2(n_1851),
.B(n_1853),
.C(n_1838),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_3339),
.A2(n_1471),
.B(n_1338),
.Y(n_3460)
);

AOI21xp5_ASAP7_75t_L g3461 ( 
.A1(n_3342),
.A2(n_1471),
.B(n_1338),
.Y(n_3461)
);

AO21x1_ASAP7_75t_L g3462 ( 
.A1(n_3402),
.A2(n_1869),
.B(n_1857),
.Y(n_3462)
);

NAND2x1p5_ASAP7_75t_L g3463 ( 
.A(n_3297),
.B(n_1934),
.Y(n_3463)
);

AOI21xp5_ASAP7_75t_L g3464 ( 
.A1(n_3348),
.A2(n_3389),
.B(n_3388),
.Y(n_3464)
);

AOI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_3369),
.A2(n_1504),
.B(n_1471),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3373),
.B(n_1500),
.Y(n_3466)
);

AOI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_3324),
.A2(n_3376),
.B(n_3306),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_3333),
.Y(n_3468)
);

NOR2xp33_ASAP7_75t_L g3469 ( 
.A(n_3316),
.B(n_2821),
.Y(n_3469)
);

HB1xp67_ASAP7_75t_L g3470 ( 
.A(n_3361),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_SL g3471 ( 
.A(n_3374),
.B(n_2825),
.Y(n_3471)
);

AOI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_3304),
.A2(n_1598),
.B(n_1504),
.Y(n_3472)
);

CKINVDCx10_ASAP7_75t_R g3473 ( 
.A(n_3372),
.Y(n_3473)
);

BUFx12f_ASAP7_75t_L g3474 ( 
.A(n_3404),
.Y(n_3474)
);

BUFx6f_ASAP7_75t_L g3475 ( 
.A(n_3300),
.Y(n_3475)
);

OAI22xp5_ASAP7_75t_L g3476 ( 
.A1(n_3307),
.A2(n_1507),
.B1(n_1508),
.B2(n_1501),
.Y(n_3476)
);

A2O1A1Ixp33_ASAP7_75t_L g3477 ( 
.A1(n_3400),
.A2(n_3309),
.B(n_3315),
.C(n_3313),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3413),
.B(n_3301),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3317),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3320),
.B(n_1511),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3322),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3326),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3330),
.B(n_3331),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_SL g3484 ( 
.A(n_3394),
.B(n_2826),
.Y(n_3484)
);

BUFx6f_ASAP7_75t_L g3485 ( 
.A(n_3321),
.Y(n_3485)
);

BUFx2_ASAP7_75t_L g3486 ( 
.A(n_3343),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3335),
.Y(n_3487)
);

AOI21xp5_ASAP7_75t_L g3488 ( 
.A1(n_3403),
.A2(n_1598),
.B(n_1504),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3344),
.Y(n_3489)
);

AND2x2_ASAP7_75t_L g3490 ( 
.A(n_3392),
.B(n_2056),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3345),
.Y(n_3491)
);

NOR2xp33_ASAP7_75t_L g3492 ( 
.A(n_3340),
.B(n_2840),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_3412),
.A2(n_1712),
.B(n_1598),
.Y(n_3493)
);

AOI21xp5_ASAP7_75t_L g3494 ( 
.A1(n_3422),
.A2(n_1964),
.B(n_1712),
.Y(n_3494)
);

BUFx4f_ASAP7_75t_L g3495 ( 
.A(n_3404),
.Y(n_3495)
);

AOI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_3298),
.A2(n_1964),
.B(n_1712),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3347),
.Y(n_3497)
);

NOR2xp33_ASAP7_75t_L g3498 ( 
.A(n_3418),
.B(n_1512),
.Y(n_3498)
);

AOI21x1_ASAP7_75t_L g3499 ( 
.A1(n_3391),
.A2(n_1877),
.B(n_1871),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_SL g3500 ( 
.A(n_3292),
.B(n_1281),
.Y(n_3500)
);

AOI21xp5_ASAP7_75t_L g3501 ( 
.A1(n_3380),
.A2(n_2008),
.B(n_1964),
.Y(n_3501)
);

AOI21x1_ASAP7_75t_L g3502 ( 
.A1(n_3382),
.A2(n_1896),
.B(n_1879),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3367),
.B(n_1516),
.Y(n_3503)
);

AOI21xp5_ASAP7_75t_L g3504 ( 
.A1(n_3357),
.A2(n_2008),
.B(n_1905),
.Y(n_3504)
);

HB1xp67_ASAP7_75t_L g3505 ( 
.A(n_3318),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3386),
.B(n_1517),
.Y(n_3506)
);

NOR2x1p5_ASAP7_75t_L g3507 ( 
.A(n_3387),
.B(n_1520),
.Y(n_3507)
);

OAI21xp5_ASAP7_75t_L g3508 ( 
.A1(n_3375),
.A2(n_1907),
.B(n_1902),
.Y(n_3508)
);

AND2x2_ASAP7_75t_L g3509 ( 
.A(n_3379),
.B(n_3323),
.Y(n_3509)
);

INVx2_ASAP7_75t_L g3510 ( 
.A(n_3338),
.Y(n_3510)
);

CKINVDCx10_ASAP7_75t_R g3511 ( 
.A(n_3411),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_3363),
.A2(n_2008),
.B(n_1916),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3386),
.B(n_1521),
.Y(n_3513)
);

AOI21x1_ASAP7_75t_L g3514 ( 
.A1(n_3384),
.A2(n_1918),
.B(n_1914),
.Y(n_3514)
);

O2A1O1Ixp33_ASAP7_75t_L g3515 ( 
.A1(n_3291),
.A2(n_1941),
.B(n_1943),
.C(n_1928),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3350),
.Y(n_3516)
);

AOI21xp5_ASAP7_75t_L g3517 ( 
.A1(n_3305),
.A2(n_1954),
.B(n_1950),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_3352),
.B(n_1525),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3353),
.B(n_1526),
.Y(n_3519)
);

OAI321xp33_ASAP7_75t_L g3520 ( 
.A1(n_3407),
.A2(n_1993),
.A3(n_1978),
.B1(n_2010),
.B2(n_1989),
.C(n_1961),
.Y(n_3520)
);

INVx1_ASAP7_75t_SL g3521 ( 
.A(n_3329),
.Y(n_3521)
);

NAND2x1_ASAP7_75t_L g3522 ( 
.A(n_3356),
.B(n_2012),
.Y(n_3522)
);

CKINVDCx5p33_ASAP7_75t_R g3523 ( 
.A(n_3396),
.Y(n_3523)
);

O2A1O1Ixp33_ASAP7_75t_L g3524 ( 
.A1(n_3354),
.A2(n_2014),
.B(n_2021),
.C(n_2013),
.Y(n_3524)
);

AOI21xp5_ASAP7_75t_L g3525 ( 
.A1(n_3351),
.A2(n_2027),
.B(n_2025),
.Y(n_3525)
);

AOI21xp5_ASAP7_75t_L g3526 ( 
.A1(n_3312),
.A2(n_3334),
.B(n_3359),
.Y(n_3526)
);

BUFx2_ASAP7_75t_SL g3527 ( 
.A(n_3395),
.Y(n_3527)
);

CKINVDCx8_ASAP7_75t_R g3528 ( 
.A(n_3401),
.Y(n_3528)
);

AOI21xp5_ASAP7_75t_L g3529 ( 
.A1(n_3360),
.A2(n_2036),
.B(n_2031),
.Y(n_3529)
);

AOI21xp5_ASAP7_75t_L g3530 ( 
.A1(n_3362),
.A2(n_2041),
.B(n_2040),
.Y(n_3530)
);

BUFx6f_ASAP7_75t_L g3531 ( 
.A(n_3327),
.Y(n_3531)
);

BUFx3_ASAP7_75t_L g3532 ( 
.A(n_3427),
.Y(n_3532)
);

INVx5_ASAP7_75t_L g3533 ( 
.A(n_3475),
.Y(n_3533)
);

BUFx2_ASAP7_75t_L g3534 ( 
.A(n_3452),
.Y(n_3534)
);

INVx2_ASAP7_75t_SL g3535 ( 
.A(n_3495),
.Y(n_3535)
);

INVx1_ASAP7_75t_SL g3536 ( 
.A(n_3486),
.Y(n_3536)
);

AOI22xp33_ASAP7_75t_L g3537 ( 
.A1(n_3425),
.A2(n_3421),
.B1(n_3346),
.B2(n_3358),
.Y(n_3537)
);

NOR2xp33_ASAP7_75t_R g3538 ( 
.A(n_3528),
.B(n_3365),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3483),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3434),
.Y(n_3540)
);

O2A1O1Ixp33_ASAP7_75t_L g3541 ( 
.A1(n_3441),
.A2(n_2054),
.B(n_2073),
.C(n_2043),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_SL g3542 ( 
.A(n_3464),
.B(n_3420),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_L g3543 ( 
.A(n_3498),
.B(n_3368),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_SL g3544 ( 
.A(n_3448),
.B(n_3416),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3430),
.Y(n_3545)
);

AOI22xp5_ASAP7_75t_L g3546 ( 
.A1(n_3469),
.A2(n_3390),
.B1(n_1529),
.B2(n_1534),
.Y(n_3546)
);

BUFx12f_ASAP7_75t_L g3547 ( 
.A(n_3429),
.Y(n_3547)
);

A2O1A1Ixp33_ASAP7_75t_L g3548 ( 
.A1(n_3454),
.A2(n_3370),
.B(n_3371),
.C(n_2074),
.Y(n_3548)
);

BUFx12f_ASAP7_75t_L g3549 ( 
.A(n_3474),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_SL g3550 ( 
.A(n_3428),
.B(n_3398),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3436),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3446),
.Y(n_3552)
);

NOR2xp33_ASAP7_75t_L g3553 ( 
.A(n_3447),
.B(n_1528),
.Y(n_3553)
);

AOI21xp5_ASAP7_75t_L g3554 ( 
.A1(n_3431),
.A2(n_3424),
.B(n_3443),
.Y(n_3554)
);

BUFx8_ASAP7_75t_L g3555 ( 
.A(n_3456),
.Y(n_3555)
);

NOR2xp33_ASAP7_75t_R g3556 ( 
.A(n_3523),
.B(n_3349),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3453),
.Y(n_3557)
);

BUFx6f_ASAP7_75t_L g3558 ( 
.A(n_3452),
.Y(n_3558)
);

NOR2xp33_ASAP7_75t_L g3559 ( 
.A(n_3439),
.B(n_1537),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3479),
.Y(n_3560)
);

INVx3_ASAP7_75t_L g3561 ( 
.A(n_3475),
.Y(n_3561)
);

AND2x2_ASAP7_75t_SL g3562 ( 
.A(n_3509),
.B(n_1710),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3440),
.B(n_1539),
.Y(n_3563)
);

AOI21xp5_ASAP7_75t_L g3564 ( 
.A1(n_3494),
.A2(n_1886),
.B(n_1836),
.Y(n_3564)
);

O2A1O1Ixp33_ASAP7_75t_L g3565 ( 
.A1(n_3451),
.A2(n_1936),
.B(n_1938),
.C(n_1889),
.Y(n_3565)
);

INVxp67_ASAP7_75t_SL g3566 ( 
.A(n_3467),
.Y(n_3566)
);

AOI22xp5_ASAP7_75t_L g3567 ( 
.A1(n_3478),
.A2(n_1541),
.B1(n_1544),
.B2(n_1540),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3477),
.B(n_1545),
.Y(n_3568)
);

INVx6_ASAP7_75t_L g3569 ( 
.A(n_3531),
.Y(n_3569)
);

O2A1O1Ixp33_ASAP7_75t_L g3570 ( 
.A1(n_3476),
.A2(n_1966),
.B(n_1988),
.C(n_1979),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_3432),
.A2(n_2005),
.B(n_1294),
.Y(n_3571)
);

BUFx2_ASAP7_75t_L g3572 ( 
.A(n_3505),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3481),
.B(n_1548),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3470),
.B(n_1557),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3435),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3482),
.B(n_1558),
.Y(n_3576)
);

O2A1O1Ixp5_ASAP7_75t_L g3577 ( 
.A1(n_3462),
.A2(n_2068),
.B(n_1463),
.C(n_3),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3487),
.B(n_1561),
.Y(n_3578)
);

BUFx4f_ASAP7_75t_L g3579 ( 
.A(n_3531),
.Y(n_3579)
);

BUFx6f_ASAP7_75t_L g3580 ( 
.A(n_3531),
.Y(n_3580)
);

AND2x2_ASAP7_75t_L g3581 ( 
.A(n_3503),
.B(n_1562),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_SL g3582 ( 
.A(n_3445),
.B(n_1293),
.Y(n_3582)
);

O2A1O1Ixp33_ASAP7_75t_L g3583 ( 
.A1(n_3520),
.A2(n_1957),
.B(n_1564),
.C(n_1565),
.Y(n_3583)
);

INVx1_ASAP7_75t_SL g3584 ( 
.A(n_3521),
.Y(n_3584)
);

NOR2xp33_ASAP7_75t_L g3585 ( 
.A(n_3444),
.B(n_1563),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3489),
.Y(n_3586)
);

INVx4_ASAP7_75t_L g3587 ( 
.A(n_3426),
.Y(n_3587)
);

OA21x2_ASAP7_75t_L g3588 ( 
.A1(n_3496),
.A2(n_1301),
.B(n_1297),
.Y(n_3588)
);

OAI22x1_ASAP7_75t_L g3589 ( 
.A1(n_3507),
.A2(n_1570),
.B1(n_1572),
.B2(n_1568),
.Y(n_3589)
);

AOI21xp5_ASAP7_75t_L g3590 ( 
.A1(n_3438),
.A2(n_1307),
.B(n_1306),
.Y(n_3590)
);

NOR3xp33_ASAP7_75t_L g3591 ( 
.A(n_3524),
.B(n_1574),
.C(n_1573),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_3465),
.A2(n_1318),
.B(n_1310),
.Y(n_3592)
);

INVx2_ASAP7_75t_L g3593 ( 
.A(n_3468),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3491),
.Y(n_3594)
);

INVx2_ASAP7_75t_L g3595 ( 
.A(n_3510),
.Y(n_3595)
);

BUFx2_ASAP7_75t_L g3596 ( 
.A(n_3475),
.Y(n_3596)
);

OAI22xp5_ASAP7_75t_SL g3597 ( 
.A1(n_3492),
.A2(n_1581),
.B1(n_1584),
.B2(n_1575),
.Y(n_3597)
);

BUFx8_ASAP7_75t_L g3598 ( 
.A(n_3490),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3488),
.A2(n_1333),
.B(n_1322),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3508),
.B(n_1585),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3449),
.B(n_1586),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3497),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_SL g3603 ( 
.A(n_3493),
.B(n_1334),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_3460),
.A2(n_1341),
.B(n_1339),
.Y(n_3604)
);

O2A1O1Ixp33_ASAP7_75t_L g3605 ( 
.A1(n_3515),
.A2(n_1590),
.B(n_1592),
.C(n_1587),
.Y(n_3605)
);

NOR2xp33_ASAP7_75t_L g3606 ( 
.A(n_3506),
.B(n_1593),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3450),
.B(n_1594),
.Y(n_3607)
);

AOI22xp33_ASAP7_75t_L g3608 ( 
.A1(n_3442),
.A2(n_1595),
.B1(n_1599),
.B2(n_1597),
.Y(n_3608)
);

AOI21x1_ASAP7_75t_L g3609 ( 
.A1(n_3501),
.A2(n_2068),
.B(n_1463),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_SL g3610 ( 
.A(n_3485),
.B(n_3512),
.Y(n_3610)
);

BUFx3_ASAP7_75t_L g3611 ( 
.A(n_3485),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_SL g3612 ( 
.A(n_3485),
.B(n_1345),
.Y(n_3612)
);

OAI22xp5_ASAP7_75t_L g3613 ( 
.A1(n_3500),
.A2(n_3457),
.B1(n_3466),
.B2(n_3480),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_3516),
.Y(n_3614)
);

OAI22xp5_ASAP7_75t_L g3615 ( 
.A1(n_3513),
.A2(n_1604),
.B1(n_1606),
.B2(n_1600),
.Y(n_3615)
);

OAI22xp5_ASAP7_75t_L g3616 ( 
.A1(n_3433),
.A2(n_1616),
.B1(n_1620),
.B2(n_1615),
.Y(n_3616)
);

AOI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_3461),
.A2(n_1358),
.B(n_1347),
.Y(n_3617)
);

O2A1O1Ixp33_ASAP7_75t_L g3618 ( 
.A1(n_3459),
.A2(n_1634),
.B(n_1639),
.C(n_1633),
.Y(n_3618)
);

NOR3xp33_ASAP7_75t_L g3619 ( 
.A(n_3522),
.B(n_3517),
.C(n_3437),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3527),
.B(n_1644),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3514),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_3499),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3529),
.B(n_1650),
.Y(n_3623)
);

NOR2xp33_ASAP7_75t_L g3624 ( 
.A(n_3511),
.B(n_1652),
.Y(n_3624)
);

INVx4_ASAP7_75t_L g3625 ( 
.A(n_3463),
.Y(n_3625)
);

NOR2xp33_ASAP7_75t_L g3626 ( 
.A(n_3471),
.B(n_1653),
.Y(n_3626)
);

BUFx2_ASAP7_75t_L g3627 ( 
.A(n_3518),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3530),
.B(n_3455),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_SL g3629 ( 
.A(n_3504),
.B(n_3525),
.Y(n_3629)
);

OAI22xp5_ASAP7_75t_L g3630 ( 
.A1(n_3519),
.A2(n_1663),
.B1(n_1667),
.B2(n_1660),
.Y(n_3630)
);

O2A1O1Ixp33_ASAP7_75t_L g3631 ( 
.A1(n_3472),
.A2(n_1670),
.B(n_1674),
.C(n_1669),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3484),
.B(n_1677),
.Y(n_3632)
);

OAI21x1_ASAP7_75t_L g3633 ( 
.A1(n_3458),
.A2(n_2068),
.B(n_1463),
.Y(n_3633)
);

INVx2_ASAP7_75t_L g3634 ( 
.A(n_3502),
.Y(n_3634)
);

NAND2x1p5_ASAP7_75t_L g3635 ( 
.A(n_3526),
.B(n_958),
.Y(n_3635)
);

OAI22xp5_ASAP7_75t_L g3636 ( 
.A1(n_3473),
.A2(n_1684),
.B1(n_1689),
.B2(n_1681),
.Y(n_3636)
);

AOI21xp5_ASAP7_75t_L g3637 ( 
.A1(n_3431),
.A2(n_1362),
.B(n_1361),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3439),
.B(n_1697),
.Y(n_3638)
);

AOI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3431),
.A2(n_1388),
.B(n_1368),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3439),
.B(n_1700),
.Y(n_3640)
);

NOR2xp33_ASAP7_75t_L g3641 ( 
.A(n_3498),
.B(n_1709),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3439),
.B(n_1711),
.Y(n_3642)
);

NAND2x1p5_ASAP7_75t_L g3643 ( 
.A(n_3427),
.B(n_960),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3439),
.B(n_1713),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3439),
.B(n_1718),
.Y(n_3645)
);

AOI21xp5_ASAP7_75t_L g3646 ( 
.A1(n_3431),
.A2(n_1402),
.B(n_1389),
.Y(n_3646)
);

A2O1A1Ixp33_ASAP7_75t_L g3647 ( 
.A1(n_3541),
.A2(n_1724),
.B(n_1725),
.C(n_1723),
.Y(n_3647)
);

OAI22xp5_ASAP7_75t_L g3648 ( 
.A1(n_3608),
.A2(n_1729),
.B1(n_1730),
.B2(n_1727),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_3539),
.B(n_1731),
.Y(n_3649)
);

OAI21x1_ASAP7_75t_L g3650 ( 
.A1(n_3609),
.A2(n_2068),
.B(n_1463),
.Y(n_3650)
);

BUFx3_ASAP7_75t_L g3651 ( 
.A(n_3532),
.Y(n_3651)
);

OR2x2_ASAP7_75t_L g3652 ( 
.A(n_3545),
.B(n_3551),
.Y(n_3652)
);

HB1xp67_ASAP7_75t_L g3653 ( 
.A(n_3572),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3552),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_SL g3655 ( 
.A(n_3549),
.B(n_1734),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3557),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3560),
.B(n_1739),
.Y(n_3657)
);

AOI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_3554),
.A2(n_1744),
.B(n_1741),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3586),
.Y(n_3659)
);

AOI21xp5_ASAP7_75t_L g3660 ( 
.A1(n_3566),
.A2(n_1756),
.B(n_1745),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3594),
.Y(n_3661)
);

INVx2_ASAP7_75t_SL g3662 ( 
.A(n_3558),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_3614),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3627),
.B(n_1757),
.Y(n_3664)
);

OAI21x1_ASAP7_75t_L g3665 ( 
.A1(n_3633),
.A2(n_2068),
.B(n_1463),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3602),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3540),
.Y(n_3667)
);

BUFx2_ASAP7_75t_L g3668 ( 
.A(n_3556),
.Y(n_3668)
);

AOI21xp5_ASAP7_75t_L g3669 ( 
.A1(n_3544),
.A2(n_1763),
.B(n_1759),
.Y(n_3669)
);

OAI22xp5_ASAP7_75t_L g3670 ( 
.A1(n_3641),
.A2(n_1774),
.B1(n_1777),
.B2(n_1772),
.Y(n_3670)
);

AO31x2_ASAP7_75t_L g3671 ( 
.A1(n_3634),
.A2(n_1412),
.A3(n_1416),
.B(n_1407),
.Y(n_3671)
);

AOI21x1_ASAP7_75t_L g3672 ( 
.A1(n_3542),
.A2(n_1780),
.B(n_1778),
.Y(n_3672)
);

OAI21x1_ASAP7_75t_L g3673 ( 
.A1(n_3629),
.A2(n_964),
.B(n_962),
.Y(n_3673)
);

INVx2_ASAP7_75t_SL g3674 ( 
.A(n_3558),
.Y(n_3674)
);

OAI21x1_ASAP7_75t_L g3675 ( 
.A1(n_3635),
.A2(n_972),
.B(n_970),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_L g3676 ( 
.A(n_3624),
.B(n_1781),
.Y(n_3676)
);

AOI21xp5_ASAP7_75t_L g3677 ( 
.A1(n_3603),
.A2(n_1786),
.B(n_1783),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3575),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3536),
.B(n_1792),
.Y(n_3679)
);

A2O1A1Ixp33_ASAP7_75t_L g3680 ( 
.A1(n_3600),
.A2(n_3605),
.B(n_3591),
.C(n_3559),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3584),
.B(n_1794),
.Y(n_3681)
);

AO21x1_ASAP7_75t_L g3682 ( 
.A1(n_3568),
.A2(n_1),
.B(n_2),
.Y(n_3682)
);

AOI21xp5_ASAP7_75t_L g3683 ( 
.A1(n_3628),
.A2(n_1807),
.B(n_1795),
.Y(n_3683)
);

O2A1O1Ixp5_ASAP7_75t_L g3684 ( 
.A1(n_3550),
.A2(n_5),
.B(n_3),
.C(n_4),
.Y(n_3684)
);

INVx1_ASAP7_75t_SL g3685 ( 
.A(n_3538),
.Y(n_3685)
);

NAND3xp33_ASAP7_75t_SL g3686 ( 
.A(n_3570),
.B(n_1809),
.C(n_1808),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3596),
.B(n_1810),
.Y(n_3687)
);

OAI21x1_ASAP7_75t_L g3688 ( 
.A1(n_3622),
.A2(n_976),
.B(n_975),
.Y(n_3688)
);

O2A1O1Ixp5_ASAP7_75t_L g3689 ( 
.A1(n_3577),
.A2(n_6),
.B(n_4),
.C(n_5),
.Y(n_3689)
);

OAI22xp5_ASAP7_75t_L g3690 ( 
.A1(n_3613),
.A2(n_1815),
.B1(n_1816),
.B2(n_1811),
.Y(n_3690)
);

OAI21x1_ASAP7_75t_L g3691 ( 
.A1(n_3599),
.A2(n_978),
.B(n_977),
.Y(n_3691)
);

A2O1A1Ixp33_ASAP7_75t_L g3692 ( 
.A1(n_3583),
.A2(n_1819),
.B(n_1822),
.C(n_1817),
.Y(n_3692)
);

OAI21x1_ASAP7_75t_L g3693 ( 
.A1(n_3621),
.A2(n_3610),
.B(n_3588),
.Y(n_3693)
);

HB1xp67_ASAP7_75t_L g3694 ( 
.A(n_3593),
.Y(n_3694)
);

AND2x2_ASAP7_75t_L g3695 ( 
.A(n_3534),
.B(n_7),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3595),
.Y(n_3696)
);

INVx3_ASAP7_75t_L g3697 ( 
.A(n_3579),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3573),
.Y(n_3698)
);

AO31x2_ASAP7_75t_L g3699 ( 
.A1(n_3564),
.A2(n_1426),
.A3(n_1427),
.B(n_1425),
.Y(n_3699)
);

NOR2xp67_ASAP7_75t_L g3700 ( 
.A(n_3533),
.B(n_7),
.Y(n_3700)
);

AO31x2_ASAP7_75t_L g3701 ( 
.A1(n_3548),
.A2(n_1441),
.A3(n_1447),
.B(n_1439),
.Y(n_3701)
);

OAI22x1_ASAP7_75t_L g3702 ( 
.A1(n_3546),
.A2(n_1826),
.B1(n_1828),
.B2(n_1824),
.Y(n_3702)
);

INVx1_ASAP7_75t_SL g3703 ( 
.A(n_3569),
.Y(n_3703)
);

OR2x2_ASAP7_75t_L g3704 ( 
.A(n_3576),
.B(n_8),
.Y(n_3704)
);

OA21x2_ASAP7_75t_L g3705 ( 
.A1(n_3571),
.A2(n_1839),
.B(n_1835),
.Y(n_3705)
);

BUFx2_ASAP7_75t_R g3706 ( 
.A(n_3611),
.Y(n_3706)
);

AOI21xp5_ASAP7_75t_L g3707 ( 
.A1(n_3582),
.A2(n_1842),
.B(n_1840),
.Y(n_3707)
);

AO31x2_ASAP7_75t_L g3708 ( 
.A1(n_3637),
.A2(n_1452),
.A3(n_1453),
.B(n_1451),
.Y(n_3708)
);

OAI21x1_ASAP7_75t_SL g3709 ( 
.A1(n_3618),
.A2(n_9),
.B(n_10),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3578),
.Y(n_3710)
);

OAI21xp5_ASAP7_75t_L g3711 ( 
.A1(n_3639),
.A2(n_1848),
.B(n_1843),
.Y(n_3711)
);

BUFx12f_ASAP7_75t_L g3712 ( 
.A(n_3555),
.Y(n_3712)
);

AO31x2_ASAP7_75t_L g3713 ( 
.A1(n_3646),
.A2(n_1472),
.A3(n_1480),
.B(n_1465),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_3574),
.B(n_1849),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3561),
.Y(n_3715)
);

BUFx6f_ASAP7_75t_L g3716 ( 
.A(n_3580),
.Y(n_3716)
);

AOI21xp5_ASAP7_75t_L g3717 ( 
.A1(n_3631),
.A2(n_1854),
.B(n_1850),
.Y(n_3717)
);

A2O1A1Ixp33_ASAP7_75t_L g3718 ( 
.A1(n_3606),
.A2(n_3565),
.B(n_3626),
.C(n_3585),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3569),
.Y(n_3719)
);

NOR2xp33_ASAP7_75t_L g3720 ( 
.A(n_3535),
.B(n_1858),
.Y(n_3720)
);

AND2x4_ASAP7_75t_L g3721 ( 
.A(n_3533),
.B(n_980),
.Y(n_3721)
);

NOR2xp33_ASAP7_75t_SL g3722 ( 
.A(n_3547),
.B(n_1861),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3563),
.B(n_1863),
.Y(n_3723)
);

AO31x2_ASAP7_75t_L g3724 ( 
.A1(n_3592),
.A2(n_1491),
.A3(n_1492),
.B(n_1488),
.Y(n_3724)
);

AO31x2_ASAP7_75t_L g3725 ( 
.A1(n_3604),
.A2(n_1502),
.A3(n_1522),
.B(n_1496),
.Y(n_3725)
);

NOR2xp33_ASAP7_75t_L g3726 ( 
.A(n_3587),
.B(n_1866),
.Y(n_3726)
);

AO31x2_ASAP7_75t_L g3727 ( 
.A1(n_3617),
.A2(n_1527),
.A3(n_1531),
.B(n_1524),
.Y(n_3727)
);

AOI21xp5_ASAP7_75t_L g3728 ( 
.A1(n_3616),
.A2(n_2058),
.B(n_2055),
.Y(n_3728)
);

OAI21x1_ASAP7_75t_L g3729 ( 
.A1(n_3590),
.A2(n_985),
.B(n_983),
.Y(n_3729)
);

NOR2x1_ASAP7_75t_SL g3730 ( 
.A(n_3533),
.B(n_9),
.Y(n_3730)
);

BUFx2_ASAP7_75t_L g3731 ( 
.A(n_3580),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3562),
.Y(n_3732)
);

BUFx6f_ASAP7_75t_L g3733 ( 
.A(n_3625),
.Y(n_3733)
);

OAI21x1_ASAP7_75t_L g3734 ( 
.A1(n_3643),
.A2(n_990),
.B(n_987),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3581),
.B(n_1870),
.Y(n_3735)
);

OAI21xp5_ASAP7_75t_SL g3736 ( 
.A1(n_3619),
.A2(n_11),
.B(n_12),
.Y(n_3736)
);

OAI21xp5_ASAP7_75t_SL g3737 ( 
.A1(n_3567),
.A2(n_14),
.B(n_15),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_L g3738 ( 
.A(n_3543),
.B(n_1872),
.Y(n_3738)
);

OAI21x1_ASAP7_75t_L g3739 ( 
.A1(n_3612),
.A2(n_993),
.B(n_992),
.Y(n_3739)
);

A2O1A1Ixp33_ASAP7_75t_L g3740 ( 
.A1(n_3623),
.A2(n_1874),
.B(n_1875),
.C(n_1873),
.Y(n_3740)
);

OAI21x1_ASAP7_75t_L g3741 ( 
.A1(n_3537),
.A2(n_997),
.B(n_994),
.Y(n_3741)
);

OAI21x1_ASAP7_75t_L g3742 ( 
.A1(n_3601),
.A2(n_1002),
.B(n_1001),
.Y(n_3742)
);

NAND3xp33_ASAP7_75t_L g3743 ( 
.A(n_3553),
.B(n_1893),
.C(n_1888),
.Y(n_3743)
);

OAI22xp5_ASAP7_75t_L g3744 ( 
.A1(n_3597),
.A2(n_1922),
.B1(n_1968),
.B2(n_1906),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3607),
.Y(n_3745)
);

NOR2x1_ASAP7_75t_SL g3746 ( 
.A(n_3652),
.B(n_3620),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3654),
.Y(n_3747)
);

O2A1O1Ixp33_ASAP7_75t_SL g3748 ( 
.A1(n_3718),
.A2(n_3638),
.B(n_3642),
.C(n_3640),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3656),
.Y(n_3749)
);

OAI22xp5_ASAP7_75t_L g3750 ( 
.A1(n_3736),
.A2(n_3644),
.B1(n_3645),
.B2(n_3636),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3663),
.Y(n_3751)
);

BUFx2_ASAP7_75t_L g3752 ( 
.A(n_3653),
.Y(n_3752)
);

OR2x2_ASAP7_75t_L g3753 ( 
.A(n_3659),
.B(n_3632),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3661),
.Y(n_3754)
);

BUFx6f_ASAP7_75t_L g3755 ( 
.A(n_3651),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3666),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3694),
.Y(n_3757)
);

OAI22xp5_ASAP7_75t_L g3758 ( 
.A1(n_3737),
.A2(n_3630),
.B1(n_3615),
.B2(n_1900),
.Y(n_3758)
);

AOI21xp5_ASAP7_75t_L g3759 ( 
.A1(n_3680),
.A2(n_3589),
.B(n_1901),
.Y(n_3759)
);

NAND3xp33_ASAP7_75t_L g3760 ( 
.A(n_3690),
.B(n_3598),
.C(n_1904),
.Y(n_3760)
);

CKINVDCx16_ASAP7_75t_R g3761 ( 
.A(n_3712),
.Y(n_3761)
);

OAI221xp5_ASAP7_75t_L g3762 ( 
.A1(n_3676),
.A2(n_1913),
.B1(n_1917),
.B2(n_1912),
.C(n_1894),
.Y(n_3762)
);

AO32x2_ASAP7_75t_L g3763 ( 
.A1(n_3662),
.A2(n_19),
.A3(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_3763)
);

OAI21x1_ASAP7_75t_L g3764 ( 
.A1(n_3650),
.A2(n_1007),
.B(n_1004),
.Y(n_3764)
);

AOI221xp5_ASAP7_75t_L g3765 ( 
.A1(n_3670),
.A2(n_3744),
.B1(n_3648),
.B2(n_3682),
.C(n_3702),
.Y(n_3765)
);

BUFx2_ASAP7_75t_L g3766 ( 
.A(n_3731),
.Y(n_3766)
);

AND2x2_ASAP7_75t_L g3767 ( 
.A(n_3695),
.B(n_18),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3667),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3678),
.Y(n_3769)
);

OAI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_3658),
.A2(n_3660),
.B(n_3683),
.Y(n_3770)
);

AOI22xp33_ASAP7_75t_SL g3771 ( 
.A1(n_3732),
.A2(n_3668),
.B1(n_3745),
.B2(n_3705),
.Y(n_3771)
);

BUFx2_ASAP7_75t_R g3772 ( 
.A(n_3738),
.Y(n_3772)
);

AND2x4_ASAP7_75t_L g3773 ( 
.A(n_3719),
.B(n_1009),
.Y(n_3773)
);

CKINVDCx11_ASAP7_75t_R g3774 ( 
.A(n_3685),
.Y(n_3774)
);

BUFx3_ASAP7_75t_L g3775 ( 
.A(n_3733),
.Y(n_3775)
);

OAI21x1_ASAP7_75t_L g3776 ( 
.A1(n_3665),
.A2(n_1014),
.B(n_1010),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3698),
.B(n_3710),
.Y(n_3777)
);

OAI21x1_ASAP7_75t_L g3778 ( 
.A1(n_3693),
.A2(n_1018),
.B(n_1016),
.Y(n_3778)
);

AOI22xp5_ASAP7_75t_L g3779 ( 
.A1(n_3686),
.A2(n_1921),
.B1(n_1924),
.B2(n_1919),
.Y(n_3779)
);

OR2x6_ASAP7_75t_L g3780 ( 
.A(n_3674),
.B(n_1020),
.Y(n_3780)
);

NOR2xp67_ASAP7_75t_L g3781 ( 
.A(n_3704),
.B(n_20),
.Y(n_3781)
);

OA21x2_ASAP7_75t_L g3782 ( 
.A1(n_3715),
.A2(n_1931),
.B(n_1927),
.Y(n_3782)
);

INVx3_ASAP7_75t_L g3783 ( 
.A(n_3716),
.Y(n_3783)
);

O2A1O1Ixp33_ASAP7_75t_L g3784 ( 
.A1(n_3647),
.A2(n_2065),
.B(n_2066),
.C(n_2062),
.Y(n_3784)
);

OAI21x1_ASAP7_75t_L g3785 ( 
.A1(n_3673),
.A2(n_1024),
.B(n_1022),
.Y(n_3785)
);

AOI21xp5_ASAP7_75t_L g3786 ( 
.A1(n_3692),
.A2(n_1937),
.B(n_1932),
.Y(n_3786)
);

AND2x4_ASAP7_75t_L g3787 ( 
.A(n_3703),
.B(n_1028),
.Y(n_3787)
);

OAI211xp5_ASAP7_75t_L g3788 ( 
.A1(n_3740),
.A2(n_1947),
.B(n_1948),
.C(n_1944),
.Y(n_3788)
);

CKINVDCx5p33_ASAP7_75t_R g3789 ( 
.A(n_3733),
.Y(n_3789)
);

OR2x6_ASAP7_75t_L g3790 ( 
.A(n_3716),
.B(n_1030),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3696),
.Y(n_3791)
);

NOR2xp33_ASAP7_75t_L g3792 ( 
.A(n_3722),
.B(n_21),
.Y(n_3792)
);

OAI21x1_ASAP7_75t_L g3793 ( 
.A1(n_3675),
.A2(n_1033),
.B(n_1031),
.Y(n_3793)
);

AO21x2_ASAP7_75t_L g3794 ( 
.A1(n_3709),
.A2(n_1554),
.B(n_1550),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3657),
.Y(n_3795)
);

NOR2x1_ASAP7_75t_SL g3796 ( 
.A(n_3672),
.B(n_21),
.Y(n_3796)
);

OAI21x1_ASAP7_75t_L g3797 ( 
.A1(n_3688),
.A2(n_1035),
.B(n_1034),
.Y(n_3797)
);

OAI21x1_ASAP7_75t_L g3798 ( 
.A1(n_3741),
.A2(n_1037),
.B(n_1036),
.Y(n_3798)
);

OR2x2_ASAP7_75t_L g3799 ( 
.A(n_3664),
.B(n_22),
.Y(n_3799)
);

INVx2_ASAP7_75t_L g3800 ( 
.A(n_3730),
.Y(n_3800)
);

INVx2_ASAP7_75t_L g3801 ( 
.A(n_3742),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3649),
.Y(n_3802)
);

OAI21x1_ASAP7_75t_L g3803 ( 
.A1(n_3729),
.A2(n_1045),
.B(n_1040),
.Y(n_3803)
);

AO21x1_ASAP7_75t_L g3804 ( 
.A1(n_3726),
.A2(n_22),
.B(n_23),
.Y(n_3804)
);

OAI21x1_ASAP7_75t_L g3805 ( 
.A1(n_3734),
.A2(n_1047),
.B(n_1046),
.Y(n_3805)
);

OAI21x1_ASAP7_75t_L g3806 ( 
.A1(n_3691),
.A2(n_3689),
.B(n_3739),
.Y(n_3806)
);

INVx2_ASAP7_75t_L g3807 ( 
.A(n_3671),
.Y(n_3807)
);

BUFx4f_ASAP7_75t_SL g3808 ( 
.A(n_3697),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3706),
.Y(n_3809)
);

AOI21xp5_ASAP7_75t_L g3810 ( 
.A1(n_3684),
.A2(n_1951),
.B(n_1949),
.Y(n_3810)
);

OAI21x1_ASAP7_75t_L g3811 ( 
.A1(n_3700),
.A2(n_1049),
.B(n_1048),
.Y(n_3811)
);

AO32x2_ASAP7_75t_L g3812 ( 
.A1(n_3671),
.A2(n_25),
.A3(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_3812)
);

INVxp67_ASAP7_75t_SL g3813 ( 
.A(n_3687),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3735),
.B(n_24),
.Y(n_3814)
);

OAI21x1_ASAP7_75t_L g3815 ( 
.A1(n_3669),
.A2(n_1051),
.B(n_1050),
.Y(n_3815)
);

AND2x4_ASAP7_75t_L g3816 ( 
.A(n_3721),
.B(n_1053),
.Y(n_3816)
);

OAI21x1_ASAP7_75t_L g3817 ( 
.A1(n_3711),
.A2(n_1056),
.B(n_1055),
.Y(n_3817)
);

OAI21x1_ASAP7_75t_L g3818 ( 
.A1(n_3677),
.A2(n_1060),
.B(n_1058),
.Y(n_3818)
);

INVx2_ASAP7_75t_L g3819 ( 
.A(n_3701),
.Y(n_3819)
);

AND2x2_ASAP7_75t_L g3820 ( 
.A(n_3720),
.B(n_27),
.Y(n_3820)
);

OR2x6_ASAP7_75t_L g3821 ( 
.A(n_3679),
.B(n_1061),
.Y(n_3821)
);

OAI21x1_ASAP7_75t_L g3822 ( 
.A1(n_3707),
.A2(n_1067),
.B(n_1065),
.Y(n_3822)
);

NOR2xp33_ASAP7_75t_SL g3823 ( 
.A(n_3655),
.B(n_1953),
.Y(n_3823)
);

NAND2x1_ASAP7_75t_L g3824 ( 
.A(n_3743),
.B(n_3681),
.Y(n_3824)
);

INVx3_ASAP7_75t_L g3825 ( 
.A(n_3755),
.Y(n_3825)
);

HB1xp67_ASAP7_75t_L g3826 ( 
.A(n_3752),
.Y(n_3826)
);

INVx3_ASAP7_75t_L g3827 ( 
.A(n_3755),
.Y(n_3827)
);

INVx2_ASAP7_75t_L g3828 ( 
.A(n_3757),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3747),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3749),
.Y(n_3830)
);

HB1xp67_ASAP7_75t_L g3831 ( 
.A(n_3766),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3754),
.Y(n_3832)
);

INVx2_ASAP7_75t_L g3833 ( 
.A(n_3751),
.Y(n_3833)
);

INVx2_ASAP7_75t_L g3834 ( 
.A(n_3769),
.Y(n_3834)
);

BUFx10_ASAP7_75t_L g3835 ( 
.A(n_3789),
.Y(n_3835)
);

OA21x2_ASAP7_75t_L g3836 ( 
.A1(n_3777),
.A2(n_3714),
.B(n_3723),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3756),
.Y(n_3837)
);

BUFx6f_ASAP7_75t_L g3838 ( 
.A(n_3775),
.Y(n_3838)
);

INVx2_ASAP7_75t_L g3839 ( 
.A(n_3768),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3791),
.Y(n_3840)
);

OAI21x1_ASAP7_75t_L g3841 ( 
.A1(n_3807),
.A2(n_3717),
.B(n_3728),
.Y(n_3841)
);

INVx4_ASAP7_75t_SL g3842 ( 
.A(n_3808),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3753),
.Y(n_3843)
);

BUFx6f_ASAP7_75t_SL g3844 ( 
.A(n_3809),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3746),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3801),
.Y(n_3846)
);

HB1xp67_ASAP7_75t_L g3847 ( 
.A(n_3813),
.Y(n_3847)
);

OR2x2_ASAP7_75t_L g3848 ( 
.A(n_3795),
.B(n_3701),
.Y(n_3848)
);

AOI22xp33_ASAP7_75t_L g3849 ( 
.A1(n_3804),
.A2(n_1959),
.B1(n_1969),
.B2(n_1956),
.Y(n_3849)
);

INVx3_ASAP7_75t_L g3850 ( 
.A(n_3783),
.Y(n_3850)
);

AOI22xp5_ASAP7_75t_L g3851 ( 
.A1(n_3750),
.A2(n_1977),
.B1(n_1980),
.B2(n_1971),
.Y(n_3851)
);

INVx4_ASAP7_75t_L g3852 ( 
.A(n_3774),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3819),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3800),
.Y(n_3854)
);

INVx6_ASAP7_75t_L g3855 ( 
.A(n_3761),
.Y(n_3855)
);

OAI22xp5_ASAP7_75t_L g3856 ( 
.A1(n_3765),
.A2(n_1982),
.B1(n_1983),
.B2(n_1981),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3802),
.Y(n_3857)
);

OAI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_3770),
.A2(n_1987),
.B1(n_1991),
.B2(n_1984),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3763),
.Y(n_3859)
);

CKINVDCx11_ASAP7_75t_R g3860 ( 
.A(n_3821),
.Y(n_3860)
);

INVx2_ASAP7_75t_L g3861 ( 
.A(n_3763),
.Y(n_3861)
);

OAI22xp33_ASAP7_75t_L g3862 ( 
.A1(n_3821),
.A2(n_2076),
.B1(n_1997),
.B2(n_2000),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3767),
.B(n_3725),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3812),
.Y(n_3864)
);

AOI22xp33_ASAP7_75t_L g3865 ( 
.A1(n_3771),
.A2(n_2001),
.B1(n_2002),
.B2(n_1996),
.Y(n_3865)
);

INVx2_ASAP7_75t_SL g3866 ( 
.A(n_3787),
.Y(n_3866)
);

AO21x1_ASAP7_75t_SL g3867 ( 
.A1(n_3814),
.A2(n_3713),
.B(n_3708),
.Y(n_3867)
);

AND2x2_ASAP7_75t_L g3868 ( 
.A(n_3820),
.B(n_3781),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3772),
.B(n_3725),
.Y(n_3869)
);

HB1xp67_ASAP7_75t_L g3870 ( 
.A(n_3799),
.Y(n_3870)
);

AND2x2_ASAP7_75t_L g3871 ( 
.A(n_3792),
.B(n_3727),
.Y(n_3871)
);

AND2x2_ASAP7_75t_L g3872 ( 
.A(n_3782),
.B(n_3727),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3812),
.Y(n_3873)
);

INVx3_ASAP7_75t_L g3874 ( 
.A(n_3773),
.Y(n_3874)
);

INVx3_ASAP7_75t_L g3875 ( 
.A(n_3780),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3778),
.Y(n_3876)
);

INVx5_ASAP7_75t_SL g3877 ( 
.A(n_3780),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3806),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3797),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3748),
.Y(n_3880)
);

INVx2_ASAP7_75t_L g3881 ( 
.A(n_3803),
.Y(n_3881)
);

INVx2_ASAP7_75t_L g3882 ( 
.A(n_3811),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3824),
.Y(n_3883)
);

INVx3_ASAP7_75t_L g3884 ( 
.A(n_3790),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3798),
.Y(n_3885)
);

HB1xp67_ASAP7_75t_L g3886 ( 
.A(n_3794),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3793),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3764),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3805),
.Y(n_3889)
);

OAI21x1_ASAP7_75t_L g3890 ( 
.A1(n_3776),
.A2(n_3817),
.B(n_3785),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3759),
.B(n_3699),
.Y(n_3891)
);

BUFx6f_ASAP7_75t_L g3892 ( 
.A(n_3816),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3790),
.Y(n_3893)
);

OAI21x1_ASAP7_75t_L g3894 ( 
.A1(n_3818),
.A2(n_3699),
.B(n_3708),
.Y(n_3894)
);

BUFx4f_ASAP7_75t_SL g3895 ( 
.A(n_3823),
.Y(n_3895)
);

HB1xp67_ASAP7_75t_L g3896 ( 
.A(n_3822),
.Y(n_3896)
);

BUFx2_ASAP7_75t_L g3897 ( 
.A(n_3815),
.Y(n_3897)
);

AOI22xp33_ASAP7_75t_L g3898 ( 
.A1(n_3758),
.A2(n_2009),
.B1(n_2011),
.B2(n_2006),
.Y(n_3898)
);

CKINVDCx20_ASAP7_75t_R g3899 ( 
.A(n_3760),
.Y(n_3899)
);

HB1xp67_ASAP7_75t_L g3900 ( 
.A(n_3796),
.Y(n_3900)
);

OAI21x1_ASAP7_75t_L g3901 ( 
.A1(n_3810),
.A2(n_3713),
.B(n_3724),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3788),
.Y(n_3902)
);

AOI22xp33_ASAP7_75t_L g3903 ( 
.A1(n_3861),
.A2(n_3786),
.B1(n_3762),
.B2(n_3779),
.Y(n_3903)
);

INVx2_ASAP7_75t_L g3904 ( 
.A(n_3846),
.Y(n_3904)
);

AOI22xp33_ASAP7_75t_L g3905 ( 
.A1(n_3859),
.A2(n_3871),
.B1(n_3873),
.B2(n_3864),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3847),
.B(n_3724),
.Y(n_3906)
);

INVx2_ASAP7_75t_L g3907 ( 
.A(n_3857),
.Y(n_3907)
);

OAI22xp5_ASAP7_75t_L g3908 ( 
.A1(n_3880),
.A2(n_3784),
.B1(n_2019),
.B2(n_2022),
.Y(n_3908)
);

AOI22xp33_ASAP7_75t_L g3909 ( 
.A1(n_3863),
.A2(n_2024),
.B1(n_2026),
.B2(n_2018),
.Y(n_3909)
);

AOI22xp33_ASAP7_75t_SL g3910 ( 
.A1(n_3869),
.A2(n_2071),
.B1(n_2044),
.B2(n_2033),
.Y(n_3910)
);

INVx3_ASAP7_75t_L g3911 ( 
.A(n_3855),
.Y(n_3911)
);

OAI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_3877),
.A2(n_2034),
.B1(n_2038),
.B2(n_2030),
.Y(n_3912)
);

BUFx4f_ASAP7_75t_SL g3913 ( 
.A(n_3852),
.Y(n_3913)
);

AOI22xp33_ASAP7_75t_L g3914 ( 
.A1(n_3872),
.A2(n_2045),
.B1(n_2050),
.B2(n_2042),
.Y(n_3914)
);

OAI22xp5_ASAP7_75t_L g3915 ( 
.A1(n_3877),
.A2(n_2070),
.B1(n_2072),
.B2(n_2069),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3854),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3829),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3830),
.Y(n_3918)
);

AOI22xp33_ASAP7_75t_SL g3919 ( 
.A1(n_3836),
.A2(n_1614),
.B1(n_1642),
.B2(n_1555),
.Y(n_3919)
);

OAI21xp33_ASAP7_75t_L g3920 ( 
.A1(n_3851),
.A2(n_28),
.B(n_29),
.Y(n_3920)
);

AOI22xp5_ASAP7_75t_L g3921 ( 
.A1(n_3883),
.A2(n_1567),
.B1(n_1576),
.B2(n_1559),
.Y(n_3921)
);

HB1xp67_ASAP7_75t_L g3922 ( 
.A(n_3826),
.Y(n_3922)
);

CKINVDCx5p33_ASAP7_75t_R g3923 ( 
.A(n_3844),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3839),
.Y(n_3924)
);

BUFx4f_ASAP7_75t_SL g3925 ( 
.A(n_3835),
.Y(n_3925)
);

AND2x2_ASAP7_75t_L g3926 ( 
.A(n_3831),
.B(n_28),
.Y(n_3926)
);

NOR2xp33_ASAP7_75t_L g3927 ( 
.A(n_3860),
.B(n_29),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3832),
.Y(n_3928)
);

AOI22xp33_ASAP7_75t_L g3929 ( 
.A1(n_3891),
.A2(n_1603),
.B1(n_1608),
.B2(n_1591),
.Y(n_3929)
);

OAI22xp5_ASAP7_75t_L g3930 ( 
.A1(n_3865),
.A2(n_1618),
.B1(n_1619),
.B2(n_1610),
.Y(n_3930)
);

CKINVDCx5p33_ASAP7_75t_R g3931 ( 
.A(n_3895),
.Y(n_3931)
);

OAI22xp33_ASAP7_75t_L g3932 ( 
.A1(n_3875),
.A2(n_1679),
.B1(n_1705),
.B2(n_1636),
.Y(n_3932)
);

AOI22xp33_ASAP7_75t_L g3933 ( 
.A1(n_3867),
.A2(n_3849),
.B1(n_3886),
.B2(n_3856),
.Y(n_3933)
);

AOI22xp33_ASAP7_75t_L g3934 ( 
.A1(n_3902),
.A2(n_1631),
.B1(n_1640),
.B2(n_1630),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3837),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3840),
.Y(n_3936)
);

INVx3_ASAP7_75t_L g3937 ( 
.A(n_3838),
.Y(n_3937)
);

AOI22xp33_ASAP7_75t_SL g3938 ( 
.A1(n_3897),
.A2(n_1695),
.B1(n_1758),
.B2(n_1651),
.Y(n_3938)
);

AOI22xp33_ASAP7_75t_L g3939 ( 
.A1(n_3848),
.A2(n_1643),
.B1(n_1664),
.B2(n_1641),
.Y(n_3939)
);

AOI22xp33_ASAP7_75t_L g3940 ( 
.A1(n_3858),
.A2(n_1678),
.B1(n_1691),
.B2(n_1673),
.Y(n_3940)
);

AOI22xp33_ASAP7_75t_L g3941 ( 
.A1(n_3900),
.A2(n_3868),
.B1(n_3901),
.B2(n_3870),
.Y(n_3941)
);

AOI22xp33_ASAP7_75t_L g3942 ( 
.A1(n_3894),
.A2(n_1693),
.B1(n_1694),
.B2(n_1692),
.Y(n_3942)
);

AOI22xp33_ASAP7_75t_L g3943 ( 
.A1(n_3862),
.A2(n_1702),
.B1(n_1707),
.B2(n_1698),
.Y(n_3943)
);

AOI22xp5_ASAP7_75t_L g3944 ( 
.A1(n_3845),
.A2(n_1737),
.B1(n_1742),
.B2(n_1708),
.Y(n_3944)
);

AOI22xp33_ASAP7_75t_L g3945 ( 
.A1(n_3882),
.A2(n_1760),
.B1(n_1761),
.B2(n_1754),
.Y(n_3945)
);

BUFx2_ASAP7_75t_L g3946 ( 
.A(n_3825),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3843),
.Y(n_3947)
);

AOI22xp33_ASAP7_75t_L g3948 ( 
.A1(n_3896),
.A2(n_1779),
.B1(n_1785),
.B2(n_1764),
.Y(n_3948)
);

INVx3_ASAP7_75t_L g3949 ( 
.A(n_3838),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3828),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3878),
.B(n_30),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3833),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3850),
.B(n_31),
.Y(n_3953)
);

AOI22xp33_ASAP7_75t_SL g3954 ( 
.A1(n_3884),
.A2(n_1860),
.B1(n_1909),
.B2(n_1801),
.Y(n_3954)
);

AOI22xp33_ASAP7_75t_L g3955 ( 
.A1(n_3876),
.A2(n_1791),
.B1(n_1793),
.B2(n_1788),
.Y(n_3955)
);

INVx3_ASAP7_75t_L g3956 ( 
.A(n_3827),
.Y(n_3956)
);

INVx2_ASAP7_75t_L g3957 ( 
.A(n_3834),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3853),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3887),
.Y(n_3959)
);

BUFx2_ASAP7_75t_L g3960 ( 
.A(n_3874),
.Y(n_3960)
);

AOI22xp33_ASAP7_75t_L g3961 ( 
.A1(n_3889),
.A2(n_1805),
.B1(n_1823),
.B2(n_1798),
.Y(n_3961)
);

AOI22xp33_ASAP7_75t_L g3962 ( 
.A1(n_3879),
.A2(n_3899),
.B1(n_3885),
.B2(n_3881),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_3866),
.B(n_33),
.Y(n_3963)
);

AOI22xp33_ASAP7_75t_L g3964 ( 
.A1(n_3893),
.A2(n_1846),
.B1(n_1852),
.B2(n_1831),
.Y(n_3964)
);

INVx8_ASAP7_75t_L g3965 ( 
.A(n_3892),
.Y(n_3965)
);

AOI22xp33_ASAP7_75t_L g3966 ( 
.A1(n_3841),
.A2(n_3888),
.B1(n_3898),
.B2(n_3890),
.Y(n_3966)
);

INVx3_ASAP7_75t_L g3967 ( 
.A(n_3892),
.Y(n_3967)
);

AOI22xp5_ASAP7_75t_L g3968 ( 
.A1(n_3842),
.A2(n_1856),
.B1(n_1867),
.B2(n_1855),
.Y(n_3968)
);

HB1xp67_ASAP7_75t_L g3969 ( 
.A(n_3842),
.Y(n_3969)
);

AOI22xp33_ASAP7_75t_L g3970 ( 
.A1(n_3861),
.A2(n_1880),
.B1(n_1881),
.B2(n_1878),
.Y(n_3970)
);

INVx4_ASAP7_75t_L g3971 ( 
.A(n_3855),
.Y(n_3971)
);

AND2x2_ASAP7_75t_L g3972 ( 
.A(n_3960),
.B(n_33),
.Y(n_3972)
);

AND2x4_ASAP7_75t_L g3973 ( 
.A(n_3946),
.B(n_34),
.Y(n_3973)
);

INVxp67_ASAP7_75t_L g3974 ( 
.A(n_3922),
.Y(n_3974)
);

NAND2x1p5_ASAP7_75t_L g3975 ( 
.A(n_3971),
.B(n_34),
.Y(n_3975)
);

XNOR2xp5_ASAP7_75t_L g3976 ( 
.A(n_3931),
.B(n_35),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3956),
.B(n_3941),
.Y(n_3977)
);

OR2x6_ASAP7_75t_L g3978 ( 
.A(n_3969),
.B(n_35),
.Y(n_3978)
);

INVxp67_ASAP7_75t_L g3979 ( 
.A(n_3906),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3917),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_3967),
.B(n_36),
.Y(n_3981)
);

NAND2xp33_ASAP7_75t_R g3982 ( 
.A(n_3923),
.B(n_38),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3959),
.B(n_37),
.Y(n_3983)
);

NAND2xp33_ASAP7_75t_R g3984 ( 
.A(n_3927),
.B(n_38),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_SL g3985 ( 
.A(n_3911),
.B(n_1885),
.Y(n_3985)
);

BUFx10_ASAP7_75t_L g3986 ( 
.A(n_3913),
.Y(n_3986)
);

INVxp67_ASAP7_75t_L g3987 ( 
.A(n_3951),
.Y(n_3987)
);

AND2x4_ASAP7_75t_L g3988 ( 
.A(n_3947),
.B(n_37),
.Y(n_3988)
);

NAND2xp33_ASAP7_75t_R g3989 ( 
.A(n_3926),
.B(n_40),
.Y(n_3989)
);

AND2x2_ASAP7_75t_L g3990 ( 
.A(n_3937),
.B(n_39),
.Y(n_3990)
);

INVx8_ASAP7_75t_L g3991 ( 
.A(n_3965),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_3904),
.Y(n_3992)
);

NAND2xp33_ASAP7_75t_R g3993 ( 
.A(n_3949),
.B(n_3953),
.Y(n_3993)
);

NOR2x1_ASAP7_75t_L g3994 ( 
.A(n_3963),
.B(n_40),
.Y(n_3994)
);

BUFx6f_ASAP7_75t_L g3995 ( 
.A(n_3965),
.Y(n_3995)
);

OR2x6_ASAP7_75t_L g3996 ( 
.A(n_3912),
.B(n_41),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_3958),
.Y(n_3997)
);

NOR2xp33_ASAP7_75t_L g3998 ( 
.A(n_3925),
.B(n_42),
.Y(n_3998)
);

NOR2xp33_ASAP7_75t_R g3999 ( 
.A(n_3903),
.B(n_42),
.Y(n_3999)
);

AND2x2_ASAP7_75t_L g4000 ( 
.A(n_3905),
.B(n_43),
.Y(n_4000)
);

NOR2xp33_ASAP7_75t_R g4001 ( 
.A(n_3933),
.B(n_43),
.Y(n_4001)
);

NOR2xp33_ASAP7_75t_R g4002 ( 
.A(n_3909),
.B(n_45),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_L g4003 ( 
.A(n_3918),
.B(n_45),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3928),
.Y(n_4004)
);

NAND2xp33_ASAP7_75t_R g4005 ( 
.A(n_3916),
.B(n_47),
.Y(n_4005)
);

AND2x4_ASAP7_75t_L g4006 ( 
.A(n_3935),
.B(n_46),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_SL g4007 ( 
.A(n_3966),
.B(n_1892),
.Y(n_4007)
);

NOR2xp33_ASAP7_75t_R g4008 ( 
.A(n_3970),
.B(n_3948),
.Y(n_4008)
);

NAND2xp33_ASAP7_75t_R g4009 ( 
.A(n_3950),
.B(n_3952),
.Y(n_4009)
);

INVxp67_ASAP7_75t_L g4010 ( 
.A(n_3924),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3907),
.Y(n_4011)
);

INVx2_ASAP7_75t_L g4012 ( 
.A(n_3936),
.Y(n_4012)
);

BUFx10_ASAP7_75t_L g4013 ( 
.A(n_3915),
.Y(n_4013)
);

AND2x2_ASAP7_75t_L g4014 ( 
.A(n_3962),
.B(n_46),
.Y(n_4014)
);

OR2x6_ASAP7_75t_L g4015 ( 
.A(n_3920),
.B(n_47),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3939),
.B(n_48),
.Y(n_4016)
);

NOR2xp33_ASAP7_75t_R g4017 ( 
.A(n_3914),
.B(n_48),
.Y(n_4017)
);

XOR2xp5_ASAP7_75t_L g4018 ( 
.A(n_3910),
.B(n_49),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3957),
.B(n_49),
.Y(n_4019)
);

AND2x4_ASAP7_75t_L g4020 ( 
.A(n_3944),
.B(n_50),
.Y(n_4020)
);

AND2x4_ASAP7_75t_L g4021 ( 
.A(n_3921),
.B(n_51),
.Y(n_4021)
);

INVxp67_ASAP7_75t_L g4022 ( 
.A(n_3919),
.Y(n_4022)
);

NOR2xp33_ASAP7_75t_R g4023 ( 
.A(n_3934),
.B(n_53),
.Y(n_4023)
);

BUFx6f_ASAP7_75t_L g4024 ( 
.A(n_3954),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_3938),
.B(n_53),
.Y(n_4025)
);

XOR2xp5_ASAP7_75t_L g4026 ( 
.A(n_3968),
.B(n_54),
.Y(n_4026)
);

NOR2xp33_ASAP7_75t_R g4027 ( 
.A(n_3942),
.B(n_54),
.Y(n_4027)
);

AND2x4_ASAP7_75t_L g4028 ( 
.A(n_3929),
.B(n_55),
.Y(n_4028)
);

NAND2xp33_ASAP7_75t_R g4029 ( 
.A(n_3932),
.B(n_56),
.Y(n_4029)
);

CKINVDCx5p33_ASAP7_75t_R g4030 ( 
.A(n_3908),
.Y(n_4030)
);

NOR2xp33_ASAP7_75t_R g4031 ( 
.A(n_3945),
.B(n_55),
.Y(n_4031)
);

BUFx3_ASAP7_75t_L g4032 ( 
.A(n_3930),
.Y(n_4032)
);

NOR2xp33_ASAP7_75t_R g4033 ( 
.A(n_3943),
.B(n_56),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3964),
.B(n_57),
.Y(n_4034)
);

NAND2xp33_ASAP7_75t_SL g4035 ( 
.A(n_3961),
.B(n_57),
.Y(n_4035)
);

BUFx6f_ASAP7_75t_L g4036 ( 
.A(n_3955),
.Y(n_4036)
);

CKINVDCx20_ASAP7_75t_R g4037 ( 
.A(n_3940),
.Y(n_4037)
);

XOR2xp5_ASAP7_75t_L g4038 ( 
.A(n_3923),
.B(n_58),
.Y(n_4038)
);

NOR2xp33_ASAP7_75t_R g4039 ( 
.A(n_3923),
.B(n_59),
.Y(n_4039)
);

NOR2xp33_ASAP7_75t_R g4040 ( 
.A(n_3923),
.B(n_60),
.Y(n_4040)
);

AND2x4_ASAP7_75t_L g4041 ( 
.A(n_3946),
.B(n_60),
.Y(n_4041)
);

NOR2xp33_ASAP7_75t_L g4042 ( 
.A(n_3913),
.B(n_61),
.Y(n_4042)
);

BUFx10_ASAP7_75t_L g4043 ( 
.A(n_3927),
.Y(n_4043)
);

BUFx10_ASAP7_75t_L g4044 ( 
.A(n_3927),
.Y(n_4044)
);

NAND2xp33_ASAP7_75t_R g4045 ( 
.A(n_3923),
.B(n_62),
.Y(n_4045)
);

AND2x4_ASAP7_75t_L g4046 ( 
.A(n_3946),
.B(n_61),
.Y(n_4046)
);

CKINVDCx5p33_ASAP7_75t_R g4047 ( 
.A(n_3931),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_3960),
.B(n_62),
.Y(n_4048)
);

NAND2xp33_ASAP7_75t_R g4049 ( 
.A(n_3923),
.B(n_64),
.Y(n_4049)
);

NAND2xp33_ASAP7_75t_R g4050 ( 
.A(n_3923),
.B(n_64),
.Y(n_4050)
);

INVxp67_ASAP7_75t_L g4051 ( 
.A(n_3922),
.Y(n_4051)
);

NOR2xp33_ASAP7_75t_R g4052 ( 
.A(n_3923),
.B(n_63),
.Y(n_4052)
);

CKINVDCx5p33_ASAP7_75t_R g4053 ( 
.A(n_3931),
.Y(n_4053)
);

CKINVDCx8_ASAP7_75t_R g4054 ( 
.A(n_3931),
.Y(n_4054)
);

INVxp67_ASAP7_75t_L g4055 ( 
.A(n_3922),
.Y(n_4055)
);

INVxp67_ASAP7_75t_L g4056 ( 
.A(n_3922),
.Y(n_4056)
);

BUFx3_ASAP7_75t_L g4057 ( 
.A(n_3931),
.Y(n_4057)
);

CKINVDCx20_ASAP7_75t_R g4058 ( 
.A(n_3913),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_3960),
.B(n_65),
.Y(n_4059)
);

BUFx4f_ASAP7_75t_L g4060 ( 
.A(n_3965),
.Y(n_4060)
);

NOR2xp33_ASAP7_75t_R g4061 ( 
.A(n_3923),
.B(n_66),
.Y(n_4061)
);

NAND2xp33_ASAP7_75t_R g4062 ( 
.A(n_3923),
.B(n_68),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3917),
.Y(n_4063)
);

BUFx3_ASAP7_75t_L g4064 ( 
.A(n_3931),
.Y(n_4064)
);

NOR2xp33_ASAP7_75t_R g4065 ( 
.A(n_3923),
.B(n_67),
.Y(n_4065)
);

NOR2xp33_ASAP7_75t_R g4066 ( 
.A(n_3923),
.B(n_67),
.Y(n_4066)
);

NOR2xp33_ASAP7_75t_L g4067 ( 
.A(n_3913),
.B(n_68),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_3906),
.B(n_69),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_3906),
.B(n_70),
.Y(n_4069)
);

BUFx3_ASAP7_75t_L g4070 ( 
.A(n_3931),
.Y(n_4070)
);

INVx2_ASAP7_75t_SL g4071 ( 
.A(n_3969),
.Y(n_4071)
);

NAND2xp33_ASAP7_75t_R g4072 ( 
.A(n_3923),
.B(n_71),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3917),
.Y(n_4073)
);

AND2x2_ASAP7_75t_L g4074 ( 
.A(n_3960),
.B(n_70),
.Y(n_4074)
);

XNOR2xp5_ASAP7_75t_L g4075 ( 
.A(n_3931),
.B(n_71),
.Y(n_4075)
);

NOR2xp33_ASAP7_75t_R g4076 ( 
.A(n_3923),
.B(n_73),
.Y(n_4076)
);

NOR2xp33_ASAP7_75t_R g4077 ( 
.A(n_3923),
.B(n_73),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_L g4078 ( 
.A(n_3906),
.B(n_74),
.Y(n_4078)
);

XNOR2xp5_ASAP7_75t_L g4079 ( 
.A(n_3931),
.B(n_74),
.Y(n_4079)
);

NAND2xp33_ASAP7_75t_R g4080 ( 
.A(n_3923),
.B(n_76),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_3906),
.B(n_75),
.Y(n_4081)
);

AND2x2_ASAP7_75t_L g4082 ( 
.A(n_3960),
.B(n_75),
.Y(n_4082)
);

NOR2xp33_ASAP7_75t_R g4083 ( 
.A(n_3923),
.B(n_76),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3906),
.B(n_77),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_3917),
.Y(n_4085)
);

NAND2xp33_ASAP7_75t_SL g4086 ( 
.A(n_3969),
.B(n_78),
.Y(n_4086)
);

BUFx10_ASAP7_75t_L g4087 ( 
.A(n_3927),
.Y(n_4087)
);

NOR2xp33_ASAP7_75t_R g4088 ( 
.A(n_3923),
.B(n_78),
.Y(n_4088)
);

AND2x2_ASAP7_75t_L g4089 ( 
.A(n_3977),
.B(n_79),
.Y(n_4089)
);

AOI21xp5_ASAP7_75t_L g4090 ( 
.A1(n_4007),
.A2(n_1915),
.B(n_1897),
.Y(n_4090)
);

CKINVDCx5p33_ASAP7_75t_R g4091 ( 
.A(n_4047),
.Y(n_4091)
);

AND2x2_ASAP7_75t_L g4092 ( 
.A(n_4071),
.B(n_79),
.Y(n_4092)
);

AND2x2_ASAP7_75t_L g4093 ( 
.A(n_3974),
.B(n_80),
.Y(n_4093)
);

OR2x2_ASAP7_75t_L g4094 ( 
.A(n_4051),
.B(n_81),
.Y(n_4094)
);

INVx2_ASAP7_75t_L g4095 ( 
.A(n_3992),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3980),
.Y(n_4096)
);

HB1xp67_ASAP7_75t_L g4097 ( 
.A(n_4055),
.Y(n_4097)
);

AND2x2_ASAP7_75t_L g4098 ( 
.A(n_4056),
.B(n_81),
.Y(n_4098)
);

AND2x4_ASAP7_75t_L g4099 ( 
.A(n_3988),
.B(n_82),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_4004),
.Y(n_4100)
);

OAI211xp5_ASAP7_75t_L g4101 ( 
.A1(n_4086),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_4101)
);

AND2x2_ASAP7_75t_L g4102 ( 
.A(n_3972),
.B(n_83),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_3987),
.B(n_84),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_4063),
.Y(n_4104)
);

NOR2xp33_ASAP7_75t_L g4105 ( 
.A(n_4058),
.B(n_85),
.Y(n_4105)
);

INVxp67_ASAP7_75t_SL g4106 ( 
.A(n_3993),
.Y(n_4106)
);

AND2x2_ASAP7_75t_L g4107 ( 
.A(n_4048),
.B(n_86),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_4073),
.Y(n_4108)
);

OR2x2_ASAP7_75t_L g4109 ( 
.A(n_4085),
.B(n_4068),
.Y(n_4109)
);

INVx3_ASAP7_75t_L g4110 ( 
.A(n_3986),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_3997),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_4012),
.Y(n_4112)
);

AND2x2_ASAP7_75t_L g4113 ( 
.A(n_4059),
.B(n_87),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_4003),
.Y(n_4114)
);

INVx2_ASAP7_75t_L g4115 ( 
.A(n_4011),
.Y(n_4115)
);

BUFx2_ASAP7_75t_L g4116 ( 
.A(n_3991),
.Y(n_4116)
);

AND2x2_ASAP7_75t_L g4117 ( 
.A(n_4074),
.B(n_87),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_4069),
.B(n_88),
.Y(n_4118)
);

OR2x6_ASAP7_75t_L g4119 ( 
.A(n_3991),
.B(n_88),
.Y(n_4119)
);

OAI211xp5_ASAP7_75t_L g4120 ( 
.A1(n_3999),
.A2(n_91),
.B(n_89),
.C(n_90),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_4078),
.Y(n_4121)
);

NAND4xp25_ASAP7_75t_L g4122 ( 
.A(n_3998),
.B(n_93),
.C(n_91),
.D(n_92),
.Y(n_4122)
);

NAND4xp25_ASAP7_75t_L g4123 ( 
.A(n_4042),
.B(n_94),
.C(n_92),
.D(n_93),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_4082),
.B(n_94),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4081),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_4006),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_4084),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3983),
.Y(n_4128)
);

OR2x2_ASAP7_75t_L g4129 ( 
.A(n_3979),
.B(n_95),
.Y(n_4129)
);

AND2x2_ASAP7_75t_L g4130 ( 
.A(n_3973),
.B(n_4041),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_4019),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_4000),
.B(n_95),
.Y(n_4132)
);

AND2x2_ASAP7_75t_L g4133 ( 
.A(n_4046),
.B(n_96),
.Y(n_4133)
);

HB1xp67_ASAP7_75t_L g4134 ( 
.A(n_4014),
.Y(n_4134)
);

CKINVDCx14_ASAP7_75t_R g4135 ( 
.A(n_4039),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_4010),
.Y(n_4136)
);

INVx2_ASAP7_75t_L g4137 ( 
.A(n_3981),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3994),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_4032),
.B(n_3990),
.Y(n_4139)
);

OR2x2_ASAP7_75t_L g4140 ( 
.A(n_4015),
.B(n_98),
.Y(n_4140)
);

AND2x4_ASAP7_75t_L g4141 ( 
.A(n_3995),
.B(n_4057),
.Y(n_4141)
);

BUFx2_ASAP7_75t_L g4142 ( 
.A(n_4060),
.Y(n_4142)
);

OR2x2_ASAP7_75t_L g4143 ( 
.A(n_4015),
.B(n_100),
.Y(n_4143)
);

OR2x2_ASAP7_75t_L g4144 ( 
.A(n_3978),
.B(n_4016),
.Y(n_4144)
);

AND2x2_ASAP7_75t_L g4145 ( 
.A(n_3995),
.B(n_100),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_3978),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_4043),
.Y(n_4147)
);

AND2x2_ASAP7_75t_L g4148 ( 
.A(n_4044),
.B(n_101),
.Y(n_4148)
);

OR2x6_ASAP7_75t_L g4149 ( 
.A(n_3975),
.B(n_101),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_4087),
.B(n_102),
.Y(n_4150)
);

HB1xp67_ASAP7_75t_L g4151 ( 
.A(n_3989),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_4064),
.B(n_102),
.Y(n_4152)
);

OR2x2_ASAP7_75t_L g4153 ( 
.A(n_3996),
.B(n_103),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_4036),
.Y(n_4154)
);

INVx3_ASAP7_75t_L g4155 ( 
.A(n_4070),
.Y(n_4155)
);

INVx2_ASAP7_75t_L g4156 ( 
.A(n_4036),
.Y(n_4156)
);

OR2x2_ASAP7_75t_L g4157 ( 
.A(n_3996),
.B(n_103),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_4021),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_4067),
.B(n_104),
.Y(n_4159)
);

OR2x2_ASAP7_75t_L g4160 ( 
.A(n_4030),
.B(n_105),
.Y(n_4160)
);

BUFx8_ASAP7_75t_L g4161 ( 
.A(n_4024),
.Y(n_4161)
);

AOI221xp5_ASAP7_75t_L g4162 ( 
.A1(n_4001),
.A2(n_1974),
.B1(n_1985),
.B2(n_1946),
.C(n_1926),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_4054),
.B(n_105),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4020),
.Y(n_4164)
);

INVx2_ASAP7_75t_SL g4165 ( 
.A(n_4053),
.Y(n_4165)
);

NOR2x1_ASAP7_75t_SL g4166 ( 
.A(n_4024),
.B(n_106),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_4025),
.Y(n_4167)
);

NAND2xp5_ASAP7_75t_L g4168 ( 
.A(n_4022),
.B(n_107),
.Y(n_4168)
);

AND2x2_ASAP7_75t_L g4169 ( 
.A(n_4013),
.B(n_107),
.Y(n_4169)
);

HB1xp67_ASAP7_75t_L g4170 ( 
.A(n_4009),
.Y(n_4170)
);

AO31x2_ASAP7_75t_L g4171 ( 
.A1(n_3982),
.A2(n_110),
.A3(n_108),
.B(n_109),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_4037),
.Y(n_4172)
);

HB1xp67_ASAP7_75t_L g4173 ( 
.A(n_4005),
.Y(n_4173)
);

AND2x2_ASAP7_75t_L g4174 ( 
.A(n_3976),
.B(n_108),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_4008),
.B(n_4034),
.Y(n_4175)
);

AND2x2_ASAP7_75t_L g4176 ( 
.A(n_4075),
.B(n_110),
.Y(n_4176)
);

NOR2xp33_ASAP7_75t_L g4177 ( 
.A(n_4026),
.B(n_111),
.Y(n_4177)
);

AND2x2_ASAP7_75t_L g4178 ( 
.A(n_4079),
.B(n_112),
.Y(n_4178)
);

INVx2_ASAP7_75t_L g4179 ( 
.A(n_4028),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_4018),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_4040),
.B(n_112),
.Y(n_4181)
);

INVx3_ASAP7_75t_L g4182 ( 
.A(n_4045),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3985),
.Y(n_4183)
);

AND2x2_ASAP7_75t_L g4184 ( 
.A(n_4052),
.B(n_113),
.Y(n_4184)
);

AND2x2_ASAP7_75t_L g4185 ( 
.A(n_4061),
.B(n_113),
.Y(n_4185)
);

NOR2xp67_ASAP7_75t_SL g4186 ( 
.A(n_4049),
.B(n_1992),
.Y(n_4186)
);

INVxp33_ASAP7_75t_L g4187 ( 
.A(n_4065),
.Y(n_4187)
);

OR2x2_ASAP7_75t_L g4188 ( 
.A(n_4038),
.B(n_115),
.Y(n_4188)
);

INVx2_ASAP7_75t_L g4189 ( 
.A(n_3984),
.Y(n_4189)
);

INVx3_ASAP7_75t_L g4190 ( 
.A(n_4050),
.Y(n_4190)
);

AND2x2_ASAP7_75t_L g4191 ( 
.A(n_4066),
.B(n_115),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_4029),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4017),
.Y(n_4193)
);

AND2x2_ASAP7_75t_L g4194 ( 
.A(n_4076),
.B(n_116),
.Y(n_4194)
);

AND2x2_ASAP7_75t_L g4195 ( 
.A(n_4077),
.B(n_116),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_4062),
.Y(n_4196)
);

OR2x2_ASAP7_75t_L g4197 ( 
.A(n_4035),
.B(n_117),
.Y(n_4197)
);

AND2x2_ASAP7_75t_L g4198 ( 
.A(n_4083),
.B(n_117),
.Y(n_4198)
);

INVxp67_ASAP7_75t_SL g4199 ( 
.A(n_4072),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_4088),
.B(n_118),
.Y(n_4200)
);

INVx2_ASAP7_75t_L g4201 ( 
.A(n_4080),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4002),
.Y(n_4202)
);

AND2x4_ASAP7_75t_L g4203 ( 
.A(n_4027),
.B(n_118),
.Y(n_4203)
);

HB1xp67_ASAP7_75t_L g4204 ( 
.A(n_4023),
.Y(n_4204)
);

INVx2_ASAP7_75t_L g4205 ( 
.A(n_4033),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4031),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_3977),
.B(n_119),
.Y(n_4207)
);

INVx2_ASAP7_75t_L g4208 ( 
.A(n_3992),
.Y(n_4208)
);

HB1xp67_ASAP7_75t_L g4209 ( 
.A(n_3974),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_3987),
.B(n_119),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_3980),
.Y(n_4211)
);

OR2x2_ASAP7_75t_L g4212 ( 
.A(n_3974),
.B(n_120),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_3987),
.B(n_120),
.Y(n_4213)
);

HB1xp67_ASAP7_75t_L g4214 ( 
.A(n_3974),
.Y(n_4214)
);

BUFx3_ASAP7_75t_L g4215 ( 
.A(n_4058),
.Y(n_4215)
);

AND2x2_ASAP7_75t_L g4216 ( 
.A(n_3977),
.B(n_121),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_3987),
.B(n_121),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_3980),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_3992),
.Y(n_4219)
);

AND2x2_ASAP7_75t_L g4220 ( 
.A(n_3977),
.B(n_122),
.Y(n_4220)
);

HB1xp67_ASAP7_75t_L g4221 ( 
.A(n_3974),
.Y(n_4221)
);

AND2x4_ASAP7_75t_L g4222 ( 
.A(n_4071),
.B(n_122),
.Y(n_4222)
);

INVxp67_ASAP7_75t_L g4223 ( 
.A(n_3982),
.Y(n_4223)
);

AND2x2_ASAP7_75t_L g4224 ( 
.A(n_3977),
.B(n_123),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_3992),
.Y(n_4225)
);

HB1xp67_ASAP7_75t_L g4226 ( 
.A(n_3974),
.Y(n_4226)
);

HB1xp67_ASAP7_75t_L g4227 ( 
.A(n_3974),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_3980),
.Y(n_4228)
);

AND2x2_ASAP7_75t_L g4229 ( 
.A(n_3977),
.B(n_124),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_3980),
.Y(n_4230)
);

OR2x2_ASAP7_75t_L g4231 ( 
.A(n_3974),
.B(n_124),
.Y(n_4231)
);

NOR2xp33_ASAP7_75t_SL g4232 ( 
.A(n_4054),
.B(n_1994),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_3977),
.B(n_125),
.Y(n_4233)
);

AND2x4_ASAP7_75t_L g4234 ( 
.A(n_4071),
.B(n_126),
.Y(n_4234)
);

OR2x2_ASAP7_75t_L g4235 ( 
.A(n_3974),
.B(n_126),
.Y(n_4235)
);

AND2x4_ASAP7_75t_SL g4236 ( 
.A(n_3986),
.B(n_127),
.Y(n_4236)
);

INVx2_ASAP7_75t_SL g4237 ( 
.A(n_3991),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_3980),
.Y(n_4238)
);

AO31x2_ASAP7_75t_L g4239 ( 
.A1(n_4068),
.A2(n_131),
.A3(n_128),
.B(n_129),
.Y(n_4239)
);

INVx3_ASAP7_75t_L g4240 ( 
.A(n_3986),
.Y(n_4240)
);

HB1xp67_ASAP7_75t_L g4241 ( 
.A(n_3974),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_3977),
.B(n_128),
.Y(n_4242)
);

BUFx6f_ASAP7_75t_L g4243 ( 
.A(n_3986),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_3980),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_3980),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_3992),
.Y(n_4246)
);

AND2x2_ASAP7_75t_L g4247 ( 
.A(n_3977),
.B(n_129),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_3980),
.Y(n_4248)
);

AOI22xp33_ASAP7_75t_L g4249 ( 
.A1(n_4170),
.A2(n_2075),
.B1(n_2063),
.B2(n_2003),
.Y(n_4249)
);

HB1xp67_ASAP7_75t_L g4250 ( 
.A(n_4097),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_4156),
.Y(n_4251)
);

AND2x4_ASAP7_75t_SL g4252 ( 
.A(n_4243),
.B(n_131),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_4121),
.B(n_132),
.Y(n_4253)
);

INVxp67_ASAP7_75t_SL g4254 ( 
.A(n_4106),
.Y(n_4254)
);

HB1xp67_ASAP7_75t_L g4255 ( 
.A(n_4209),
.Y(n_4255)
);

BUFx2_ASAP7_75t_L g4256 ( 
.A(n_4110),
.Y(n_4256)
);

AND2x2_ASAP7_75t_L g4257 ( 
.A(n_4147),
.B(n_133),
.Y(n_4257)
);

AND2x2_ASAP7_75t_L g4258 ( 
.A(n_4130),
.B(n_133),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_4146),
.Y(n_4259)
);

INVx2_ASAP7_75t_L g4260 ( 
.A(n_4154),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4096),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4100),
.Y(n_4262)
);

AND2x2_ASAP7_75t_L g4263 ( 
.A(n_4240),
.B(n_134),
.Y(n_4263)
);

HB1xp67_ASAP7_75t_L g4264 ( 
.A(n_4214),
.Y(n_4264)
);

INVx2_ASAP7_75t_L g4265 ( 
.A(n_4189),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_4104),
.Y(n_4266)
);

INVx2_ASAP7_75t_L g4267 ( 
.A(n_4196),
.Y(n_4267)
);

AND2x2_ASAP7_75t_L g4268 ( 
.A(n_4221),
.B(n_136),
.Y(n_4268)
);

INVx2_ASAP7_75t_L g4269 ( 
.A(n_4201),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4108),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4211),
.Y(n_4271)
);

INVxp67_ASAP7_75t_L g4272 ( 
.A(n_4199),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4218),
.Y(n_4273)
);

OAI22xp5_ASAP7_75t_L g4274 ( 
.A1(n_4139),
.A2(n_2004),
.B1(n_2015),
.B2(n_1998),
.Y(n_4274)
);

OR2x2_ASAP7_75t_L g4275 ( 
.A(n_4109),
.B(n_137),
.Y(n_4275)
);

AND2x4_ASAP7_75t_L g4276 ( 
.A(n_4155),
.B(n_138),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_L g4277 ( 
.A(n_4125),
.B(n_4127),
.Y(n_4277)
);

OR2x2_ASAP7_75t_L g4278 ( 
.A(n_4226),
.B(n_139),
.Y(n_4278)
);

NOR2xp33_ASAP7_75t_L g4279 ( 
.A(n_4135),
.B(n_139),
.Y(n_4279)
);

OR2x2_ASAP7_75t_L g4280 ( 
.A(n_4227),
.B(n_140),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4228),
.Y(n_4281)
);

INVx2_ASAP7_75t_L g4282 ( 
.A(n_4151),
.Y(n_4282)
);

AND2x2_ASAP7_75t_L g4283 ( 
.A(n_4241),
.B(n_141),
.Y(n_4283)
);

AND2x2_ASAP7_75t_L g4284 ( 
.A(n_4114),
.B(n_142),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4230),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_4128),
.B(n_142),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_4138),
.B(n_143),
.Y(n_4287)
);

NOR2xp67_ASAP7_75t_L g4288 ( 
.A(n_4182),
.B(n_143),
.Y(n_4288)
);

AND2x2_ASAP7_75t_L g4289 ( 
.A(n_4116),
.B(n_144),
.Y(n_4289)
);

AND2x4_ASAP7_75t_L g4290 ( 
.A(n_4137),
.B(n_144),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4238),
.Y(n_4291)
);

AND2x2_ASAP7_75t_L g4292 ( 
.A(n_4092),
.B(n_145),
.Y(n_4292)
);

AND2x4_ASAP7_75t_L g4293 ( 
.A(n_4141),
.B(n_145),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4244),
.Y(n_4294)
);

BUFx2_ASAP7_75t_L g4295 ( 
.A(n_4243),
.Y(n_4295)
);

AND2x4_ASAP7_75t_L g4296 ( 
.A(n_4237),
.B(n_146),
.Y(n_4296)
);

AND2x4_ASAP7_75t_L g4297 ( 
.A(n_4126),
.B(n_146),
.Y(n_4297)
);

NOR2xp33_ASAP7_75t_L g4298 ( 
.A(n_4187),
.B(n_147),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4245),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4248),
.Y(n_4300)
);

HB1xp67_ASAP7_75t_L g4301 ( 
.A(n_4134),
.Y(n_4301)
);

INVxp67_ASAP7_75t_SL g4302 ( 
.A(n_4190),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4136),
.Y(n_4303)
);

HB1xp67_ASAP7_75t_L g4304 ( 
.A(n_4239),
.Y(n_4304)
);

HB1xp67_ASAP7_75t_L g4305 ( 
.A(n_4239),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4094),
.Y(n_4306)
);

OR2x2_ASAP7_75t_L g4307 ( 
.A(n_4129),
.B(n_147),
.Y(n_4307)
);

AND2x4_ASAP7_75t_L g4308 ( 
.A(n_4142),
.B(n_148),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_4222),
.B(n_149),
.Y(n_4309)
);

INVx2_ASAP7_75t_L g4310 ( 
.A(n_4172),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4167),
.B(n_4089),
.Y(n_4311)
);

AND2x2_ASAP7_75t_L g4312 ( 
.A(n_4234),
.B(n_149),
.Y(n_4312)
);

AND2x4_ASAP7_75t_L g4313 ( 
.A(n_4215),
.B(n_150),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_4212),
.Y(n_4314)
);

BUFx3_ASAP7_75t_L g4315 ( 
.A(n_4236),
.Y(n_4315)
);

INVx2_ASAP7_75t_L g4316 ( 
.A(n_4173),
.Y(n_4316)
);

NOR2xp67_ASAP7_75t_SL g4317 ( 
.A(n_4140),
.B(n_2029),
.Y(n_4317)
);

OR2x2_ASAP7_75t_L g4318 ( 
.A(n_4231),
.B(n_151),
.Y(n_4318)
);

HB1xp67_ASAP7_75t_L g4319 ( 
.A(n_4235),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_4158),
.Y(n_4320)
);

AND2x2_ASAP7_75t_L g4321 ( 
.A(n_4093),
.B(n_151),
.Y(n_4321)
);

AND2x2_ASAP7_75t_L g4322 ( 
.A(n_4098),
.B(n_152),
.Y(n_4322)
);

OR2x2_ASAP7_75t_SL g4323 ( 
.A(n_4144),
.B(n_152),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4207),
.B(n_4216),
.Y(n_4324)
);

INVx2_ASAP7_75t_L g4325 ( 
.A(n_4192),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4103),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_4220),
.B(n_153),
.Y(n_4327)
);

AND2x2_ASAP7_75t_L g4328 ( 
.A(n_4224),
.B(n_153),
.Y(n_4328)
);

OR2x2_ASAP7_75t_L g4329 ( 
.A(n_4131),
.B(n_154),
.Y(n_4329)
);

AND2x4_ASAP7_75t_L g4330 ( 
.A(n_4099),
.B(n_154),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4210),
.Y(n_4331)
);

BUFx2_ASAP7_75t_L g4332 ( 
.A(n_4119),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4213),
.Y(n_4333)
);

AND2x2_ASAP7_75t_L g4334 ( 
.A(n_4229),
.B(n_155),
.Y(n_4334)
);

AND2x2_ASAP7_75t_L g4335 ( 
.A(n_4233),
.B(n_4242),
.Y(n_4335)
);

INVx2_ASAP7_75t_L g4336 ( 
.A(n_4171),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4247),
.B(n_155),
.Y(n_4337)
);

AND2x2_ASAP7_75t_L g4338 ( 
.A(n_4102),
.B(n_156),
.Y(n_4338)
);

NOR2xp33_ASAP7_75t_L g4339 ( 
.A(n_4223),
.B(n_158),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4217),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4115),
.Y(n_4341)
);

AND2x2_ASAP7_75t_L g4342 ( 
.A(n_4107),
.B(n_4113),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_4117),
.B(n_159),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_4124),
.B(n_160),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4164),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4118),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4179),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_4133),
.B(n_161),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_SL g4349 ( 
.A(n_4160),
.B(n_2049),
.Y(n_4349)
);

INVx2_ASAP7_75t_L g4350 ( 
.A(n_4171),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_4165),
.B(n_161),
.Y(n_4351)
);

OR2x2_ASAP7_75t_L g4352 ( 
.A(n_4132),
.B(n_164),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_4169),
.B(n_165),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4095),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_4119),
.B(n_165),
.Y(n_4355)
);

INVxp67_ASAP7_75t_L g4356 ( 
.A(n_4204),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4111),
.Y(n_4357)
);

AND2x6_ASAP7_75t_L g4358 ( 
.A(n_4184),
.B(n_166),
.Y(n_4358)
);

INVx2_ASAP7_75t_L g4359 ( 
.A(n_4112),
.Y(n_4359)
);

AND2x4_ASAP7_75t_L g4360 ( 
.A(n_4148),
.B(n_168),
.Y(n_4360)
);

INVx2_ASAP7_75t_SL g4361 ( 
.A(n_4091),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4208),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_4150),
.B(n_168),
.Y(n_4363)
);

AND2x4_ASAP7_75t_L g4364 ( 
.A(n_4152),
.B(n_169),
.Y(n_4364)
);

OR2x2_ASAP7_75t_L g4365 ( 
.A(n_4246),
.B(n_170),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4219),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4225),
.Y(n_4367)
);

INVx2_ASAP7_75t_L g4368 ( 
.A(n_4153),
.Y(n_4368)
);

AND2x2_ASAP7_75t_L g4369 ( 
.A(n_4159),
.B(n_171),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4143),
.Y(n_4370)
);

AND2x2_ASAP7_75t_L g4371 ( 
.A(n_4145),
.B(n_172),
.Y(n_4371)
);

AND2x2_ASAP7_75t_L g4372 ( 
.A(n_4149),
.B(n_172),
.Y(n_4372)
);

AND2x2_ASAP7_75t_L g4373 ( 
.A(n_4149),
.B(n_173),
.Y(n_4373)
);

BUFx2_ASAP7_75t_L g4374 ( 
.A(n_4163),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4168),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4157),
.Y(n_4376)
);

AND2x4_ASAP7_75t_L g4377 ( 
.A(n_4183),
.B(n_173),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_4185),
.B(n_174),
.Y(n_4378)
);

INVx2_ASAP7_75t_L g4379 ( 
.A(n_4161),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4197),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_4193),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4180),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4175),
.Y(n_4383)
);

BUFx2_ASAP7_75t_L g4384 ( 
.A(n_4191),
.Y(n_4384)
);

AND2x2_ASAP7_75t_L g4385 ( 
.A(n_4105),
.B(n_174),
.Y(n_4385)
);

BUFx2_ASAP7_75t_L g4386 ( 
.A(n_4194),
.Y(n_4386)
);

INVxp67_ASAP7_75t_SL g4387 ( 
.A(n_4181),
.Y(n_4387)
);

INVx2_ASAP7_75t_L g4388 ( 
.A(n_4202),
.Y(n_4388)
);

INVx2_ASAP7_75t_L g4389 ( 
.A(n_4206),
.Y(n_4389)
);

HB1xp67_ASAP7_75t_L g4390 ( 
.A(n_4188),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4205),
.Y(n_4391)
);

INVx2_ASAP7_75t_L g4392 ( 
.A(n_4166),
.Y(n_4392)
);

AND2x2_ASAP7_75t_L g4393 ( 
.A(n_4174),
.B(n_175),
.Y(n_4393)
);

NOR2x1_ASAP7_75t_SL g4394 ( 
.A(n_4101),
.B(n_175),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4195),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4198),
.Y(n_4396)
);

INVx2_ASAP7_75t_L g4397 ( 
.A(n_4203),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_4200),
.B(n_176),
.Y(n_4398)
);

INVx2_ASAP7_75t_L g4399 ( 
.A(n_4176),
.Y(n_4399)
);

AND2x2_ASAP7_75t_L g4400 ( 
.A(n_4178),
.B(n_177),
.Y(n_4400)
);

INVx2_ASAP7_75t_L g4401 ( 
.A(n_4177),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4123),
.Y(n_4402)
);

AND2x2_ASAP7_75t_L g4403 ( 
.A(n_4232),
.B(n_177),
.Y(n_4403)
);

AND2x2_ASAP7_75t_L g4404 ( 
.A(n_4186),
.B(n_178),
.Y(n_4404)
);

INVxp67_ASAP7_75t_L g4405 ( 
.A(n_4122),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_4120),
.B(n_178),
.Y(n_4406)
);

CKINVDCx5p33_ASAP7_75t_R g4407 ( 
.A(n_4090),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4162),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4096),
.Y(n_4409)
);

BUFx2_ASAP7_75t_L g4410 ( 
.A(n_4110),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_L g4411 ( 
.A(n_4121),
.B(n_180),
.Y(n_4411)
);

INVx2_ASAP7_75t_L g4412 ( 
.A(n_4156),
.Y(n_4412)
);

AND2x2_ASAP7_75t_L g4413 ( 
.A(n_4106),
.B(n_180),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4106),
.B(n_181),
.Y(n_4414)
);

INVx2_ASAP7_75t_L g4415 ( 
.A(n_4156),
.Y(n_4415)
);

NAND2xp5_ASAP7_75t_L g4416 ( 
.A(n_4121),
.B(n_181),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4096),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4096),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_SL g4419 ( 
.A(n_4139),
.B(n_2057),
.Y(n_4419)
);

AND2x2_ASAP7_75t_L g4420 ( 
.A(n_4106),
.B(n_182),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4096),
.Y(n_4421)
);

INVx3_ASAP7_75t_L g4422 ( 
.A(n_4243),
.Y(n_4422)
);

NAND2xp5_ASAP7_75t_L g4423 ( 
.A(n_4121),
.B(n_183),
.Y(n_4423)
);

AND2x2_ASAP7_75t_L g4424 ( 
.A(n_4106),
.B(n_183),
.Y(n_4424)
);

HB1xp67_ASAP7_75t_L g4425 ( 
.A(n_4097),
.Y(n_4425)
);

HB1xp67_ASAP7_75t_L g4426 ( 
.A(n_4097),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4096),
.Y(n_4427)
);

INVx2_ASAP7_75t_L g4428 ( 
.A(n_4156),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_4121),
.B(n_184),
.Y(n_4429)
);

HB1xp67_ASAP7_75t_L g4430 ( 
.A(n_4097),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_L g4431 ( 
.A(n_4121),
.B(n_184),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4106),
.B(n_185),
.Y(n_4432)
);

NOR2x1_ASAP7_75t_L g4433 ( 
.A(n_4155),
.B(n_185),
.Y(n_4433)
);

OR2x2_ASAP7_75t_L g4434 ( 
.A(n_4109),
.B(n_186),
.Y(n_4434)
);

AND2x2_ASAP7_75t_L g4435 ( 
.A(n_4106),
.B(n_186),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4096),
.Y(n_4436)
);

BUFx2_ASAP7_75t_L g4437 ( 
.A(n_4110),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_4096),
.Y(n_4438)
);

NOR2x1_ASAP7_75t_SL g4439 ( 
.A(n_4149),
.B(n_187),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_L g4440 ( 
.A(n_4121),
.B(n_188),
.Y(n_4440)
);

INVx2_ASAP7_75t_L g4441 ( 
.A(n_4156),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4096),
.Y(n_4442)
);

AND2x2_ASAP7_75t_L g4443 ( 
.A(n_4256),
.B(n_189),
.Y(n_4443)
);

AND2x2_ASAP7_75t_L g4444 ( 
.A(n_4410),
.B(n_189),
.Y(n_4444)
);

NAND2xp5_ASAP7_75t_L g4445 ( 
.A(n_4390),
.B(n_190),
.Y(n_4445)
);

AND2x2_ASAP7_75t_L g4446 ( 
.A(n_4437),
.B(n_190),
.Y(n_4446)
);

INVx2_ASAP7_75t_L g4447 ( 
.A(n_4342),
.Y(n_4447)
);

BUFx2_ASAP7_75t_L g4448 ( 
.A(n_4295),
.Y(n_4448)
);

OR2x2_ASAP7_75t_L g4449 ( 
.A(n_4301),
.B(n_192),
.Y(n_4449)
);

INVx3_ASAP7_75t_L g4450 ( 
.A(n_4315),
.Y(n_4450)
);

OR2x2_ASAP7_75t_L g4451 ( 
.A(n_4282),
.B(n_193),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_4250),
.Y(n_4452)
);

AND2x4_ASAP7_75t_L g4453 ( 
.A(n_4379),
.B(n_194),
.Y(n_4453)
);

BUFx2_ASAP7_75t_L g4454 ( 
.A(n_4422),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4255),
.Y(n_4455)
);

AND2x2_ASAP7_75t_L g4456 ( 
.A(n_4254),
.B(n_194),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4264),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_4332),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_4374),
.B(n_195),
.Y(n_4459)
);

HB1xp67_ASAP7_75t_L g4460 ( 
.A(n_4272),
.Y(n_4460)
);

AND2x2_ASAP7_75t_L g4461 ( 
.A(n_4413),
.B(n_195),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_R g4462 ( 
.A(n_4361),
.B(n_196),
.Y(n_4462)
);

HB1xp67_ASAP7_75t_L g4463 ( 
.A(n_4316),
.Y(n_4463)
);

AOI22xp33_ASAP7_75t_L g4464 ( 
.A1(n_4265),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_4464)
);

OR2x2_ASAP7_75t_L g4465 ( 
.A(n_4425),
.B(n_197),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4426),
.Y(n_4466)
);

HB1xp67_ASAP7_75t_L g4467 ( 
.A(n_4430),
.Y(n_4467)
);

OR2x2_ASAP7_75t_L g4468 ( 
.A(n_4383),
.B(n_198),
.Y(n_4468)
);

INVx1_ASAP7_75t_L g4469 ( 
.A(n_4277),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4382),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_L g4471 ( 
.A(n_4414),
.B(n_199),
.Y(n_4471)
);

AND2x2_ASAP7_75t_L g4472 ( 
.A(n_4420),
.B(n_200),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4261),
.Y(n_4473)
);

NOR2xp33_ASAP7_75t_L g4474 ( 
.A(n_4405),
.B(n_200),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4262),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_4424),
.B(n_201),
.Y(n_4476)
);

INVx2_ASAP7_75t_L g4477 ( 
.A(n_4324),
.Y(n_4477)
);

AND2x2_ASAP7_75t_L g4478 ( 
.A(n_4432),
.B(n_201),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_4435),
.B(n_202),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4266),
.Y(n_4480)
);

AND2x4_ASAP7_75t_L g4481 ( 
.A(n_4302),
.B(n_202),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_4399),
.B(n_4384),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4270),
.Y(n_4483)
);

OR2x2_ASAP7_75t_L g4484 ( 
.A(n_4346),
.B(n_203),
.Y(n_4484)
);

HB1xp67_ASAP7_75t_L g4485 ( 
.A(n_4356),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_4335),
.Y(n_4486)
);

OR2x6_ASAP7_75t_SL g4487 ( 
.A(n_4381),
.B(n_203),
.Y(n_4487)
);

AND2x4_ASAP7_75t_L g4488 ( 
.A(n_4258),
.B(n_204),
.Y(n_4488)
);

NOR2xp33_ASAP7_75t_L g4489 ( 
.A(n_4275),
.B(n_205),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4257),
.B(n_206),
.Y(n_4490)
);

AND2x4_ASAP7_75t_L g4491 ( 
.A(n_4388),
.B(n_208),
.Y(n_4491)
);

AND2x2_ASAP7_75t_L g4492 ( 
.A(n_4268),
.B(n_4283),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4271),
.Y(n_4493)
);

AND2x2_ASAP7_75t_L g4494 ( 
.A(n_4289),
.B(n_208),
.Y(n_4494)
);

AND2x2_ASAP7_75t_L g4495 ( 
.A(n_4319),
.B(n_4389),
.Y(n_4495)
);

OR2x2_ASAP7_75t_L g4496 ( 
.A(n_4306),
.B(n_209),
.Y(n_4496)
);

OR2x2_ASAP7_75t_L g4497 ( 
.A(n_4314),
.B(n_210),
.Y(n_4497)
);

AND2x2_ASAP7_75t_L g4498 ( 
.A(n_4263),
.B(n_210),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4273),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_4281),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4296),
.B(n_211),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_4386),
.B(n_211),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4285),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4291),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4294),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4299),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4300),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_4387),
.B(n_4395),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4303),
.B(n_212),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4409),
.Y(n_4510)
);

BUFx2_ASAP7_75t_L g4511 ( 
.A(n_4433),
.Y(n_4511)
);

AND2x2_ASAP7_75t_L g4512 ( 
.A(n_4345),
.B(n_213),
.Y(n_4512)
);

INVxp67_ASAP7_75t_SL g4513 ( 
.A(n_4439),
.Y(n_4513)
);

INVx4_ASAP7_75t_L g4514 ( 
.A(n_4313),
.Y(n_4514)
);

OR2x2_ASAP7_75t_L g4515 ( 
.A(n_4434),
.B(n_213),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_L g4516 ( 
.A(n_4396),
.B(n_4370),
.Y(n_4516)
);

AND2x4_ASAP7_75t_L g4517 ( 
.A(n_4364),
.B(n_214),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4417),
.Y(n_4518)
);

AND2x2_ASAP7_75t_L g4519 ( 
.A(n_4402),
.B(n_215),
.Y(n_4519)
);

AND2x2_ASAP7_75t_L g4520 ( 
.A(n_4351),
.B(n_215),
.Y(n_4520)
);

INVx3_ASAP7_75t_L g4521 ( 
.A(n_4308),
.Y(n_4521)
);

OR2x2_ASAP7_75t_L g4522 ( 
.A(n_4326),
.B(n_218),
.Y(n_4522)
);

OR2x2_ASAP7_75t_L g4523 ( 
.A(n_4331),
.B(n_218),
.Y(n_4523)
);

INVxp67_ASAP7_75t_SL g4524 ( 
.A(n_4394),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_4418),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4421),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4323),
.Y(n_4527)
);

INVx1_ASAP7_75t_L g4528 ( 
.A(n_4427),
.Y(n_4528)
);

NAND4xp25_ASAP7_75t_L g4529 ( 
.A(n_4249),
.B(n_222),
.C(n_219),
.D(n_220),
.Y(n_4529)
);

INVx2_ASAP7_75t_L g4530 ( 
.A(n_4365),
.Y(n_4530)
);

AND2x2_ASAP7_75t_L g4531 ( 
.A(n_4376),
.B(n_219),
.Y(n_4531)
);

AND2x4_ASAP7_75t_L g4532 ( 
.A(n_4397),
.B(n_222),
.Y(n_4532)
);

AOI22xp33_ASAP7_75t_L g4533 ( 
.A1(n_4325),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_4533)
);

AND2x2_ASAP7_75t_L g4534 ( 
.A(n_4276),
.B(n_227),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4436),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4438),
.Y(n_4536)
);

OR2x2_ASAP7_75t_L g4537 ( 
.A(n_4333),
.B(n_228),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4442),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4278),
.Y(n_4539)
);

INVx2_ASAP7_75t_L g4540 ( 
.A(n_4310),
.Y(n_4540)
);

AND2x2_ASAP7_75t_L g4541 ( 
.A(n_4293),
.B(n_228),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_L g4542 ( 
.A(n_4284),
.B(n_229),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_4392),
.Y(n_4543)
);

INVxp67_ASAP7_75t_L g4544 ( 
.A(n_4358),
.Y(n_4544)
);

INVx1_ASAP7_75t_L g4545 ( 
.A(n_4280),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4368),
.B(n_229),
.Y(n_4546)
);

HB1xp67_ASAP7_75t_L g4547 ( 
.A(n_4391),
.Y(n_4547)
);

INVx2_ASAP7_75t_L g4548 ( 
.A(n_4329),
.Y(n_4548)
);

AND2x2_ASAP7_75t_L g4549 ( 
.A(n_4340),
.B(n_230),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4341),
.Y(n_4550)
);

INVx3_ASAP7_75t_L g4551 ( 
.A(n_4377),
.Y(n_4551)
);

BUFx2_ASAP7_75t_L g4552 ( 
.A(n_4287),
.Y(n_4552)
);

BUFx2_ASAP7_75t_L g4553 ( 
.A(n_4385),
.Y(n_4553)
);

INVx2_ASAP7_75t_L g4554 ( 
.A(n_4267),
.Y(n_4554)
);

HB1xp67_ASAP7_75t_L g4555 ( 
.A(n_4311),
.Y(n_4555)
);

AND2x4_ASAP7_75t_SL g4556 ( 
.A(n_4330),
.B(n_230),
.Y(n_4556)
);

AND2x2_ASAP7_75t_L g4557 ( 
.A(n_4321),
.B(n_231),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4304),
.Y(n_4558)
);

BUFx2_ASAP7_75t_L g4559 ( 
.A(n_4286),
.Y(n_4559)
);

INVx2_ASAP7_75t_L g4560 ( 
.A(n_4269),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_4305),
.Y(n_4561)
);

AND2x2_ASAP7_75t_L g4562 ( 
.A(n_4322),
.B(n_231),
.Y(n_4562)
);

OR2x2_ASAP7_75t_L g4563 ( 
.A(n_4253),
.B(n_232),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4347),
.Y(n_4564)
);

AND2x2_ASAP7_75t_L g4565 ( 
.A(n_4292),
.B(n_233),
.Y(n_4565)
);

AND2x2_ASAP7_75t_L g4566 ( 
.A(n_4369),
.B(n_234),
.Y(n_4566)
);

AND2x4_ASAP7_75t_L g4567 ( 
.A(n_4338),
.B(n_234),
.Y(n_4567)
);

NAND2xp5_ASAP7_75t_L g4568 ( 
.A(n_4375),
.B(n_235),
.Y(n_4568)
);

OR2x2_ASAP7_75t_L g4569 ( 
.A(n_4411),
.B(n_235),
.Y(n_4569)
);

INVx4_ASAP7_75t_L g4570 ( 
.A(n_4252),
.Y(n_4570)
);

AND2x2_ASAP7_75t_L g4571 ( 
.A(n_4348),
.B(n_4344),
.Y(n_4571)
);

NOR2xp33_ASAP7_75t_L g4572 ( 
.A(n_4279),
.B(n_237),
.Y(n_4572)
);

INVx2_ASAP7_75t_L g4573 ( 
.A(n_4259),
.Y(n_4573)
);

AND2x4_ASAP7_75t_L g4574 ( 
.A(n_4371),
.B(n_237),
.Y(n_4574)
);

AND2x2_ASAP7_75t_L g4575 ( 
.A(n_4309),
.B(n_238),
.Y(n_4575)
);

NAND2x1p5_ASAP7_75t_L g4576 ( 
.A(n_4288),
.B(n_239),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_L g4577 ( 
.A(n_4380),
.B(n_240),
.Y(n_4577)
);

AND2x2_ASAP7_75t_L g4578 ( 
.A(n_4312),
.B(n_241),
.Y(n_4578)
);

INVx2_ASAP7_75t_L g4579 ( 
.A(n_4360),
.Y(n_4579)
);

AND2x4_ASAP7_75t_L g4580 ( 
.A(n_4570),
.B(n_4372),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4467),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4485),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4460),
.Y(n_4583)
);

AND2x2_ASAP7_75t_L g4584 ( 
.A(n_4513),
.B(n_4355),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4553),
.B(n_4401),
.Y(n_4585)
);

INVx3_ASAP7_75t_L g4586 ( 
.A(n_4514),
.Y(n_4586)
);

OAI21xp5_ASAP7_75t_L g4587 ( 
.A1(n_4524),
.A2(n_4406),
.B(n_4339),
.Y(n_4587)
);

AND2x4_ASAP7_75t_L g4588 ( 
.A(n_4450),
.B(n_4571),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_4448),
.B(n_4260),
.Y(n_4589)
);

INVxp67_ASAP7_75t_SL g4590 ( 
.A(n_4511),
.Y(n_4590)
);

AND2x2_ASAP7_75t_L g4591 ( 
.A(n_4454),
.B(n_4373),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4558),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4561),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4445),
.Y(n_4594)
);

AND2x2_ASAP7_75t_L g4595 ( 
.A(n_4492),
.B(n_4328),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_L g4596 ( 
.A(n_4559),
.B(n_4334),
.Y(n_4596)
);

AND2x2_ASAP7_75t_L g4597 ( 
.A(n_4447),
.B(n_4337),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_4456),
.B(n_4393),
.Y(n_4598)
);

AND2x2_ASAP7_75t_L g4599 ( 
.A(n_4477),
.B(n_4486),
.Y(n_4599)
);

BUFx2_ASAP7_75t_L g4600 ( 
.A(n_4521),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4459),
.Y(n_4601)
);

AND2x2_ASAP7_75t_L g4602 ( 
.A(n_4555),
.B(n_4298),
.Y(n_4602)
);

AND2x4_ASAP7_75t_L g4603 ( 
.A(n_4551),
.B(n_4363),
.Y(n_4603)
);

AND2x2_ASAP7_75t_L g4604 ( 
.A(n_4495),
.B(n_4416),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_4576),
.Y(n_4605)
);

AND2x2_ASAP7_75t_L g4606 ( 
.A(n_4458),
.B(n_4443),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4465),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4552),
.B(n_4400),
.Y(n_4608)
);

OR2x2_ASAP7_75t_L g4609 ( 
.A(n_4482),
.B(n_4423),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_4548),
.B(n_4549),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_4444),
.B(n_4429),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_4446),
.B(n_4463),
.Y(n_4612)
);

AND2x2_ASAP7_75t_L g4613 ( 
.A(n_4481),
.B(n_4431),
.Y(n_4613)
);

NAND4xp25_ASAP7_75t_L g4614 ( 
.A(n_4452),
.B(n_4440),
.C(n_4343),
.D(n_4274),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4449),
.Y(n_4615)
);

AND2x2_ASAP7_75t_SL g4616 ( 
.A(n_4527),
.B(n_4297),
.Y(n_4616)
);

NOR2xp33_ASAP7_75t_L g4617 ( 
.A(n_4487),
.B(n_4349),
.Y(n_4617)
);

NAND2x1p5_ASAP7_75t_L g4618 ( 
.A(n_4574),
.B(n_4317),
.Y(n_4618)
);

AND2x4_ASAP7_75t_SL g4619 ( 
.A(n_4453),
.B(n_4290),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_L g4620 ( 
.A(n_4531),
.B(n_4358),
.Y(n_4620)
);

OR2x2_ASAP7_75t_L g4621 ( 
.A(n_4516),
.B(n_4318),
.Y(n_4621)
);

AND2x4_ASAP7_75t_SL g4622 ( 
.A(n_4488),
.B(n_4403),
.Y(n_4622)
);

INVx2_ASAP7_75t_L g4623 ( 
.A(n_4515),
.Y(n_4623)
);

HB1xp67_ASAP7_75t_L g4624 ( 
.A(n_4547),
.Y(n_4624)
);

AND2x2_ASAP7_75t_L g4625 ( 
.A(n_4509),
.B(n_4419),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4508),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_4539),
.B(n_4358),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4455),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_L g4629 ( 
.A(n_4545),
.B(n_4408),
.Y(n_4629)
);

INVx2_ASAP7_75t_L g4630 ( 
.A(n_4491),
.Y(n_4630)
);

OR2x2_ASAP7_75t_L g4631 ( 
.A(n_4457),
.B(n_4307),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4466),
.Y(n_4632)
);

AND2x2_ASAP7_75t_L g4633 ( 
.A(n_4470),
.B(n_4412),
.Y(n_4633)
);

INVx1_ASAP7_75t_SL g4634 ( 
.A(n_4556),
.Y(n_4634)
);

OR2x2_ASAP7_75t_L g4635 ( 
.A(n_4502),
.B(n_4352),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4519),
.Y(n_4636)
);

AND2x2_ASAP7_75t_L g4637 ( 
.A(n_4512),
.B(n_4415),
.Y(n_4637)
);

AND2x2_ASAP7_75t_L g4638 ( 
.A(n_4469),
.B(n_4428),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4489),
.B(n_4327),
.Y(n_4639)
);

AND2x2_ASAP7_75t_L g4640 ( 
.A(n_4494),
.B(n_4441),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4496),
.Y(n_4641)
);

AND2x4_ASAP7_75t_L g4642 ( 
.A(n_4567),
.B(n_4320),
.Y(n_4642)
);

AND2x2_ASAP7_75t_L g4643 ( 
.A(n_4520),
.B(n_4251),
.Y(n_4643)
);

OR2x2_ASAP7_75t_L g4644 ( 
.A(n_4568),
.B(n_4378),
.Y(n_4644)
);

INVx2_ASAP7_75t_L g4645 ( 
.A(n_4451),
.Y(n_4645)
);

AND2x2_ASAP7_75t_L g4646 ( 
.A(n_4490),
.B(n_4407),
.Y(n_4646)
);

INVxp67_ASAP7_75t_L g4647 ( 
.A(n_4572),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_L g4648 ( 
.A(n_4461),
.B(n_4336),
.Y(n_4648)
);

INVx2_ASAP7_75t_L g4649 ( 
.A(n_4579),
.Y(n_4649)
);

AND2x2_ASAP7_75t_L g4650 ( 
.A(n_4474),
.B(n_4353),
.Y(n_4650)
);

AND2x2_ASAP7_75t_L g4651 ( 
.A(n_4472),
.B(n_4398),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_4476),
.B(n_4478),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4498),
.B(n_4404),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4497),
.Y(n_4654)
);

HB1xp67_ASAP7_75t_L g4655 ( 
.A(n_4577),
.Y(n_4655)
);

AND2x2_ASAP7_75t_L g4656 ( 
.A(n_4501),
.B(n_4350),
.Y(n_4656)
);

NAND2xp5_ASAP7_75t_SL g4657 ( 
.A(n_4468),
.B(n_4359),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4564),
.Y(n_4658)
);

NAND2xp5_ASAP7_75t_L g4659 ( 
.A(n_4484),
.B(n_4354),
.Y(n_4659)
);

INVx1_ASAP7_75t_SL g4660 ( 
.A(n_4566),
.Y(n_4660)
);

NAND2xp5_ASAP7_75t_SL g4661 ( 
.A(n_4522),
.B(n_4357),
.Y(n_4661)
);

OR2x2_ASAP7_75t_L g4662 ( 
.A(n_4546),
.B(n_4366),
.Y(n_4662)
);

AND2x2_ASAP7_75t_L g4663 ( 
.A(n_4473),
.B(n_4362),
.Y(n_4663)
);

AND2x4_ASAP7_75t_L g4664 ( 
.A(n_4575),
.B(n_4578),
.Y(n_4664)
);

AND2x4_ASAP7_75t_L g4665 ( 
.A(n_4557),
.B(n_4367),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4475),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_4480),
.Y(n_4667)
);

AND2x4_ASAP7_75t_L g4668 ( 
.A(n_4562),
.B(n_242),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4483),
.Y(n_4669)
);

AND2x2_ASAP7_75t_L g4670 ( 
.A(n_4493),
.B(n_4499),
.Y(n_4670)
);

INVx2_ASAP7_75t_L g4671 ( 
.A(n_4532),
.Y(n_4671)
);

OR2x2_ASAP7_75t_L g4672 ( 
.A(n_4550),
.B(n_243),
.Y(n_4672)
);

OR2x2_ASAP7_75t_L g4673 ( 
.A(n_4608),
.B(n_4585),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4624),
.Y(n_4674)
);

XOR2xp5_ASAP7_75t_L g4675 ( 
.A(n_4664),
.B(n_4517),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4655),
.Y(n_4676)
);

INVx3_ASAP7_75t_L g4677 ( 
.A(n_4588),
.Y(n_4677)
);

OR2x2_ASAP7_75t_L g4678 ( 
.A(n_4596),
.B(n_4500),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4581),
.Y(n_4679)
);

OR2x2_ASAP7_75t_L g4680 ( 
.A(n_4590),
.B(n_4503),
.Y(n_4680)
);

NOR2xp33_ASAP7_75t_SL g4681 ( 
.A(n_4660),
.B(n_4544),
.Y(n_4681)
);

AND2x2_ASAP7_75t_L g4682 ( 
.A(n_4591),
.B(n_4504),
.Y(n_4682)
);

AND2x2_ASAP7_75t_L g4683 ( 
.A(n_4595),
.B(n_4505),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_4600),
.B(n_4506),
.Y(n_4684)
);

AND2x2_ASAP7_75t_L g4685 ( 
.A(n_4584),
.B(n_4580),
.Y(n_4685)
);

INVx2_ASAP7_75t_L g4686 ( 
.A(n_4652),
.Y(n_4686)
);

INVx2_ASAP7_75t_L g4687 ( 
.A(n_4616),
.Y(n_4687)
);

AND2x4_ASAP7_75t_L g4688 ( 
.A(n_4603),
.B(n_4534),
.Y(n_4688)
);

OR2x2_ASAP7_75t_L g4689 ( 
.A(n_4621),
.B(n_4507),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_L g4690 ( 
.A(n_4651),
.B(n_4523),
.Y(n_4690)
);

INVxp67_ASAP7_75t_L g4691 ( 
.A(n_4612),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4582),
.Y(n_4692)
);

HB1xp67_ASAP7_75t_L g4693 ( 
.A(n_4598),
.Y(n_4693)
);

OAI21xp5_ASAP7_75t_SL g4694 ( 
.A1(n_4606),
.A2(n_4518),
.B(n_4510),
.Y(n_4694)
);

HB1xp67_ASAP7_75t_L g4695 ( 
.A(n_4597),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_4602),
.B(n_4537),
.Y(n_4696)
);

AND2x4_ASAP7_75t_L g4697 ( 
.A(n_4586),
.B(n_4541),
.Y(n_4697)
);

AND2x2_ASAP7_75t_L g4698 ( 
.A(n_4589),
.B(n_4525),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_L g4699 ( 
.A(n_4601),
.B(n_4565),
.Y(n_4699)
);

AND2x2_ASAP7_75t_L g4700 ( 
.A(n_4599),
.B(n_4526),
.Y(n_4700)
);

INVx1_ASAP7_75t_SL g4701 ( 
.A(n_4646),
.Y(n_4701)
);

AND2x2_ASAP7_75t_L g4702 ( 
.A(n_4634),
.B(n_4528),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4583),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_4604),
.B(n_4535),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4613),
.B(n_4536),
.Y(n_4705)
);

AND2x2_ASAP7_75t_L g4706 ( 
.A(n_4611),
.B(n_4538),
.Y(n_4706)
);

AND2x2_ASAP7_75t_L g4707 ( 
.A(n_4626),
.B(n_4471),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_4640),
.B(n_4540),
.Y(n_4708)
);

OAI22xp5_ASAP7_75t_L g4709 ( 
.A1(n_4587),
.A2(n_4479),
.B1(n_4569),
.B2(n_4563),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4643),
.B(n_4542),
.Y(n_4710)
);

AND2x2_ASAP7_75t_L g4711 ( 
.A(n_4631),
.B(n_4543),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4629),
.Y(n_4712)
);

NAND2xp5_ASAP7_75t_L g4713 ( 
.A(n_4636),
.B(n_4554),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4607),
.Y(n_4714)
);

AND2x2_ASAP7_75t_L g4715 ( 
.A(n_4670),
.B(n_4530),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4615),
.Y(n_4716)
);

AND2x2_ASAP7_75t_L g4717 ( 
.A(n_4625),
.B(n_4633),
.Y(n_4717)
);

AND2x2_ASAP7_75t_L g4718 ( 
.A(n_4609),
.B(n_4560),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4672),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4641),
.Y(n_4720)
);

INVx3_ASAP7_75t_L g4721 ( 
.A(n_4668),
.Y(n_4721)
);

INVx2_ASAP7_75t_SL g4722 ( 
.A(n_4619),
.Y(n_4722)
);

AND2x2_ASAP7_75t_SL g4723 ( 
.A(n_4622),
.B(n_4573),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4654),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4665),
.B(n_4464),
.Y(n_4725)
);

NOR2xp33_ASAP7_75t_SL g4726 ( 
.A(n_4617),
.B(n_4529),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_SL g4727 ( 
.A(n_4653),
.B(n_4533),
.Y(n_4727)
);

INVx2_ASAP7_75t_SL g4728 ( 
.A(n_4638),
.Y(n_4728)
);

OR2x2_ASAP7_75t_L g4729 ( 
.A(n_4628),
.B(n_4462),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4663),
.Y(n_4730)
);

OR2x2_ASAP7_75t_L g4731 ( 
.A(n_4632),
.B(n_243),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4610),
.Y(n_4732)
);

AND2x2_ASAP7_75t_L g4733 ( 
.A(n_4650),
.B(n_244),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_4695),
.Y(n_4734)
);

INVx1_ASAP7_75t_L g4735 ( 
.A(n_4733),
.Y(n_4735)
);

NAND2xp5_ASAP7_75t_L g4736 ( 
.A(n_4717),
.B(n_4637),
.Y(n_4736)
);

OR2x2_ASAP7_75t_L g4737 ( 
.A(n_4691),
.B(n_4614),
.Y(n_4737)
);

HB1xp67_ASAP7_75t_L g4738 ( 
.A(n_4677),
.Y(n_4738)
);

OR2x2_ASAP7_75t_L g4739 ( 
.A(n_4686),
.B(n_4594),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4706),
.B(n_4704),
.Y(n_4740)
);

INVx2_ASAP7_75t_L g4741 ( 
.A(n_4723),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4693),
.Y(n_4742)
);

INVx2_ASAP7_75t_L g4743 ( 
.A(n_4685),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4728),
.B(n_4647),
.Y(n_4744)
);

AND2x2_ASAP7_75t_SL g4745 ( 
.A(n_4697),
.B(n_4635),
.Y(n_4745)
);

AND2x2_ASAP7_75t_L g4746 ( 
.A(n_4688),
.B(n_4618),
.Y(n_4746)
);

AND2x4_ASAP7_75t_L g4747 ( 
.A(n_4722),
.B(n_4642),
.Y(n_4747)
);

INVx2_ASAP7_75t_SL g4748 ( 
.A(n_4715),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4718),
.B(n_4656),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4690),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4705),
.B(n_4623),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_L g4752 ( 
.A(n_4683),
.B(n_4639),
.Y(n_4752)
);

OAI22xp5_ASAP7_75t_L g4753 ( 
.A1(n_4675),
.A2(n_4620),
.B1(n_4627),
.B2(n_4605),
.Y(n_4753)
);

OAI32xp33_ASAP7_75t_L g4754 ( 
.A1(n_4680),
.A2(n_4648),
.A3(n_4593),
.B1(n_4592),
.B2(n_4658),
.Y(n_4754)
);

AND2x2_ASAP7_75t_L g4755 ( 
.A(n_4701),
.B(n_4666),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4689),
.Y(n_4756)
);

HB1xp67_ASAP7_75t_L g4757 ( 
.A(n_4721),
.Y(n_4757)
);

AND2x2_ASAP7_75t_L g4758 ( 
.A(n_4698),
.B(n_4667),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4707),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4700),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4682),
.B(n_4661),
.Y(n_4761)
);

OR2x6_ASAP7_75t_L g4762 ( 
.A(n_4687),
.B(n_4649),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4730),
.B(n_4630),
.Y(n_4763)
);

NAND2xp5_ASAP7_75t_L g4764 ( 
.A(n_4711),
.B(n_4644),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4684),
.B(n_4657),
.Y(n_4765)
);

AND2x2_ASAP7_75t_L g4766 ( 
.A(n_4702),
.B(n_4669),
.Y(n_4766)
);

AND2x2_ASAP7_75t_L g4767 ( 
.A(n_4681),
.B(n_4671),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4731),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4699),
.Y(n_4769)
);

AOI21xp5_ASAP7_75t_L g4770 ( 
.A1(n_4727),
.A2(n_4659),
.B(n_4662),
.Y(n_4770)
);

AND2x4_ASAP7_75t_L g4771 ( 
.A(n_4676),
.B(n_4645),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_SL g4772 ( 
.A(n_4726),
.B(n_244),
.Y(n_4772)
);

NAND4xp25_ASAP7_75t_L g4773 ( 
.A(n_4673),
.B(n_4732),
.C(n_4694),
.D(n_4674),
.Y(n_4773)
);

NAND2xp5_ASAP7_75t_SL g4774 ( 
.A(n_4696),
.B(n_4710),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_L g4775 ( 
.A(n_4719),
.B(n_245),
.Y(n_4775)
);

INVx3_ASAP7_75t_R g4776 ( 
.A(n_4729),
.Y(n_4776)
);

AND2x2_ASAP7_75t_L g4777 ( 
.A(n_4712),
.B(n_246),
.Y(n_4777)
);

NAND2x1p5_ASAP7_75t_L g4778 ( 
.A(n_4692),
.B(n_246),
.Y(n_4778)
);

AOI22xp5_ASAP7_75t_L g4779 ( 
.A1(n_4709),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.Y(n_4779)
);

NAND3xp33_ASAP7_75t_L g4780 ( 
.A(n_4679),
.B(n_247),
.C(n_248),
.Y(n_4780)
);

AOI21xp5_ASAP7_75t_L g4781 ( 
.A1(n_4770),
.A2(n_4708),
.B(n_4725),
.Y(n_4781)
);

NOR3xp33_ASAP7_75t_L g4782 ( 
.A(n_4764),
.B(n_4713),
.C(n_4714),
.Y(n_4782)
);

CKINVDCx16_ASAP7_75t_R g4783 ( 
.A(n_4767),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4738),
.Y(n_4784)
);

AOI22xp5_ASAP7_75t_L g4785 ( 
.A1(n_4762),
.A2(n_4720),
.B1(n_4724),
.B2(n_4716),
.Y(n_4785)
);

XNOR2xp5_ASAP7_75t_L g4786 ( 
.A(n_4745),
.B(n_4678),
.Y(n_4786)
);

AOI21xp33_ASAP7_75t_L g4787 ( 
.A1(n_4749),
.A2(n_4703),
.B(n_249),
.Y(n_4787)
);

NOR2xp33_ASAP7_75t_L g4788 ( 
.A(n_4736),
.B(n_250),
.Y(n_4788)
);

OAI21xp5_ASAP7_75t_L g4789 ( 
.A1(n_4740),
.A2(n_251),
.B(n_253),
.Y(n_4789)
);

OAI21xp5_ASAP7_75t_L g4790 ( 
.A1(n_4748),
.A2(n_251),
.B(n_253),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_L g4791 ( 
.A(n_4735),
.B(n_254),
.Y(n_4791)
);

OAI21xp5_ASAP7_75t_L g4792 ( 
.A1(n_4765),
.A2(n_254),
.B(n_255),
.Y(n_4792)
);

AOI22xp33_ASAP7_75t_L g4793 ( 
.A1(n_4768),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_4793)
);

AND2x4_ASAP7_75t_L g4794 ( 
.A(n_4747),
.B(n_256),
.Y(n_4794)
);

OAI21xp5_ASAP7_75t_L g4795 ( 
.A1(n_4761),
.A2(n_258),
.B(n_259),
.Y(n_4795)
);

AOI22xp5_ASAP7_75t_L g4796 ( 
.A1(n_4762),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_4796)
);

AOI211xp5_ASAP7_75t_L g4797 ( 
.A1(n_4754),
.A2(n_263),
.B(n_260),
.C(n_262),
.Y(n_4797)
);

NAND2xp5_ASAP7_75t_L g4798 ( 
.A(n_4758),
.B(n_4766),
.Y(n_4798)
);

OAI211xp5_ASAP7_75t_SL g4799 ( 
.A1(n_4752),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_4799)
);

OAI21xp5_ASAP7_75t_L g4800 ( 
.A1(n_4757),
.A2(n_264),
.B(n_265),
.Y(n_4800)
);

AOI21xp5_ASAP7_75t_L g4801 ( 
.A1(n_4772),
.A2(n_265),
.B(n_266),
.Y(n_4801)
);

INVx2_ASAP7_75t_L g4802 ( 
.A(n_4778),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_4751),
.Y(n_4803)
);

OA22x2_ASAP7_75t_L g4804 ( 
.A1(n_4741),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_4804)
);

HB1xp67_ASAP7_75t_L g4805 ( 
.A(n_4743),
.Y(n_4805)
);

NOR3xp33_ASAP7_75t_L g4806 ( 
.A(n_4774),
.B(n_269),
.C(n_271),
.Y(n_4806)
);

OAI221xp5_ASAP7_75t_SL g4807 ( 
.A1(n_4739),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.C(n_274),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4777),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4759),
.Y(n_4809)
);

HB1xp67_ASAP7_75t_L g4810 ( 
.A(n_4760),
.Y(n_4810)
);

AOI21xp5_ASAP7_75t_L g4811 ( 
.A1(n_4773),
.A2(n_272),
.B(n_274),
.Y(n_4811)
);

BUFx12f_ASAP7_75t_L g4812 ( 
.A(n_4746),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4755),
.Y(n_4813)
);

OAI22xp5_ASAP7_75t_L g4814 ( 
.A1(n_4756),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4734),
.Y(n_4815)
);

AOI211xp5_ASAP7_75t_L g4816 ( 
.A1(n_4753),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_4816)
);

OAI21xp5_ASAP7_75t_L g4817 ( 
.A1(n_4742),
.A2(n_278),
.B(n_279),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4771),
.Y(n_4818)
);

AOI22xp5_ASAP7_75t_L g4819 ( 
.A1(n_4750),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_4819)
);

NOR3xp33_ASAP7_75t_L g4820 ( 
.A(n_4775),
.B(n_280),
.C(n_283),
.Y(n_4820)
);

INVx2_ASAP7_75t_L g4821 ( 
.A(n_4737),
.Y(n_4821)
);

INVx1_ASAP7_75t_SL g4822 ( 
.A(n_4763),
.Y(n_4822)
);

XNOR2xp5_ASAP7_75t_L g4823 ( 
.A(n_4779),
.B(n_283),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_4744),
.Y(n_4824)
);

OAI21xp33_ASAP7_75t_SL g4825 ( 
.A1(n_4769),
.A2(n_284),
.B(n_285),
.Y(n_4825)
);

INVx1_ASAP7_75t_SL g4826 ( 
.A(n_4780),
.Y(n_4826)
);

AOI22xp33_ASAP7_75t_SL g4827 ( 
.A1(n_4776),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_4827)
);

INVx1_ASAP7_75t_L g4828 ( 
.A(n_4764),
.Y(n_4828)
);

NOR2xp33_ASAP7_75t_L g4829 ( 
.A(n_4783),
.B(n_286),
.Y(n_4829)
);

OAI22xp5_ASAP7_75t_L g4830 ( 
.A1(n_4786),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_4830)
);

AOI32xp33_ASAP7_75t_L g4831 ( 
.A1(n_4782),
.A2(n_289),
.A3(n_287),
.B1(n_288),
.B2(n_290),
.Y(n_4831)
);

NOR3xp33_ASAP7_75t_L g4832 ( 
.A(n_4787),
.B(n_291),
.C(n_292),
.Y(n_4832)
);

AND2x2_ASAP7_75t_L g4833 ( 
.A(n_4805),
.B(n_292),
.Y(n_4833)
);

AOI21xp5_ASAP7_75t_L g4834 ( 
.A1(n_4781),
.A2(n_295),
.B(n_294),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_SL g4835 ( 
.A(n_4812),
.B(n_4798),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_4804),
.Y(n_4836)
);

OAI21xp5_ASAP7_75t_SL g4837 ( 
.A1(n_4822),
.A2(n_293),
.B(n_294),
.Y(n_4837)
);

INVxp67_ASAP7_75t_L g4838 ( 
.A(n_4810),
.Y(n_4838)
);

OAI22xp33_ASAP7_75t_SL g4839 ( 
.A1(n_4808),
.A2(n_296),
.B1(n_293),
.B2(n_295),
.Y(n_4839)
);

AOI21xp33_ASAP7_75t_L g4840 ( 
.A1(n_4825),
.A2(n_296),
.B(n_297),
.Y(n_4840)
);

OAI21xp33_ASAP7_75t_L g4841 ( 
.A1(n_4818),
.A2(n_297),
.B(n_298),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4813),
.Y(n_4842)
);

OAI21xp5_ASAP7_75t_L g4843 ( 
.A1(n_4811),
.A2(n_298),
.B(n_300),
.Y(n_4843)
);

NOR2x1_ASAP7_75t_L g4844 ( 
.A(n_4794),
.B(n_301),
.Y(n_4844)
);

OR2x2_ASAP7_75t_L g4845 ( 
.A(n_4784),
.B(n_302),
.Y(n_4845)
);

OAI22xp33_ASAP7_75t_L g4846 ( 
.A1(n_4826),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.Y(n_4846)
);

AND2x4_ASAP7_75t_L g4847 ( 
.A(n_4794),
.B(n_305),
.Y(n_4847)
);

OAI221xp5_ASAP7_75t_L g4848 ( 
.A1(n_4785),
.A2(n_4802),
.B1(n_4797),
.B2(n_4827),
.C(n_4792),
.Y(n_4848)
);

NAND2xp5_ASAP7_75t_L g4849 ( 
.A(n_4788),
.B(n_308),
.Y(n_4849)
);

AOI22xp5_ASAP7_75t_L g4850 ( 
.A1(n_4820),
.A2(n_4821),
.B1(n_4799),
.B2(n_4806),
.Y(n_4850)
);

O2A1O1Ixp33_ASAP7_75t_L g4851 ( 
.A1(n_4816),
.A2(n_310),
.B(n_308),
.C(n_309),
.Y(n_4851)
);

OAI22xp5_ASAP7_75t_L g4852 ( 
.A1(n_4828),
.A2(n_312),
.B1(n_309),
.B2(n_311),
.Y(n_4852)
);

INVxp33_ASAP7_75t_L g4853 ( 
.A(n_4823),
.Y(n_4853)
);

AND2x2_ASAP7_75t_L g4854 ( 
.A(n_4803),
.B(n_312),
.Y(n_4854)
);

INVx2_ASAP7_75t_L g4855 ( 
.A(n_4824),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4801),
.B(n_313),
.Y(n_4856)
);

AOI221xp5_ASAP7_75t_L g4857 ( 
.A1(n_4795),
.A2(n_333),
.B1(n_343),
.B2(n_323),
.C(n_313),
.Y(n_4857)
);

OAI221xp5_ASAP7_75t_L g4858 ( 
.A1(n_4791),
.A2(n_318),
.B1(n_314),
.B2(n_317),
.C(n_319),
.Y(n_4858)
);

AND2x4_ASAP7_75t_L g4859 ( 
.A(n_4815),
.B(n_317),
.Y(n_4859)
);

NAND2x1_ASAP7_75t_L g4860 ( 
.A(n_4809),
.B(n_318),
.Y(n_4860)
);

NOR2xp33_ASAP7_75t_L g4861 ( 
.A(n_4807),
.B(n_319),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4796),
.B(n_320),
.Y(n_4862)
);

INVx2_ASAP7_75t_L g4863 ( 
.A(n_4819),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4814),
.Y(n_4864)
);

INVx1_ASAP7_75t_SL g4865 ( 
.A(n_4789),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_L g4866 ( 
.A(n_4793),
.B(n_320),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4817),
.Y(n_4867)
);

XNOR2xp5_ASAP7_75t_L g4868 ( 
.A(n_4790),
.B(n_321),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4800),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4805),
.Y(n_4870)
);

INVx1_ASAP7_75t_L g4871 ( 
.A(n_4805),
.Y(n_4871)
);

HB1xp67_ASAP7_75t_L g4872 ( 
.A(n_4783),
.Y(n_4872)
);

AOI211xp5_ASAP7_75t_L g4873 ( 
.A1(n_4786),
.A2(n_325),
.B(n_322),
.C(n_323),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4805),
.Y(n_4874)
);

INVxp67_ASAP7_75t_L g4875 ( 
.A(n_4805),
.Y(n_4875)
);

OAI21xp5_ASAP7_75t_L g4876 ( 
.A1(n_4786),
.A2(n_326),
.B(n_327),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4805),
.Y(n_4877)
);

INVx2_ASAP7_75t_L g4878 ( 
.A(n_4783),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4783),
.B(n_326),
.Y(n_4879)
);

NAND2x1p5_ASAP7_75t_L g4880 ( 
.A(n_4794),
.B(n_327),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4783),
.B(n_329),
.Y(n_4881)
);

INVx1_ASAP7_75t_L g4882 ( 
.A(n_4805),
.Y(n_4882)
);

INVx1_ASAP7_75t_SL g4883 ( 
.A(n_4783),
.Y(n_4883)
);

AND2x2_ASAP7_75t_L g4884 ( 
.A(n_4783),
.B(n_329),
.Y(n_4884)
);

NAND3xp33_ASAP7_75t_L g4885 ( 
.A(n_4797),
.B(n_330),
.C(n_331),
.Y(n_4885)
);

AOI21xp5_ASAP7_75t_L g4886 ( 
.A1(n_4786),
.A2(n_332),
.B(n_331),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4805),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4805),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4872),
.Y(n_4889)
);

HB1xp67_ASAP7_75t_L g4890 ( 
.A(n_4883),
.Y(n_4890)
);

AOI22xp5_ASAP7_75t_L g4891 ( 
.A1(n_4878),
.A2(n_333),
.B1(n_330),
.B2(n_332),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4884),
.Y(n_4892)
);

AOI21xp5_ASAP7_75t_L g4893 ( 
.A1(n_4835),
.A2(n_334),
.B(n_335),
.Y(n_4893)
);

OR2x2_ASAP7_75t_L g4894 ( 
.A(n_4879),
.B(n_334),
.Y(n_4894)
);

AOI22xp33_ASAP7_75t_L g4895 ( 
.A1(n_4840),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_4895)
);

HB1xp67_ASAP7_75t_L g4896 ( 
.A(n_4880),
.Y(n_4896)
);

AND2x2_ASAP7_75t_L g4897 ( 
.A(n_4875),
.B(n_338),
.Y(n_4897)
);

A2O1A1Ixp33_ASAP7_75t_L g4898 ( 
.A1(n_4834),
.A2(n_343),
.B(n_341),
.C(n_342),
.Y(n_4898)
);

AOI21xp33_ASAP7_75t_L g4899 ( 
.A1(n_4853),
.A2(n_4836),
.B(n_4865),
.Y(n_4899)
);

NAND2xp5_ASAP7_75t_L g4900 ( 
.A(n_4847),
.B(n_344),
.Y(n_4900)
);

NOR3xp33_ASAP7_75t_SL g4901 ( 
.A(n_4848),
.B(n_344),
.C(n_345),
.Y(n_4901)
);

INVx1_ASAP7_75t_SL g4902 ( 
.A(n_4833),
.Y(n_4902)
);

O2A1O1Ixp33_ASAP7_75t_SL g4903 ( 
.A1(n_4838),
.A2(n_348),
.B(n_345),
.C(n_346),
.Y(n_4903)
);

BUFx2_ASAP7_75t_SL g4904 ( 
.A(n_4870),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4881),
.Y(n_4905)
);

AND2x2_ASAP7_75t_L g4906 ( 
.A(n_4871),
.B(n_346),
.Y(n_4906)
);

INVx1_ASAP7_75t_L g4907 ( 
.A(n_4844),
.Y(n_4907)
);

OAI21xp5_ASAP7_75t_SL g4908 ( 
.A1(n_4874),
.A2(n_349),
.B(n_350),
.Y(n_4908)
);

AOI22xp33_ASAP7_75t_L g4909 ( 
.A1(n_4863),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.Y(n_4909)
);

AOI221xp5_ASAP7_75t_L g4910 ( 
.A1(n_4876),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.C(n_357),
.Y(n_4910)
);

AOI21xp5_ASAP7_75t_L g4911 ( 
.A1(n_4860),
.A2(n_354),
.B(n_355),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4829),
.Y(n_4912)
);

OAI222xp33_ASAP7_75t_L g4913 ( 
.A1(n_4850),
.A2(n_4888),
.B1(n_4882),
.B2(n_4887),
.C1(n_4877),
.C2(n_4864),
.Y(n_4913)
);

NOR2xp33_ASAP7_75t_L g4914 ( 
.A(n_4837),
.B(n_357),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4854),
.Y(n_4915)
);

XNOR2x1_ASAP7_75t_L g4916 ( 
.A(n_4868),
.B(n_358),
.Y(n_4916)
);

AND2x2_ASAP7_75t_L g4917 ( 
.A(n_4842),
.B(n_358),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_L g4918 ( 
.A(n_4847),
.B(n_360),
.Y(n_4918)
);

OAI21xp5_ASAP7_75t_L g4919 ( 
.A1(n_4886),
.A2(n_360),
.B(n_361),
.Y(n_4919)
);

INVxp67_ASAP7_75t_L g4920 ( 
.A(n_4849),
.Y(n_4920)
);

OAI21xp33_ASAP7_75t_L g4921 ( 
.A1(n_4869),
.A2(n_4867),
.B(n_4855),
.Y(n_4921)
);

AOI21xp5_ASAP7_75t_L g4922 ( 
.A1(n_4856),
.A2(n_361),
.B(n_362),
.Y(n_4922)
);

NOR2xp33_ASAP7_75t_SL g4923 ( 
.A(n_4841),
.B(n_362),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4859),
.Y(n_4924)
);

OAI21xp5_ASAP7_75t_L g4925 ( 
.A1(n_4885),
.A2(n_363),
.B(n_364),
.Y(n_4925)
);

OAI22xp33_ASAP7_75t_L g4926 ( 
.A1(n_4845),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_4926)
);

INVxp67_ASAP7_75t_SL g4927 ( 
.A(n_4873),
.Y(n_4927)
);

INVx1_ASAP7_75t_L g4928 ( 
.A(n_4859),
.Y(n_4928)
);

NAND2xp33_ASAP7_75t_R g4929 ( 
.A(n_4861),
.B(n_367),
.Y(n_4929)
);

AND2x2_ASAP7_75t_L g4930 ( 
.A(n_4843),
.B(n_367),
.Y(n_4930)
);

NAND2xp5_ASAP7_75t_L g4931 ( 
.A(n_4831),
.B(n_369),
.Y(n_4931)
);

INVx2_ASAP7_75t_L g4932 ( 
.A(n_4862),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4839),
.Y(n_4933)
);

AND2x2_ASAP7_75t_L g4934 ( 
.A(n_4830),
.B(n_4832),
.Y(n_4934)
);

NOR2x1_ASAP7_75t_L g4935 ( 
.A(n_4846),
.B(n_370),
.Y(n_4935)
);

AOI21xp5_ASAP7_75t_L g4936 ( 
.A1(n_4851),
.A2(n_370),
.B(n_372),
.Y(n_4936)
);

OAI22xp33_ASAP7_75t_L g4937 ( 
.A1(n_4866),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_4937)
);

INVx2_ASAP7_75t_SL g4938 ( 
.A(n_4852),
.Y(n_4938)
);

A2O1A1Ixp33_ASAP7_75t_L g4939 ( 
.A1(n_4857),
.A2(n_377),
.B(n_375),
.C(n_376),
.Y(n_4939)
);

AND2x2_ASAP7_75t_L g4940 ( 
.A(n_4858),
.B(n_375),
.Y(n_4940)
);

AOI22xp5_ASAP7_75t_L g4941 ( 
.A1(n_4883),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_4941)
);

NAND2xp5_ASAP7_75t_SL g4942 ( 
.A(n_4883),
.B(n_378),
.Y(n_4942)
);

NAND2xp5_ASAP7_75t_L g4943 ( 
.A(n_4883),
.B(n_379),
.Y(n_4943)
);

NAND2xp33_ASAP7_75t_SL g4944 ( 
.A(n_4872),
.B(n_380),
.Y(n_4944)
);

AND2x4_ASAP7_75t_L g4945 ( 
.A(n_4878),
.B(n_380),
.Y(n_4945)
);

NOR2xp33_ASAP7_75t_L g4946 ( 
.A(n_4883),
.B(n_381),
.Y(n_4946)
);

OAI211xp5_ASAP7_75t_SL g4947 ( 
.A1(n_4883),
.A2(n_383),
.B(n_381),
.C(n_382),
.Y(n_4947)
);

AOI21xp33_ASAP7_75t_L g4948 ( 
.A1(n_4853),
.A2(n_382),
.B(n_384),
.Y(n_4948)
);

AND2x2_ASAP7_75t_L g4949 ( 
.A(n_4872),
.B(n_385),
.Y(n_4949)
);

AOI22xp33_ASAP7_75t_L g4950 ( 
.A1(n_4840),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_4950)
);

OAI221xp5_ASAP7_75t_L g4951 ( 
.A1(n_4883),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.C(n_390),
.Y(n_4951)
);

NOR2xp33_ASAP7_75t_L g4952 ( 
.A(n_4883),
.B(n_388),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_L g4953 ( 
.A(n_4883),
.B(n_391),
.Y(n_4953)
);

INVxp67_ASAP7_75t_SL g4954 ( 
.A(n_4872),
.Y(n_4954)
);

AOI221xp5_ASAP7_75t_SL g4955 ( 
.A1(n_4875),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.C(n_395),
.Y(n_4955)
);

NAND3xp33_ASAP7_75t_L g4956 ( 
.A(n_4872),
.B(n_401),
.C(n_392),
.Y(n_4956)
);

AOI31xp33_ASAP7_75t_L g4957 ( 
.A1(n_4872),
.A2(n_396),
.A3(n_393),
.B(n_394),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4872),
.Y(n_4958)
);

HB1xp67_ASAP7_75t_L g4959 ( 
.A(n_4872),
.Y(n_4959)
);

INVx2_ASAP7_75t_L g4960 ( 
.A(n_4880),
.Y(n_4960)
);

OAI22xp5_ASAP7_75t_L g4961 ( 
.A1(n_4883),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4872),
.Y(n_4962)
);

AND2x2_ASAP7_75t_L g4963 ( 
.A(n_4872),
.B(n_397),
.Y(n_4963)
);

NOR2xp33_ASAP7_75t_R g4964 ( 
.A(n_4883),
.B(n_399),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4872),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4872),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4872),
.Y(n_4967)
);

OAI21xp5_ASAP7_75t_L g4968 ( 
.A1(n_4872),
.A2(n_398),
.B(n_400),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4872),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4872),
.Y(n_4970)
);

OR2x2_ASAP7_75t_L g4971 ( 
.A(n_4883),
.B(n_400),
.Y(n_4971)
);

NOR2x1_ASAP7_75t_L g4972 ( 
.A(n_4878),
.B(n_402),
.Y(n_4972)
);

AOI31xp33_ASAP7_75t_L g4973 ( 
.A1(n_4872),
.A2(n_404),
.A3(n_402),
.B(n_403),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4872),
.Y(n_4974)
);

AOI211xp5_ASAP7_75t_L g4975 ( 
.A1(n_4883),
.A2(n_405),
.B(n_403),
.C(n_404),
.Y(n_4975)
);

OAI21xp33_ASAP7_75t_L g4976 ( 
.A1(n_4883),
.A2(n_406),
.B(n_407),
.Y(n_4976)
);

XNOR2xp5_ASAP7_75t_L g4977 ( 
.A(n_4872),
.B(n_406),
.Y(n_4977)
);

OAI32xp33_ASAP7_75t_L g4978 ( 
.A1(n_4883),
.A2(n_409),
.A3(n_407),
.B1(n_408),
.B2(n_410),
.Y(n_4978)
);

XNOR2xp5_ASAP7_75t_L g4979 ( 
.A(n_4872),
.B(n_408),
.Y(n_4979)
);

AOI21xp5_ASAP7_75t_L g4980 ( 
.A1(n_4883),
.A2(n_409),
.B(n_410),
.Y(n_4980)
);

INVx1_ASAP7_75t_SL g4981 ( 
.A(n_4964),
.Y(n_4981)
);

AOI221xp5_ASAP7_75t_L g4982 ( 
.A1(n_4944),
.A2(n_413),
.B1(n_411),
.B2(n_412),
.C(n_414),
.Y(n_4982)
);

AOI211xp5_ASAP7_75t_L g4983 ( 
.A1(n_4954),
.A2(n_415),
.B(n_411),
.C(n_414),
.Y(n_4983)
);

NOR2xp33_ASAP7_75t_SL g4984 ( 
.A(n_4890),
.B(n_415),
.Y(n_4984)
);

NOR2xp33_ASAP7_75t_L g4985 ( 
.A(n_4947),
.B(n_4957),
.Y(n_4985)
);

NOR2xp33_ASAP7_75t_L g4986 ( 
.A(n_4973),
.B(n_416),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4959),
.Y(n_4987)
);

AOI211xp5_ASAP7_75t_L g4988 ( 
.A1(n_4913),
.A2(n_4921),
.B(n_4899),
.C(n_4889),
.Y(n_4988)
);

NOR2xp33_ASAP7_75t_L g4989 ( 
.A(n_4907),
.B(n_416),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4945),
.B(n_417),
.Y(n_4990)
);

INVx1_ASAP7_75t_L g4991 ( 
.A(n_4977),
.Y(n_4991)
);

O2A1O1Ixp33_ASAP7_75t_L g4992 ( 
.A1(n_4896),
.A2(n_419),
.B(n_417),
.C(n_418),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_SL g4993 ( 
.A(n_4945),
.B(n_418),
.Y(n_4993)
);

NAND2xp33_ASAP7_75t_L g4994 ( 
.A(n_4958),
.B(n_419),
.Y(n_4994)
);

AOI22xp5_ASAP7_75t_L g4995 ( 
.A1(n_4892),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_4995)
);

NAND2xp5_ASAP7_75t_L g4996 ( 
.A(n_4902),
.B(n_420),
.Y(n_4996)
);

NAND3xp33_ASAP7_75t_SL g4997 ( 
.A(n_4962),
.B(n_422),
.C(n_424),
.Y(n_4997)
);

AOI221xp5_ASAP7_75t_L g4998 ( 
.A1(n_4905),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.C(n_428),
.Y(n_4998)
);

INVx2_ASAP7_75t_L g4999 ( 
.A(n_4916),
.Y(n_4999)
);

NOR2xp33_ASAP7_75t_SL g5000 ( 
.A(n_4949),
.B(n_426),
.Y(n_5000)
);

NOR3x1_ASAP7_75t_L g5001 ( 
.A(n_4908),
.B(n_428),
.C(n_430),
.Y(n_5001)
);

NAND3xp33_ASAP7_75t_L g5002 ( 
.A(n_4901),
.B(n_430),
.C(n_431),
.Y(n_5002)
);

NAND3xp33_ASAP7_75t_L g5003 ( 
.A(n_4972),
.B(n_431),
.C(n_432),
.Y(n_5003)
);

NAND2xp5_ASAP7_75t_SL g5004 ( 
.A(n_4955),
.B(n_433),
.Y(n_5004)
);

NAND4xp25_ASAP7_75t_L g5005 ( 
.A(n_4965),
.B(n_435),
.C(n_436),
.D(n_434),
.Y(n_5005)
);

NOR2xp33_ASAP7_75t_L g5006 ( 
.A(n_4924),
.B(n_433),
.Y(n_5006)
);

NAND3xp33_ASAP7_75t_L g5007 ( 
.A(n_4975),
.B(n_434),
.C(n_435),
.Y(n_5007)
);

NOR3x1_ASAP7_75t_L g5008 ( 
.A(n_4968),
.B(n_436),
.C(n_437),
.Y(n_5008)
);

INVx1_ASAP7_75t_L g5009 ( 
.A(n_4979),
.Y(n_5009)
);

NAND2xp5_ASAP7_75t_L g5010 ( 
.A(n_4911),
.B(n_438),
.Y(n_5010)
);

NAND3xp33_ASAP7_75t_SL g5011 ( 
.A(n_4966),
.B(n_438),
.C(n_439),
.Y(n_5011)
);

OR2x2_ASAP7_75t_L g5012 ( 
.A(n_4904),
.B(n_439),
.Y(n_5012)
);

AND2x2_ASAP7_75t_L g5013 ( 
.A(n_4963),
.B(n_441),
.Y(n_5013)
);

OR2x2_ASAP7_75t_L g5014 ( 
.A(n_4971),
.B(n_441),
.Y(n_5014)
);

NOR4xp75_ASAP7_75t_L g5015 ( 
.A(n_4942),
.B(n_444),
.C(n_442),
.D(n_443),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_L g5016 ( 
.A(n_4928),
.B(n_442),
.Y(n_5016)
);

NOR2xp33_ASAP7_75t_L g5017 ( 
.A(n_4903),
.B(n_443),
.Y(n_5017)
);

NAND3xp33_ASAP7_75t_L g5018 ( 
.A(n_4946),
.B(n_4952),
.C(n_4967),
.Y(n_5018)
);

AO22x2_ASAP7_75t_L g5019 ( 
.A1(n_4933),
.A2(n_447),
.B1(n_445),
.B2(n_446),
.Y(n_5019)
);

INVx1_ASAP7_75t_L g5020 ( 
.A(n_4900),
.Y(n_5020)
);

AOI221xp5_ASAP7_75t_L g5021 ( 
.A1(n_4912),
.A2(n_448),
.B1(n_445),
.B2(n_446),
.C(n_449),
.Y(n_5021)
);

NAND2xp5_ASAP7_75t_L g5022 ( 
.A(n_4960),
.B(n_449),
.Y(n_5022)
);

OA22x2_ASAP7_75t_L g5023 ( 
.A1(n_4969),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.Y(n_5023)
);

OR2x2_ASAP7_75t_L g5024 ( 
.A(n_4943),
.B(n_451),
.Y(n_5024)
);

AOI221xp5_ASAP7_75t_L g5025 ( 
.A1(n_4922),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.C(n_455),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4918),
.Y(n_5026)
);

AOI21xp5_ASAP7_75t_L g5027 ( 
.A1(n_4980),
.A2(n_453),
.B(n_455),
.Y(n_5027)
);

NOR2xp33_ASAP7_75t_L g5028 ( 
.A(n_4978),
.B(n_456),
.Y(n_5028)
);

AOI211xp5_ASAP7_75t_L g5029 ( 
.A1(n_4970),
.A2(n_460),
.B(n_456),
.C(n_458),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4917),
.Y(n_5030)
);

INVx1_ASAP7_75t_SL g5031 ( 
.A(n_4906),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_4894),
.Y(n_5032)
);

NOR2xp33_ASAP7_75t_L g5033 ( 
.A(n_4915),
.B(n_458),
.Y(n_5033)
);

INVx1_ASAP7_75t_L g5034 ( 
.A(n_4897),
.Y(n_5034)
);

AOI21xp33_ASAP7_75t_L g5035 ( 
.A1(n_4929),
.A2(n_460),
.B(n_461),
.Y(n_5035)
);

INVxp67_ASAP7_75t_SL g5036 ( 
.A(n_4914),
.Y(n_5036)
);

NOR3xp33_ASAP7_75t_L g5037 ( 
.A(n_4974),
.B(n_462),
.C(n_463),
.Y(n_5037)
);

INVx2_ASAP7_75t_L g5038 ( 
.A(n_4930),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_L g5039 ( 
.A(n_4920),
.B(n_462),
.Y(n_5039)
);

NAND4xp25_ASAP7_75t_L g5040 ( 
.A(n_4934),
.B(n_466),
.C(n_469),
.D(n_465),
.Y(n_5040)
);

NAND2xp33_ASAP7_75t_L g5041 ( 
.A(n_4953),
.B(n_464),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_4927),
.B(n_464),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_4898),
.B(n_465),
.Y(n_5043)
);

INVx2_ASAP7_75t_SL g5044 ( 
.A(n_4935),
.Y(n_5044)
);

AOI211xp5_ASAP7_75t_L g5045 ( 
.A1(n_4893),
.A2(n_4956),
.B(n_4976),
.C(n_4919),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_4931),
.Y(n_5046)
);

NAND2xp5_ASAP7_75t_L g5047 ( 
.A(n_4895),
.B(n_466),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4941),
.Y(n_5048)
);

NAND3xp33_ASAP7_75t_L g5049 ( 
.A(n_4950),
.B(n_469),
.C(n_470),
.Y(n_5049)
);

NOR2xp33_ASAP7_75t_L g5050 ( 
.A(n_4923),
.B(n_470),
.Y(n_5050)
);

AND2x2_ASAP7_75t_L g5051 ( 
.A(n_4940),
.B(n_471),
.Y(n_5051)
);

NAND2xp5_ASAP7_75t_L g5052 ( 
.A(n_4926),
.B(n_471),
.Y(n_5052)
);

NOR3xp33_ASAP7_75t_SL g5053 ( 
.A(n_4951),
.B(n_473),
.C(n_474),
.Y(n_5053)
);

NAND2xp5_ASAP7_75t_L g5054 ( 
.A(n_4936),
.B(n_473),
.Y(n_5054)
);

AOI221xp5_ASAP7_75t_L g5055 ( 
.A1(n_4932),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.C(n_479),
.Y(n_5055)
);

OAI21xp33_ASAP7_75t_SL g5056 ( 
.A1(n_4938),
.A2(n_475),
.B(n_477),
.Y(n_5056)
);

NAND3xp33_ASAP7_75t_L g5057 ( 
.A(n_4910),
.B(n_479),
.C(n_480),
.Y(n_5057)
);

NOR2xp33_ASAP7_75t_L g5058 ( 
.A(n_4948),
.B(n_480),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_L g5059 ( 
.A(n_4909),
.B(n_481),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_4961),
.Y(n_5060)
);

OAI22xp5_ASAP7_75t_L g5061 ( 
.A1(n_4891),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_4937),
.B(n_483),
.Y(n_5062)
);

AOI221xp5_ASAP7_75t_L g5063 ( 
.A1(n_4925),
.A2(n_486),
.B1(n_484),
.B2(n_485),
.C(n_489),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_4939),
.Y(n_5064)
);

INVx2_ASAP7_75t_L g5065 ( 
.A(n_4916),
.Y(n_5065)
);

NAND2xp5_ASAP7_75t_SL g5066 ( 
.A(n_4945),
.B(n_484),
.Y(n_5066)
);

AOI21xp5_ASAP7_75t_L g5067 ( 
.A1(n_4954),
.A2(n_485),
.B(n_490),
.Y(n_5067)
);

NOR3xp33_ASAP7_75t_L g5068 ( 
.A(n_4899),
.B(n_490),
.C(n_491),
.Y(n_5068)
);

OAI211xp5_ASAP7_75t_L g5069 ( 
.A1(n_4988),
.A2(n_493),
.B(n_491),
.C(n_492),
.Y(n_5069)
);

AOI22xp5_ASAP7_75t_L g5070 ( 
.A1(n_4981),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.Y(n_5070)
);

AOI22xp5_ASAP7_75t_L g5071 ( 
.A1(n_4985),
.A2(n_497),
.B1(n_494),
.B2(n_495),
.Y(n_5071)
);

OAI221xp5_ASAP7_75t_L g5072 ( 
.A1(n_4984),
.A2(n_498),
.B1(n_495),
.B2(n_497),
.C(n_499),
.Y(n_5072)
);

NAND2xp5_ASAP7_75t_L g5073 ( 
.A(n_5013),
.B(n_498),
.Y(n_5073)
);

AOI21xp5_ASAP7_75t_L g5074 ( 
.A1(n_4994),
.A2(n_5004),
.B(n_4987),
.Y(n_5074)
);

AOI221xp5_ASAP7_75t_L g5075 ( 
.A1(n_5035),
.A2(n_5046),
.B1(n_5027),
.B2(n_5018),
.C(n_5031),
.Y(n_5075)
);

NOR4xp25_ASAP7_75t_L g5076 ( 
.A(n_5044),
.B(n_501),
.C(n_499),
.D(n_500),
.Y(n_5076)
);

OAI21xp5_ASAP7_75t_SL g5077 ( 
.A1(n_5068),
.A2(n_502),
.B(n_503),
.Y(n_5077)
);

OAI211xp5_ASAP7_75t_L g5078 ( 
.A1(n_5056),
.A2(n_504),
.B(n_502),
.C(n_503),
.Y(n_5078)
);

OAI22xp33_ASAP7_75t_L g5079 ( 
.A1(n_5012),
.A2(n_506),
.B1(n_504),
.B2(n_505),
.Y(n_5079)
);

AOI221xp5_ASAP7_75t_L g5080 ( 
.A1(n_5020),
.A2(n_5026),
.B1(n_5045),
.B2(n_5048),
.C(n_5030),
.Y(n_5080)
);

OAI22xp5_ASAP7_75t_L g5081 ( 
.A1(n_5060),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_5081)
);

NAND4xp25_ASAP7_75t_L g5082 ( 
.A(n_5001),
.B(n_5008),
.C(n_5002),
.D(n_5007),
.Y(n_5082)
);

AOI22xp33_ASAP7_75t_L g5083 ( 
.A1(n_5032),
.A2(n_510),
.B1(n_508),
.B2(n_509),
.Y(n_5083)
);

OAI221xp5_ASAP7_75t_L g5084 ( 
.A1(n_5017),
.A2(n_510),
.B1(n_508),
.B2(n_509),
.C(n_511),
.Y(n_5084)
);

NOR3xp33_ASAP7_75t_L g5085 ( 
.A(n_4999),
.B(n_512),
.C(n_514),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_5019),
.Y(n_5086)
);

NAND3xp33_ASAP7_75t_L g5087 ( 
.A(n_5000),
.B(n_515),
.C(n_514),
.Y(n_5087)
);

AOI21xp5_ASAP7_75t_L g5088 ( 
.A1(n_5067),
.A2(n_512),
.B(n_515),
.Y(n_5088)
);

NAND3xp33_ASAP7_75t_L g5089 ( 
.A(n_4986),
.B(n_518),
.C(n_517),
.Y(n_5089)
);

AOI21xp5_ASAP7_75t_L g5090 ( 
.A1(n_4992),
.A2(n_516),
.B(n_517),
.Y(n_5090)
);

AOI211xp5_ASAP7_75t_L g5091 ( 
.A1(n_4997),
.A2(n_520),
.B(n_518),
.C(n_519),
.Y(n_5091)
);

AOI21xp5_ASAP7_75t_L g5092 ( 
.A1(n_5011),
.A2(n_520),
.B(n_521),
.Y(n_5092)
);

NOR3xp33_ASAP7_75t_L g5093 ( 
.A(n_5065),
.B(n_521),
.C(n_522),
.Y(n_5093)
);

HB1xp67_ASAP7_75t_L g5094 ( 
.A(n_5015),
.Y(n_5094)
);

OAI221xp5_ASAP7_75t_SL g5095 ( 
.A1(n_4991),
.A2(n_524),
.B1(n_522),
.B2(n_523),
.C(n_525),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_5019),
.Y(n_5096)
);

O2A1O1Ixp33_ASAP7_75t_L g5097 ( 
.A1(n_4996),
.A2(n_526),
.B(n_524),
.C(n_525),
.Y(n_5097)
);

AOI211xp5_ASAP7_75t_L g5098 ( 
.A1(n_5028),
.A2(n_529),
.B(n_527),
.C(n_528),
.Y(n_5098)
);

AOI311xp33_ASAP7_75t_L g5099 ( 
.A1(n_5034),
.A2(n_529),
.A3(n_527),
.B(n_528),
.C(n_530),
.Y(n_5099)
);

AOI221xp5_ASAP7_75t_L g5100 ( 
.A1(n_5003),
.A2(n_533),
.B1(n_530),
.B2(n_531),
.C(n_534),
.Y(n_5100)
);

NAND2xp5_ASAP7_75t_SL g5101 ( 
.A(n_4982),
.B(n_531),
.Y(n_5101)
);

AND2x2_ASAP7_75t_L g5102 ( 
.A(n_5053),
.B(n_536),
.Y(n_5102)
);

NOR2xp67_ASAP7_75t_L g5103 ( 
.A(n_5005),
.B(n_5040),
.Y(n_5103)
);

NOR2xp33_ASAP7_75t_L g5104 ( 
.A(n_4993),
.B(n_537),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_5023),
.Y(n_5105)
);

AOI211xp5_ASAP7_75t_SL g5106 ( 
.A1(n_5009),
.A2(n_540),
.B(n_538),
.C(n_539),
.Y(n_5106)
);

AOI22xp5_ASAP7_75t_L g5107 ( 
.A1(n_5036),
.A2(n_541),
.B1(n_539),
.B2(n_540),
.Y(n_5107)
);

OAI22xp5_ASAP7_75t_L g5108 ( 
.A1(n_4995),
.A2(n_543),
.B1(n_541),
.B2(n_542),
.Y(n_5108)
);

OAI211xp5_ASAP7_75t_L g5109 ( 
.A1(n_5029),
.A2(n_545),
.B(n_542),
.C(n_543),
.Y(n_5109)
);

NAND3xp33_ASAP7_75t_SL g5110 ( 
.A(n_5014),
.B(n_545),
.C(n_546),
.Y(n_5110)
);

O2A1O1Ixp33_ASAP7_75t_L g5111 ( 
.A1(n_5042),
.A2(n_548),
.B(n_546),
.C(n_547),
.Y(n_5111)
);

OAI211xp5_ASAP7_75t_L g5112 ( 
.A1(n_4983),
.A2(n_550),
.B(n_548),
.C(n_549),
.Y(n_5112)
);

OAI21xp5_ASAP7_75t_L g5113 ( 
.A1(n_5033),
.A2(n_549),
.B(n_552),
.Y(n_5113)
);

NOR2xp67_ASAP7_75t_L g5114 ( 
.A(n_4989),
.B(n_552),
.Y(n_5114)
);

NAND4xp25_ASAP7_75t_SL g5115 ( 
.A(n_5063),
.B(n_555),
.C(n_553),
.D(n_554),
.Y(n_5115)
);

NAND5xp2_ASAP7_75t_L g5116 ( 
.A(n_5064),
.B(n_556),
.C(n_559),
.D(n_555),
.E(n_557),
.Y(n_5116)
);

AOI221xp5_ASAP7_75t_L g5117 ( 
.A1(n_5041),
.A2(n_560),
.B1(n_554),
.B2(n_559),
.C(n_561),
.Y(n_5117)
);

AOI221xp5_ASAP7_75t_L g5118 ( 
.A1(n_5059),
.A2(n_564),
.B1(n_561),
.B2(n_562),
.C(n_565),
.Y(n_5118)
);

NAND2xp5_ASAP7_75t_SL g5119 ( 
.A(n_4990),
.B(n_564),
.Y(n_5119)
);

OAI21xp33_ASAP7_75t_L g5120 ( 
.A1(n_5022),
.A2(n_565),
.B(n_566),
.Y(n_5120)
);

OAI21xp5_ASAP7_75t_L g5121 ( 
.A1(n_5057),
.A2(n_566),
.B(n_567),
.Y(n_5121)
);

NAND2xp5_ASAP7_75t_L g5122 ( 
.A(n_5066),
.B(n_5006),
.Y(n_5122)
);

NOR3xp33_ASAP7_75t_L g5123 ( 
.A(n_5016),
.B(n_567),
.C(n_568),
.Y(n_5123)
);

AOI221xp5_ASAP7_75t_L g5124 ( 
.A1(n_5038),
.A2(n_570),
.B1(n_568),
.B2(n_569),
.C(n_571),
.Y(n_5124)
);

NAND4xp25_ASAP7_75t_L g5125 ( 
.A(n_5050),
.B(n_573),
.C(n_571),
.D(n_572),
.Y(n_5125)
);

NAND2xp5_ASAP7_75t_SL g5126 ( 
.A(n_5025),
.B(n_5037),
.Y(n_5126)
);

NOR2xp33_ASAP7_75t_R g5127 ( 
.A(n_5062),
.B(n_572),
.Y(n_5127)
);

AOI222xp33_ASAP7_75t_L g5128 ( 
.A1(n_5054),
.A2(n_575),
.B1(n_577),
.B2(n_573),
.C1(n_574),
.C2(n_576),
.Y(n_5128)
);

NAND2xp33_ASAP7_75t_R g5129 ( 
.A(n_5051),
.B(n_574),
.Y(n_5129)
);

OAI21xp5_ASAP7_75t_L g5130 ( 
.A1(n_5049),
.A2(n_576),
.B(n_577),
.Y(n_5130)
);

AOI21xp33_ASAP7_75t_SL g5131 ( 
.A1(n_5024),
.A2(n_578),
.B(n_579),
.Y(n_5131)
);

A2O1A1Ixp33_ASAP7_75t_L g5132 ( 
.A1(n_5058),
.A2(n_5010),
.B(n_5043),
.C(n_5047),
.Y(n_5132)
);

NAND4xp25_ASAP7_75t_SL g5133 ( 
.A(n_4998),
.B(n_5021),
.C(n_5055),
.D(n_5039),
.Y(n_5133)
);

O2A1O1Ixp5_ASAP7_75t_L g5134 ( 
.A1(n_5061),
.A2(n_580),
.B(n_578),
.C(n_579),
.Y(n_5134)
);

OAI22xp5_ASAP7_75t_L g5135 ( 
.A1(n_5052),
.A2(n_583),
.B1(n_580),
.B2(n_581),
.Y(n_5135)
);

AOI222xp33_ASAP7_75t_L g5136 ( 
.A1(n_4981),
.A2(n_585),
.B1(n_587),
.B2(n_581),
.C1(n_583),
.C2(n_586),
.Y(n_5136)
);

NAND3xp33_ASAP7_75t_L g5137 ( 
.A(n_4988),
.B(n_590),
.C(n_589),
.Y(n_5137)
);

AOI22xp5_ASAP7_75t_L g5138 ( 
.A1(n_4981),
.A2(n_592),
.B1(n_585),
.B2(n_591),
.Y(n_5138)
);

OAI221xp5_ASAP7_75t_L g5139 ( 
.A1(n_4988),
.A2(n_593),
.B1(n_591),
.B2(n_592),
.C(n_594),
.Y(n_5139)
);

AOI221x1_ASAP7_75t_L g5140 ( 
.A1(n_5068),
.A2(n_595),
.B1(n_593),
.B2(n_594),
.C(n_596),
.Y(n_5140)
);

NOR2xp33_ASAP7_75t_L g5141 ( 
.A(n_5056),
.B(n_595),
.Y(n_5141)
);

AOI21xp33_ASAP7_75t_L g5142 ( 
.A1(n_4981),
.A2(n_596),
.B(n_597),
.Y(n_5142)
);

NAND3xp33_ASAP7_75t_SL g5143 ( 
.A(n_4988),
.B(n_597),
.C(n_598),
.Y(n_5143)
);

OAI21xp33_ASAP7_75t_L g5144 ( 
.A1(n_4985),
.A2(n_598),
.B(n_599),
.Y(n_5144)
);

AOI21xp5_ASAP7_75t_L g5145 ( 
.A1(n_4988),
.A2(n_599),
.B(n_600),
.Y(n_5145)
);

AOI21xp5_ASAP7_75t_L g5146 ( 
.A1(n_4988),
.A2(n_600),
.B(n_601),
.Y(n_5146)
);

AOI21xp5_ASAP7_75t_L g5147 ( 
.A1(n_4988),
.A2(n_601),
.B(n_602),
.Y(n_5147)
);

NAND2xp5_ASAP7_75t_L g5148 ( 
.A(n_4985),
.B(n_602),
.Y(n_5148)
);

XNOR2x1_ASAP7_75t_L g5149 ( 
.A(n_4981),
.B(n_603),
.Y(n_5149)
);

NAND3xp33_ASAP7_75t_SL g5150 ( 
.A(n_4988),
.B(n_604),
.C(n_605),
.Y(n_5150)
);

OAI211xp5_ASAP7_75t_SL g5151 ( 
.A1(n_4988),
.A2(n_608),
.B(n_606),
.C(n_607),
.Y(n_5151)
);

AOI22xp33_ASAP7_75t_L g5152 ( 
.A1(n_5032),
.A2(n_609),
.B1(n_607),
.B2(n_608),
.Y(n_5152)
);

NAND2xp5_ASAP7_75t_L g5153 ( 
.A(n_4985),
.B(n_609),
.Y(n_5153)
);

AOI211xp5_ASAP7_75t_L g5154 ( 
.A1(n_4987),
.A2(n_612),
.B(n_610),
.C(n_611),
.Y(n_5154)
);

NAND2xp5_ASAP7_75t_L g5155 ( 
.A(n_4985),
.B(n_610),
.Y(n_5155)
);

OAI22xp5_ASAP7_75t_L g5156 ( 
.A1(n_5137),
.A2(n_614),
.B1(n_612),
.B2(n_613),
.Y(n_5156)
);

OAI21xp5_ASAP7_75t_L g5157 ( 
.A1(n_5074),
.A2(n_613),
.B(n_614),
.Y(n_5157)
);

NAND3xp33_ASAP7_75t_L g5158 ( 
.A(n_5075),
.B(n_615),
.C(n_616),
.Y(n_5158)
);

NAND3xp33_ASAP7_75t_L g5159 ( 
.A(n_5080),
.B(n_616),
.C(n_618),
.Y(n_5159)
);

OAI22xp5_ASAP7_75t_L g5160 ( 
.A1(n_5139),
.A2(n_621),
.B1(n_619),
.B2(n_620),
.Y(n_5160)
);

O2A1O1Ixp33_ASAP7_75t_L g5161 ( 
.A1(n_5143),
.A2(n_621),
.B(n_619),
.C(n_620),
.Y(n_5161)
);

AOI221xp5_ASAP7_75t_L g5162 ( 
.A1(n_5150),
.A2(n_624),
.B1(n_622),
.B2(n_623),
.C(n_625),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_SL g5163 ( 
.A(n_5076),
.B(n_624),
.Y(n_5163)
);

AOI21xp5_ASAP7_75t_L g5164 ( 
.A1(n_5145),
.A2(n_625),
.B(n_626),
.Y(n_5164)
);

OAI21xp33_ASAP7_75t_L g5165 ( 
.A1(n_5151),
.A2(n_626),
.B(n_628),
.Y(n_5165)
);

AOI211xp5_ASAP7_75t_L g5166 ( 
.A1(n_5069),
.A2(n_633),
.B(n_628),
.C(n_632),
.Y(n_5166)
);

AOI22xp33_ASAP7_75t_L g5167 ( 
.A1(n_5086),
.A2(n_634),
.B1(n_632),
.B2(n_633),
.Y(n_5167)
);

NAND3xp33_ASAP7_75t_L g5168 ( 
.A(n_5096),
.B(n_634),
.C(n_635),
.Y(n_5168)
);

AOI321xp33_ASAP7_75t_L g5169 ( 
.A1(n_5105),
.A2(n_638),
.A3(n_641),
.B1(n_635),
.B2(n_636),
.C(n_639),
.Y(n_5169)
);

NAND4xp25_ASAP7_75t_SL g5170 ( 
.A(n_5146),
.B(n_641),
.C(n_638),
.D(n_639),
.Y(n_5170)
);

AOI211xp5_ASAP7_75t_L g5171 ( 
.A1(n_5147),
.A2(n_645),
.B(n_643),
.C(n_644),
.Y(n_5171)
);

OA21x2_ASAP7_75t_L g5172 ( 
.A1(n_5148),
.A2(n_643),
.B(n_646),
.Y(n_5172)
);

AOI21xp5_ASAP7_75t_L g5173 ( 
.A1(n_5092),
.A2(n_647),
.B(n_649),
.Y(n_5173)
);

AOI221xp5_ASAP7_75t_L g5174 ( 
.A1(n_5133),
.A2(n_650),
.B1(n_647),
.B2(n_649),
.C(n_651),
.Y(n_5174)
);

NAND2xp5_ASAP7_75t_L g5175 ( 
.A(n_5094),
.B(n_5106),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_L g5176 ( 
.A(n_5141),
.B(n_652),
.Y(n_5176)
);

INVx2_ASAP7_75t_L g5177 ( 
.A(n_5149),
.Y(n_5177)
);

NOR3x1_ASAP7_75t_L g5178 ( 
.A(n_5077),
.B(n_659),
.C(n_651),
.Y(n_5178)
);

AOI311xp33_ASAP7_75t_L g5179 ( 
.A1(n_5098),
.A2(n_654),
.A3(n_652),
.B(n_653),
.C(n_655),
.Y(n_5179)
);

OAI21xp5_ASAP7_75t_L g5180 ( 
.A1(n_5103),
.A2(n_655),
.B(n_656),
.Y(n_5180)
);

NOR4xp25_ASAP7_75t_SL g5181 ( 
.A(n_5129),
.B(n_659),
.C(n_657),
.D(n_658),
.Y(n_5181)
);

NOR4xp25_ASAP7_75t_L g5182 ( 
.A(n_5132),
.B(n_5082),
.C(n_5122),
.D(n_5126),
.Y(n_5182)
);

AOI21xp33_ASAP7_75t_SL g5183 ( 
.A1(n_5079),
.A2(n_660),
.B(n_661),
.Y(n_5183)
);

NOR3xp33_ASAP7_75t_L g5184 ( 
.A(n_5153),
.B(n_663),
.C(n_664),
.Y(n_5184)
);

OAI21xp33_ASAP7_75t_L g5185 ( 
.A1(n_5155),
.A2(n_663),
.B(n_664),
.Y(n_5185)
);

AOI21xp5_ASAP7_75t_L g5186 ( 
.A1(n_5072),
.A2(n_665),
.B(n_666),
.Y(n_5186)
);

AOI21xp5_ASAP7_75t_L g5187 ( 
.A1(n_5084),
.A2(n_5144),
.B(n_5108),
.Y(n_5187)
);

NAND3xp33_ASAP7_75t_L g5188 ( 
.A(n_5123),
.B(n_667),
.C(n_668),
.Y(n_5188)
);

O2A1O1Ixp33_ASAP7_75t_L g5189 ( 
.A1(n_5111),
.A2(n_672),
.B(n_669),
.C(n_670),
.Y(n_5189)
);

OAI21xp5_ASAP7_75t_L g5190 ( 
.A1(n_5134),
.A2(n_670),
.B(n_673),
.Y(n_5190)
);

O2A1O1Ixp33_ASAP7_75t_SL g5191 ( 
.A1(n_5154),
.A2(n_676),
.B(n_673),
.C(n_674),
.Y(n_5191)
);

OAI21xp5_ASAP7_75t_SL g5192 ( 
.A1(n_5112),
.A2(n_674),
.B(n_677),
.Y(n_5192)
);

CKINVDCx14_ASAP7_75t_R g5193 ( 
.A(n_5127),
.Y(n_5193)
);

A2O1A1Ixp33_ASAP7_75t_L g5194 ( 
.A1(n_5097),
.A2(n_679),
.B(n_677),
.C(n_678),
.Y(n_5194)
);

NAND3xp33_ASAP7_75t_SL g5195 ( 
.A(n_5091),
.B(n_680),
.C(n_681),
.Y(n_5195)
);

NOR2xp33_ASAP7_75t_L g5196 ( 
.A(n_5116),
.B(n_680),
.Y(n_5196)
);

AOI221x1_ASAP7_75t_L g5197 ( 
.A1(n_5081),
.A2(n_683),
.B1(n_681),
.B2(n_682),
.C(n_684),
.Y(n_5197)
);

AOI22xp33_ASAP7_75t_L g5198 ( 
.A1(n_5114),
.A2(n_685),
.B1(n_682),
.B2(n_684),
.Y(n_5198)
);

NOR2xp33_ASAP7_75t_SL g5199 ( 
.A(n_5095),
.B(n_685),
.Y(n_5199)
);

NOR2xp33_ASAP7_75t_L g5200 ( 
.A(n_5078),
.B(n_686),
.Y(n_5200)
);

A2O1A1Ixp33_ASAP7_75t_L g5201 ( 
.A1(n_5088),
.A2(n_688),
.B(n_686),
.C(n_687),
.Y(n_5201)
);

NOR2xp33_ASAP7_75t_SL g5202 ( 
.A(n_5125),
.B(n_687),
.Y(n_5202)
);

NAND3xp33_ASAP7_75t_SL g5203 ( 
.A(n_5131),
.B(n_688),
.C(n_689),
.Y(n_5203)
);

AOI22xp5_ASAP7_75t_L g5204 ( 
.A1(n_5104),
.A2(n_692),
.B1(n_690),
.B2(n_691),
.Y(n_5204)
);

AOI211xp5_ASAP7_75t_L g5205 ( 
.A1(n_5109),
.A2(n_694),
.B(n_690),
.C(n_693),
.Y(n_5205)
);

HB1xp67_ASAP7_75t_L g5206 ( 
.A(n_5073),
.Y(n_5206)
);

NAND3xp33_ASAP7_75t_SL g5207 ( 
.A(n_5128),
.B(n_693),
.C(n_694),
.Y(n_5207)
);

NOR2xp33_ASAP7_75t_L g5208 ( 
.A(n_5110),
.B(n_695),
.Y(n_5208)
);

NAND4xp25_ASAP7_75t_SL g5209 ( 
.A(n_5136),
.B(n_698),
.C(n_696),
.D(n_697),
.Y(n_5209)
);

AOI211x1_ASAP7_75t_SL g5210 ( 
.A1(n_5121),
.A2(n_699),
.B(n_697),
.C(n_698),
.Y(n_5210)
);

OAI21xp5_ASAP7_75t_SL g5211 ( 
.A1(n_5089),
.A2(n_700),
.B(n_701),
.Y(n_5211)
);

NAND4xp25_ASAP7_75t_L g5212 ( 
.A(n_5099),
.B(n_704),
.C(n_702),
.D(n_703),
.Y(n_5212)
);

AOI211xp5_ASAP7_75t_SL g5213 ( 
.A1(n_5142),
.A2(n_705),
.B(n_703),
.C(n_704),
.Y(n_5213)
);

AOI21xp5_ASAP7_75t_L g5214 ( 
.A1(n_5101),
.A2(n_705),
.B(n_706),
.Y(n_5214)
);

OAI211xp5_ASAP7_75t_SL g5215 ( 
.A1(n_5100),
.A2(n_709),
.B(n_707),
.C(n_708),
.Y(n_5215)
);

NAND2xp5_ASAP7_75t_L g5216 ( 
.A(n_5102),
.B(n_708),
.Y(n_5216)
);

AOI221xp5_ASAP7_75t_L g5217 ( 
.A1(n_5090),
.A2(n_710),
.B1(n_707),
.B2(n_709),
.C(n_711),
.Y(n_5217)
);

NOR2xp33_ASAP7_75t_L g5218 ( 
.A(n_5087),
.B(n_5119),
.Y(n_5218)
);

AOI221xp5_ASAP7_75t_L g5219 ( 
.A1(n_5130),
.A2(n_712),
.B1(n_710),
.B2(n_711),
.C(n_713),
.Y(n_5219)
);

NOR2x1_ASAP7_75t_L g5220 ( 
.A(n_5135),
.B(n_712),
.Y(n_5220)
);

OAI221xp5_ASAP7_75t_L g5221 ( 
.A1(n_5113),
.A2(n_715),
.B1(n_713),
.B2(n_714),
.C(n_716),
.Y(n_5221)
);

AOI21x1_ASAP7_75t_L g5222 ( 
.A1(n_5140),
.A2(n_714),
.B(n_715),
.Y(n_5222)
);

AOI21xp5_ASAP7_75t_L g5223 ( 
.A1(n_5124),
.A2(n_716),
.B(n_717),
.Y(n_5223)
);

NOR4xp25_ASAP7_75t_L g5224 ( 
.A(n_5120),
.B(n_720),
.C(n_718),
.D(n_719),
.Y(n_5224)
);

INVx1_ASAP7_75t_L g5225 ( 
.A(n_5070),
.Y(n_5225)
);

AOI221xp5_ASAP7_75t_L g5226 ( 
.A1(n_5115),
.A2(n_5085),
.B1(n_5093),
.B2(n_5118),
.C(n_5117),
.Y(n_5226)
);

NOR2xp33_ASAP7_75t_L g5227 ( 
.A(n_5138),
.B(n_719),
.Y(n_5227)
);

OAI221xp5_ASAP7_75t_L g5228 ( 
.A1(n_5071),
.A2(n_722),
.B1(n_720),
.B2(n_721),
.C(n_723),
.Y(n_5228)
);

NAND3xp33_ASAP7_75t_SL g5229 ( 
.A(n_5152),
.B(n_722),
.C(n_725),
.Y(n_5229)
);

NAND2xp5_ASAP7_75t_SL g5230 ( 
.A(n_5083),
.B(n_726),
.Y(n_5230)
);

AOI211xp5_ASAP7_75t_L g5231 ( 
.A1(n_5107),
.A2(n_729),
.B(n_727),
.C(n_728),
.Y(n_5231)
);

AOI221xp5_ASAP7_75t_L g5232 ( 
.A1(n_5074),
.A2(n_730),
.B1(n_727),
.B2(n_729),
.C(n_732),
.Y(n_5232)
);

A2O1A1Ixp33_ASAP7_75t_L g5233 ( 
.A1(n_5227),
.A2(n_733),
.B(n_730),
.C(n_732),
.Y(n_5233)
);

AOI21xp5_ASAP7_75t_L g5234 ( 
.A1(n_5175),
.A2(n_734),
.B(n_735),
.Y(n_5234)
);

NAND2xp5_ASAP7_75t_L g5235 ( 
.A(n_5210),
.B(n_734),
.Y(n_5235)
);

XOR2xp5_ASAP7_75t_L g5236 ( 
.A(n_5193),
.B(n_735),
.Y(n_5236)
);

AOI211xp5_ASAP7_75t_L g5237 ( 
.A1(n_5212),
.A2(n_739),
.B(n_741),
.C(n_737),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_L g5238 ( 
.A(n_5196),
.B(n_736),
.Y(n_5238)
);

O2A1O1Ixp33_ASAP7_75t_L g5239 ( 
.A1(n_5163),
.A2(n_742),
.B(n_737),
.C(n_739),
.Y(n_5239)
);

AOI211xp5_ASAP7_75t_L g5240 ( 
.A1(n_5209),
.A2(n_744),
.B(n_745),
.C(n_743),
.Y(n_5240)
);

AOI211xp5_ASAP7_75t_L g5241 ( 
.A1(n_5157),
.A2(n_747),
.B(n_748),
.C(n_746),
.Y(n_5241)
);

AOI311xp33_ASAP7_75t_L g5242 ( 
.A1(n_5225),
.A2(n_763),
.A3(n_771),
.B(n_755),
.C(n_742),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_5222),
.Y(n_5243)
);

OAI211xp5_ASAP7_75t_L g5244 ( 
.A1(n_5182),
.A2(n_750),
.B(n_746),
.C(n_747),
.Y(n_5244)
);

AOI221xp5_ASAP7_75t_L g5245 ( 
.A1(n_5173),
.A2(n_753),
.B1(n_751),
.B2(n_752),
.C(n_754),
.Y(n_5245)
);

OAI22xp33_ASAP7_75t_L g5246 ( 
.A1(n_5216),
.A2(n_755),
.B1(n_752),
.B2(n_753),
.Y(n_5246)
);

OAI211xp5_ASAP7_75t_SL g5247 ( 
.A1(n_5177),
.A2(n_758),
.B(n_756),
.C(n_757),
.Y(n_5247)
);

NOR2x1_ASAP7_75t_L g5248 ( 
.A(n_5159),
.B(n_756),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_5172),
.Y(n_5249)
);

OAI221xp5_ASAP7_75t_L g5250 ( 
.A1(n_5180),
.A2(n_759),
.B1(n_757),
.B2(n_758),
.C(n_760),
.Y(n_5250)
);

AOI21xp5_ASAP7_75t_SL g5251 ( 
.A1(n_5161),
.A2(n_759),
.B(n_761),
.Y(n_5251)
);

AOI211xp5_ASAP7_75t_L g5252 ( 
.A1(n_5170),
.A2(n_765),
.B(n_766),
.C(n_764),
.Y(n_5252)
);

AOI222xp33_ASAP7_75t_L g5253 ( 
.A1(n_5207),
.A2(n_768),
.B1(n_770),
.B2(n_762),
.C1(n_767),
.C2(n_769),
.Y(n_5253)
);

NAND4xp25_ASAP7_75t_L g5254 ( 
.A(n_5179),
.B(n_769),
.C(n_762),
.D(n_767),
.Y(n_5254)
);

NOR4xp25_ASAP7_75t_L g5255 ( 
.A(n_5158),
.B(n_5192),
.C(n_5195),
.D(n_5211),
.Y(n_5255)
);

AOI21xp5_ASAP7_75t_L g5256 ( 
.A1(n_5191),
.A2(n_770),
.B(n_771),
.Y(n_5256)
);

AND2x2_ASAP7_75t_L g5257 ( 
.A(n_5178),
.B(n_772),
.Y(n_5257)
);

NAND3xp33_ASAP7_75t_L g5258 ( 
.A(n_5168),
.B(n_773),
.C(n_774),
.Y(n_5258)
);

AOI22xp33_ASAP7_75t_L g5259 ( 
.A1(n_5206),
.A2(n_776),
.B1(n_774),
.B2(n_775),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_SL g5260 ( 
.A(n_5169),
.B(n_775),
.Y(n_5260)
);

O2A1O1Ixp33_ASAP7_75t_L g5261 ( 
.A1(n_5176),
.A2(n_778),
.B(n_776),
.C(n_777),
.Y(n_5261)
);

NOR2x1_ASAP7_75t_L g5262 ( 
.A(n_5221),
.B(n_777),
.Y(n_5262)
);

AOI221x1_ASAP7_75t_L g5263 ( 
.A1(n_5223),
.A2(n_780),
.B1(n_778),
.B2(n_779),
.C(n_781),
.Y(n_5263)
);

AOI222xp33_ASAP7_75t_L g5264 ( 
.A1(n_5203),
.A2(n_784),
.B1(n_786),
.B2(n_780),
.C1(n_783),
.C2(n_785),
.Y(n_5264)
);

AOI211xp5_ASAP7_75t_SL g5265 ( 
.A1(n_5200),
.A2(n_786),
.B(n_783),
.C(n_785),
.Y(n_5265)
);

AOI211xp5_ASAP7_75t_L g5266 ( 
.A1(n_5160),
.A2(n_789),
.B(n_790),
.C(n_788),
.Y(n_5266)
);

AOI211xp5_ASAP7_75t_SL g5267 ( 
.A1(n_5208),
.A2(n_789),
.B(n_787),
.C(n_788),
.Y(n_5267)
);

OAI221xp5_ASAP7_75t_L g5268 ( 
.A1(n_5162),
.A2(n_793),
.B1(n_791),
.B2(n_792),
.C(n_794),
.Y(n_5268)
);

AOI21xp5_ASAP7_75t_L g5269 ( 
.A1(n_5232),
.A2(n_793),
.B(n_794),
.Y(n_5269)
);

NAND4xp25_ASAP7_75t_L g5270 ( 
.A(n_5202),
.B(n_797),
.C(n_795),
.D(n_796),
.Y(n_5270)
);

NAND2xp5_ASAP7_75t_L g5271 ( 
.A(n_5213),
.B(n_795),
.Y(n_5271)
);

NOR3x1_ASAP7_75t_L g5272 ( 
.A(n_5228),
.B(n_796),
.C(n_797),
.Y(n_5272)
);

AOI221x1_ASAP7_75t_L g5273 ( 
.A1(n_5214),
.A2(n_800),
.B1(n_798),
.B2(n_799),
.C(n_801),
.Y(n_5273)
);

O2A1O1Ixp33_ASAP7_75t_L g5274 ( 
.A1(n_5194),
.A2(n_802),
.B(n_798),
.C(n_799),
.Y(n_5274)
);

AOI21xp5_ASAP7_75t_L g5275 ( 
.A1(n_5174),
.A2(n_802),
.B(n_803),
.Y(n_5275)
);

AOI221x1_ASAP7_75t_L g5276 ( 
.A1(n_5186),
.A2(n_805),
.B1(n_803),
.B2(n_804),
.C(n_807),
.Y(n_5276)
);

OAI221xp5_ASAP7_75t_SL g5277 ( 
.A1(n_5165),
.A2(n_809),
.B1(n_812),
.B2(n_808),
.C(n_810),
.Y(n_5277)
);

AND2x2_ASAP7_75t_L g5278 ( 
.A(n_5190),
.B(n_804),
.Y(n_5278)
);

AOI211xp5_ASAP7_75t_SL g5279 ( 
.A1(n_5164),
.A2(n_5218),
.B(n_5199),
.C(n_5156),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_L g5280 ( 
.A(n_5224),
.B(n_808),
.Y(n_5280)
);

OAI211xp5_ASAP7_75t_L g5281 ( 
.A1(n_5171),
.A2(n_813),
.B(n_809),
.C(n_812),
.Y(n_5281)
);

AOI21xp5_ASAP7_75t_L g5282 ( 
.A1(n_5230),
.A2(n_5189),
.B(n_5187),
.Y(n_5282)
);

AOI221xp5_ASAP7_75t_L g5283 ( 
.A1(n_5226),
.A2(n_815),
.B1(n_813),
.B2(n_814),
.C(n_816),
.Y(n_5283)
);

AOI22xp5_ASAP7_75t_L g5284 ( 
.A1(n_5184),
.A2(n_816),
.B1(n_814),
.B2(n_815),
.Y(n_5284)
);

OAI211xp5_ASAP7_75t_SL g5285 ( 
.A1(n_5220),
.A2(n_819),
.B(n_817),
.C(n_818),
.Y(n_5285)
);

NOR4xp25_ASAP7_75t_L g5286 ( 
.A(n_5185),
.B(n_821),
.C(n_817),
.D(n_820),
.Y(n_5286)
);

OAI211xp5_ASAP7_75t_SL g5287 ( 
.A1(n_5166),
.A2(n_822),
.B(n_820),
.C(n_821),
.Y(n_5287)
);

AOI211xp5_ASAP7_75t_SL g5288 ( 
.A1(n_5229),
.A2(n_824),
.B(n_822),
.C(n_823),
.Y(n_5288)
);

NOR2x1_ASAP7_75t_L g5289 ( 
.A(n_5243),
.B(n_5188),
.Y(n_5289)
);

NOR2xp33_ASAP7_75t_L g5290 ( 
.A(n_5285),
.B(n_5172),
.Y(n_5290)
);

NOR4xp75_ASAP7_75t_L g5291 ( 
.A(n_5260),
.B(n_5181),
.C(n_5183),
.D(n_5205),
.Y(n_5291)
);

NAND3xp33_ASAP7_75t_L g5292 ( 
.A(n_5249),
.B(n_5198),
.C(n_5167),
.Y(n_5292)
);

NOR2x1_ASAP7_75t_L g5293 ( 
.A(n_5244),
.B(n_5201),
.Y(n_5293)
);

INVx2_ASAP7_75t_L g5294 ( 
.A(n_5257),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_5256),
.B(n_5197),
.Y(n_5295)
);

NOR3xp33_ASAP7_75t_L g5296 ( 
.A(n_5238),
.B(n_5270),
.C(n_5271),
.Y(n_5296)
);

NOR2xp67_ASAP7_75t_L g5297 ( 
.A(n_5254),
.B(n_5204),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_5236),
.Y(n_5298)
);

NOR2xp67_ASAP7_75t_L g5299 ( 
.A(n_5250),
.B(n_5231),
.Y(n_5299)
);

INVx2_ASAP7_75t_L g5300 ( 
.A(n_5278),
.Y(n_5300)
);

OAI22xp5_ASAP7_75t_SL g5301 ( 
.A1(n_5235),
.A2(n_5219),
.B1(n_5215),
.B2(n_5217),
.Y(n_5301)
);

OAI22xp5_ASAP7_75t_SL g5302 ( 
.A1(n_5280),
.A2(n_827),
.B1(n_823),
.B2(n_826),
.Y(n_5302)
);

NOR3xp33_ASAP7_75t_SL g5303 ( 
.A(n_5282),
.B(n_826),
.C(n_827),
.Y(n_5303)
);

NAND2xp33_ASAP7_75t_L g5304 ( 
.A(n_5242),
.B(n_828),
.Y(n_5304)
);

NOR2x1_ASAP7_75t_L g5305 ( 
.A(n_5234),
.B(n_829),
.Y(n_5305)
);

NAND4xp75_ASAP7_75t_L g5306 ( 
.A(n_5248),
.B(n_832),
.C(n_830),
.D(n_831),
.Y(n_5306)
);

OAI211xp5_ASAP7_75t_L g5307 ( 
.A1(n_5264),
.A2(n_832),
.B(n_830),
.C(n_831),
.Y(n_5307)
);

AO22x2_ASAP7_75t_L g5308 ( 
.A1(n_5276),
.A2(n_835),
.B1(n_833),
.B2(n_834),
.Y(n_5308)
);

AND2x2_ASAP7_75t_L g5309 ( 
.A(n_5237),
.B(n_834),
.Y(n_5309)
);

NAND4xp25_ASAP7_75t_L g5310 ( 
.A(n_5265),
.B(n_837),
.C(n_835),
.D(n_836),
.Y(n_5310)
);

AOI22xp5_ASAP7_75t_L g5311 ( 
.A1(n_5262),
.A2(n_839),
.B1(n_836),
.B2(n_838),
.Y(n_5311)
);

OR2x2_ASAP7_75t_L g5312 ( 
.A(n_5286),
.B(n_838),
.Y(n_5312)
);

BUFx4_ASAP7_75t_R g5313 ( 
.A(n_5255),
.Y(n_5313)
);

AND2x2_ASAP7_75t_SL g5314 ( 
.A(n_5272),
.B(n_839),
.Y(n_5314)
);

NOR3xp33_ASAP7_75t_L g5315 ( 
.A(n_5246),
.B(n_840),
.C(n_841),
.Y(n_5315)
);

NAND3xp33_ASAP7_75t_L g5316 ( 
.A(n_5267),
.B(n_841),
.C(n_842),
.Y(n_5316)
);

NOR3xp33_ASAP7_75t_L g5317 ( 
.A(n_5261),
.B(n_842),
.C(n_843),
.Y(n_5317)
);

INVxp67_ASAP7_75t_SL g5318 ( 
.A(n_5239),
.Y(n_5318)
);

NAND4xp25_ASAP7_75t_L g5319 ( 
.A(n_5288),
.B(n_845),
.C(n_843),
.D(n_844),
.Y(n_5319)
);

NAND4xp75_ASAP7_75t_L g5320 ( 
.A(n_5263),
.B(n_848),
.C(n_846),
.D(n_847),
.Y(n_5320)
);

NOR3xp33_ASAP7_75t_L g5321 ( 
.A(n_5247),
.B(n_846),
.C(n_849),
.Y(n_5321)
);

NOR3xp33_ASAP7_75t_L g5322 ( 
.A(n_5283),
.B(n_849),
.C(n_850),
.Y(n_5322)
);

INVx1_ASAP7_75t_L g5323 ( 
.A(n_5273),
.Y(n_5323)
);

NOR2x1_ASAP7_75t_L g5324 ( 
.A(n_5289),
.B(n_5251),
.Y(n_5324)
);

NAND4xp75_ASAP7_75t_L g5325 ( 
.A(n_5298),
.B(n_5275),
.C(n_5269),
.D(n_5245),
.Y(n_5325)
);

NOR3xp33_ASAP7_75t_L g5326 ( 
.A(n_5294),
.B(n_5281),
.C(n_5258),
.Y(n_5326)
);

NAND2x1p5_ASAP7_75t_L g5327 ( 
.A(n_5323),
.B(n_5305),
.Y(n_5327)
);

AND2x2_ASAP7_75t_L g5328 ( 
.A(n_5303),
.B(n_5253),
.Y(n_5328)
);

OR2x2_ASAP7_75t_L g5329 ( 
.A(n_5310),
.B(n_5277),
.Y(n_5329)
);

AND3x4_ASAP7_75t_L g5330 ( 
.A(n_5291),
.B(n_5279),
.C(n_5240),
.Y(n_5330)
);

NOR3xp33_ASAP7_75t_L g5331 ( 
.A(n_5300),
.B(n_5292),
.C(n_5302),
.Y(n_5331)
);

NOR2x1_ASAP7_75t_L g5332 ( 
.A(n_5304),
.B(n_5233),
.Y(n_5332)
);

AND2x2_ASAP7_75t_L g5333 ( 
.A(n_5309),
.B(n_5252),
.Y(n_5333)
);

AND2x4_ASAP7_75t_L g5334 ( 
.A(n_5318),
.B(n_5284),
.Y(n_5334)
);

NAND2xp5_ASAP7_75t_L g5335 ( 
.A(n_5314),
.B(n_5241),
.Y(n_5335)
);

NOR2x1_ASAP7_75t_L g5336 ( 
.A(n_5312),
.B(n_5287),
.Y(n_5336)
);

NAND2xp5_ASAP7_75t_L g5337 ( 
.A(n_5290),
.B(n_5259),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_5308),
.Y(n_5338)
);

NAND2xp33_ASAP7_75t_L g5339 ( 
.A(n_5317),
.B(n_5268),
.Y(n_5339)
);

NOR2x1_ASAP7_75t_L g5340 ( 
.A(n_5306),
.B(n_5274),
.Y(n_5340)
);

INVx2_ASAP7_75t_L g5341 ( 
.A(n_5327),
.Y(n_5341)
);

OAI21xp5_ASAP7_75t_SL g5342 ( 
.A1(n_5324),
.A2(n_5311),
.B(n_5307),
.Y(n_5342)
);

OR2x2_ASAP7_75t_L g5343 ( 
.A(n_5338),
.B(n_5319),
.Y(n_5343)
);

NAND4xp75_ASAP7_75t_L g5344 ( 
.A(n_5332),
.B(n_5293),
.C(n_5297),
.D(n_5295),
.Y(n_5344)
);

NAND2xp5_ASAP7_75t_L g5345 ( 
.A(n_5336),
.B(n_5308),
.Y(n_5345)
);

AND2x2_ASAP7_75t_SL g5346 ( 
.A(n_5331),
.B(n_5326),
.Y(n_5346)
);

AND2x4_ASAP7_75t_L g5347 ( 
.A(n_5334),
.B(n_5296),
.Y(n_5347)
);

NAND2x1_ASAP7_75t_L g5348 ( 
.A(n_5328),
.B(n_5316),
.Y(n_5348)
);

NAND3xp33_ASAP7_75t_SL g5349 ( 
.A(n_5330),
.B(n_5315),
.C(n_5266),
.Y(n_5349)
);

OAI221xp5_ASAP7_75t_SL g5350 ( 
.A1(n_5337),
.A2(n_5322),
.B1(n_5321),
.B2(n_5313),
.C(n_5320),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_5335),
.Y(n_5351)
);

NAND3xp33_ASAP7_75t_L g5352 ( 
.A(n_5341),
.B(n_5339),
.C(n_5333),
.Y(n_5352)
);

NAND3xp33_ASAP7_75t_L g5353 ( 
.A(n_5345),
.B(n_5340),
.C(n_5329),
.Y(n_5353)
);

NOR2xp33_ASAP7_75t_R g5354 ( 
.A(n_5349),
.B(n_850),
.Y(n_5354)
);

NOR2xp33_ASAP7_75t_R g5355 ( 
.A(n_5346),
.B(n_851),
.Y(n_5355)
);

NAND2xp33_ASAP7_75t_SL g5356 ( 
.A(n_5343),
.B(n_5301),
.Y(n_5356)
);

NAND3xp33_ASAP7_75t_L g5357 ( 
.A(n_5348),
.B(n_5299),
.C(n_5325),
.Y(n_5357)
);

NOR2xp33_ASAP7_75t_R g5358 ( 
.A(n_5351),
.B(n_851),
.Y(n_5358)
);

INVx1_ASAP7_75t_L g5359 ( 
.A(n_5357),
.Y(n_5359)
);

INVx1_ASAP7_75t_L g5360 ( 
.A(n_5352),
.Y(n_5360)
);

INVx2_ASAP7_75t_L g5361 ( 
.A(n_5353),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_5355),
.Y(n_5362)
);

OA22x2_ASAP7_75t_L g5363 ( 
.A1(n_5356),
.A2(n_5342),
.B1(n_5347),
.B2(n_5344),
.Y(n_5363)
);

INVx2_ASAP7_75t_L g5364 ( 
.A(n_5361),
.Y(n_5364)
);

AOI22xp5_ASAP7_75t_L g5365 ( 
.A1(n_5360),
.A2(n_5354),
.B1(n_5350),
.B2(n_5358),
.Y(n_5365)
);

INVx1_ASAP7_75t_L g5366 ( 
.A(n_5364),
.Y(n_5366)
);

XNOR2xp5_ASAP7_75t_L g5367 ( 
.A(n_5366),
.B(n_5363),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_5367),
.Y(n_5368)
);

OAI211xp5_ASAP7_75t_L g5369 ( 
.A1(n_5368),
.A2(n_5365),
.B(n_5359),
.C(n_5362),
.Y(n_5369)
);

OAI322xp33_ASAP7_75t_L g5370 ( 
.A1(n_5369),
.A2(n_858),
.A3(n_856),
.B1(n_854),
.B2(n_852),
.C1(n_853),
.C2(n_855),
.Y(n_5370)
);

AOI21xp33_ASAP7_75t_L g5371 ( 
.A1(n_5370),
.A2(n_854),
.B(n_855),
.Y(n_5371)
);

NAND2xp5_ASAP7_75t_L g5372 ( 
.A(n_5370),
.B(n_856),
.Y(n_5372)
);

OA21x2_ASAP7_75t_L g5373 ( 
.A1(n_5372),
.A2(n_859),
.B(n_860),
.Y(n_5373)
);

OAI21xp5_ASAP7_75t_SL g5374 ( 
.A1(n_5371),
.A2(n_861),
.B(n_862),
.Y(n_5374)
);

OAI321xp33_ASAP7_75t_L g5375 ( 
.A1(n_5373),
.A2(n_863),
.A3(n_865),
.B1(n_861),
.B2(n_862),
.C(n_864),
.Y(n_5375)
);

NAND2xp5_ASAP7_75t_L g5376 ( 
.A(n_5375),
.B(n_5374),
.Y(n_5376)
);

AOI21xp5_ASAP7_75t_L g5377 ( 
.A1(n_5376),
.A2(n_865),
.B(n_866),
.Y(n_5377)
);

AOI211xp5_ASAP7_75t_L g5378 ( 
.A1(n_5377),
.A2(n_869),
.B(n_867),
.C(n_868),
.Y(n_5378)
);


endmodule