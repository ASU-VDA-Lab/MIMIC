module fake_ariane_1628_n_1810 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_410, n_379, n_445, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_439, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_413, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_257, n_148, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_430, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_425, n_431, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_1810);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_410;
input n_379;
input n_445;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_439;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_413;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_430;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_425;
input n_431;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_1810;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_995;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_1751;
wire n_533;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1396;
wire n_1230;
wire n_612;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_1716;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_489;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1674;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_1467;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1208;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_1521;
wire n_1694;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_519;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_1687;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_765;
wire n_1809;
wire n_1268;
wire n_917;
wire n_1271;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1344;
wire n_1390;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_954;
wire n_596;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_1063;
wire n_537;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_946;
wire n_757;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_1569;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_849;
wire n_1251;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g448 ( 
.A(n_93),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_112),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_186),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_155),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_199),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_55),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_217),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_387),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_147),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_3),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_430),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_304),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_433),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_32),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_446),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_59),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_174),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_417),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_428),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_398),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_116),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_203),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_109),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_343),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_333),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_291),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_272),
.Y(n_474)
);

CKINVDCx11_ASAP7_75t_R g475 ( 
.A(n_172),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_231),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_271),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_122),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_330),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_286),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_437),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_440),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_424),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_225),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_146),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_184),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_423),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_382),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_405),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_245),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_289),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_404),
.Y(n_492)
);

INVx4_ASAP7_75t_R g493 ( 
.A(n_264),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_420),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_43),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_24),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_345),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_431),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_388),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_27),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_67),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_92),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_39),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_12),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_160),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_157),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_323),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_419),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_152),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_37),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_51),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_110),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_88),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_212),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_332),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_435),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_159),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_391),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_364),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_246),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_299),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_270),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_305),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_261),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_142),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_15),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_86),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_281),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_406),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_403),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_17),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_68),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_294),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_22),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_421),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_196),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_243),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_383),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_341),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_111),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_182),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_42),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_130),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_18),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_368),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_377),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_19),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_150),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_170),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_61),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_280),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_273),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_413),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_63),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_434),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_279),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_237),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_293),
.Y(n_559)
);

BUFx10_ASAP7_75t_L g560 ( 
.A(n_211),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_251),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_426),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_357),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_65),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_319),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_6),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_379),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_429),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_17),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_392),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_60),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_353),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_267),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_168),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_44),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_136),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_325),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_104),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_432),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_165),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_311),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_176),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_19),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_194),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_49),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_409),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_25),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_32),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_355),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_167),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_188),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_306),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_354),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_401),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_439),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_198),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_162),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_81),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_54),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_381),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_375),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_55),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_197),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_94),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_436),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_39),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_438),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_64),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_258),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_277),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_300),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_324),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_7),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_260),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_284),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_295),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_40),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_2),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_117),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_69),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_76),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_427),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_500),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_500),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_495),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_548),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_569),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_583),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_587),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_618),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_544),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_517),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_496),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_546),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_461),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_560),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_560),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_475),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_578),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_453),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_448),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_452),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_458),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_462),
.Y(n_644)
);

CKINVDCx16_ASAP7_75t_R g645 ( 
.A(n_489),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_465),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_476),
.Y(n_647)
);

CKINVDCx16_ASAP7_75t_R g648 ( 
.A(n_520),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_468),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_486),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_517),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_530),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_473),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_483),
.Y(n_654)
);

INVx1_ASAP7_75t_SL g655 ( 
.A(n_599),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_488),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_530),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_502),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_490),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_554),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_507),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_578),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_578),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_513),
.Y(n_664)
);

CKINVDCx16_ASAP7_75t_R g665 ( 
.A(n_525),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_523),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_491),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_492),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_457),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_536),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_494),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_540),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_554),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_497),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_501),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_508),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_509),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_547),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_519),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_527),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_529),
.Y(n_681)
);

INVxp67_ASAP7_75t_SL g682 ( 
.A(n_557),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_539),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_503),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_542),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_622),
.B(n_0),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_551),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_556),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_557),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_563),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_580),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_572),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_581),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_582),
.Y(n_694)
);

INVxp67_ASAP7_75t_SL g695 ( 
.A(n_593),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_586),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_593),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_597),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_578),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_589),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_504),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_592),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_591),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_595),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_598),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_604),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_597),
.Y(n_707)
);

INVxp67_ASAP7_75t_SL g708 ( 
.A(n_449),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_615),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_621),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_510),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_526),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_532),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_605),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_535),
.Y(n_715)
);

NOR2xp67_ASAP7_75t_L g716 ( 
.A(n_543),
.B(n_0),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_545),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_566),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_575),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_585),
.Y(n_720)
);

INVxp33_ASAP7_75t_SL g721 ( 
.A(n_588),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_602),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_606),
.Y(n_723)
);

OA21x2_ASAP7_75t_L g724 ( 
.A1(n_641),
.A2(n_594),
.B(n_449),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_655),
.B(n_613),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_645),
.B(n_594),
.Y(n_726)
);

INVx5_ASAP7_75t_L g727 ( 
.A(n_639),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_636),
.B(n_600),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_635),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_635),
.Y(n_730)
);

INVx5_ASAP7_75t_L g731 ( 
.A(n_639),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_639),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_662),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_647),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_662),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_682),
.B(n_474),
.Y(n_736)
);

OA21x2_ASAP7_75t_L g737 ( 
.A1(n_642),
.A2(n_601),
.B(n_600),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_662),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_682),
.B(n_608),
.Y(n_739)
);

INVx5_ASAP7_75t_L g740 ( 
.A(n_663),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_663),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_712),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_663),
.Y(n_743)
);

INVx6_ASAP7_75t_L g744 ( 
.A(n_648),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_699),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_695),
.B(n_601),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_699),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_625),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_699),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_632),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_643),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_651),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_652),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_626),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_660),
.Y(n_755)
);

OAI21x1_ASAP7_75t_L g756 ( 
.A1(n_644),
.A2(n_499),
.B(n_481),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_695),
.B(n_518),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_650),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_673),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_637),
.B(n_522),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_634),
.B(n_562),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_657),
.B(n_479),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_689),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_697),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_627),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_698),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_707),
.Y(n_767)
);

BUFx8_ASAP7_75t_L g768 ( 
.A(n_630),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_665),
.A2(n_511),
.B1(n_617),
.B2(n_541),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_623),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_684),
.B(n_450),
.Y(n_771)
);

AND2x2_ASAP7_75t_SL g772 ( 
.A(n_686),
.B(n_669),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_SL g773 ( 
.A(n_655),
.B(n_638),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_624),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_646),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_711),
.B(n_451),
.Y(n_776)
);

CKINVDCx6p67_ASAP7_75t_R g777 ( 
.A(n_664),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_628),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_649),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_629),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_653),
.Y(n_781)
);

OA21x2_ASAP7_75t_L g782 ( 
.A1(n_654),
.A2(n_455),
.B(n_454),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_633),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_656),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_631),
.B(n_456),
.Y(n_785)
);

INVxp33_ASAP7_75t_SL g786 ( 
.A(n_658),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_659),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_640),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_661),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_667),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_721),
.A2(n_640),
.B1(n_701),
.B2(n_716),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_713),
.B(n_459),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_668),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_715),
.B(n_1),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_671),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_666),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_674),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_675),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_676),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_717),
.B(n_460),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_677),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_679),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_680),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_681),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_683),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_685),
.Y(n_806)
);

BUFx8_ASAP7_75t_SL g807 ( 
.A(n_702),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_687),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_690),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_767),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_779),
.B(n_708),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_770),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_750),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_744),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_750),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_759),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_724),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_729),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_724),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_787),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_759),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_764),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_774),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_778),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_729),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_730),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_762),
.B(n_708),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_780),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_764),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_752),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_753),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_761),
.B(n_785),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_773),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_755),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_763),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_766),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_787),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_733),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_725),
.B(n_718),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_751),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_751),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_736),
.B(n_719),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_732),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_790),
.Y(n_844)
);

OA21x2_ASAP7_75t_L g845 ( 
.A1(n_756),
.A2(n_693),
.B(n_692),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_775),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_741),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_790),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_796),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_761),
.B(n_720),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_747),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_772),
.A2(n_723),
.B1(n_722),
.B2(n_696),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_744),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_732),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_785),
.B(n_694),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_735),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_749),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_738),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_735),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_739),
.B(n_700),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_737),
.Y(n_861)
);

INVx6_ASAP7_75t_L g862 ( 
.A(n_789),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_775),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_801),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_738),
.Y(n_865)
);

AND2x6_ASAP7_75t_L g866 ( 
.A(n_800),
.B(n_703),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_792),
.B(n_704),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_743),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_734),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_743),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_801),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_745),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_808),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_808),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_809),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_745),
.Y(n_876)
);

INVx6_ASAP7_75t_L g877 ( 
.A(n_795),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_809),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_748),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_795),
.Y(n_880)
);

BUFx8_ASAP7_75t_L g881 ( 
.A(n_796),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_788),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_781),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_737),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_797),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_798),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_788),
.B(n_670),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_799),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_784),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_760),
.B(n_705),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_754),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_799),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_793),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_805),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_802),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_771),
.B(n_672),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_802),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_765),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_803),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_804),
.Y(n_900)
);

AND2x6_ASAP7_75t_L g901 ( 
.A(n_800),
.B(n_706),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_804),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_840),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_814),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_830),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_841),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_825),
.B(n_786),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_835),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_826),
.B(n_678),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_853),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_849),
.B(n_688),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_833),
.B(n_691),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_818),
.B(n_714),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_881),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_882),
.B(n_742),
.Y(n_915)
);

BUFx4f_ASAP7_75t_L g916 ( 
.A(n_862),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_846),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_863),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_864),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_855),
.B(n_832),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_871),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_862),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_836),
.Y(n_923)
);

BUFx8_ASAP7_75t_SL g924 ( 
.A(n_869),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_843),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_883),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_873),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_887),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_874),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_855),
.B(n_777),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_877),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_875),
.Y(n_932)
);

INVx5_ASAP7_75t_L g933 ( 
.A(n_866),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_881),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_878),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_867),
.B(n_746),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_832),
.B(n_771),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_839),
.B(n_769),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_866),
.A2(n_791),
.B1(n_776),
.B2(n_782),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_877),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_880),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_852),
.B(n_757),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_885),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_SL g944 ( 
.A(n_866),
.B(n_807),
.Y(n_944)
);

NAND2xp33_ASAP7_75t_L g945 ( 
.A(n_866),
.B(n_794),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_889),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_811),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_885),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_893),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_842),
.B(n_806),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_827),
.B(n_728),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_896),
.B(n_726),
.Y(n_952)
);

INVx3_ASAP7_75t_R g953 ( 
.A(n_850),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_813),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_811),
.B(n_728),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_886),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_890),
.B(n_760),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_894),
.Y(n_958)
);

INVx4_ASAP7_75t_SL g959 ( 
.A(n_901),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_880),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_860),
.B(n_806),
.Y(n_961)
);

OR2x6_ASAP7_75t_L g962 ( 
.A(n_890),
.B(n_758),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_813),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_880),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_810),
.B(n_782),
.Y(n_965)
);

BUFx10_ASAP7_75t_L g966 ( 
.A(n_850),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_L g967 ( 
.A(n_901),
.B(n_463),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_895),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_831),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_895),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_886),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_813),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_820),
.B(n_783),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_895),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_902),
.Y(n_975)
);

NAND2xp33_ASAP7_75t_SL g976 ( 
.A(n_899),
.B(n_783),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_902),
.B(n_709),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_899),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_821),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_902),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_820),
.B(n_837),
.Y(n_981)
);

INVxp67_ASAP7_75t_SL g982 ( 
.A(n_817),
.Y(n_982)
);

BUFx10_ASAP7_75t_L g983 ( 
.A(n_901),
.Y(n_983)
);

INVxp67_ASAP7_75t_SL g984 ( 
.A(n_817),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_837),
.B(n_710),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_879),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_844),
.B(n_727),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_821),
.Y(n_988)
);

OR2x6_ASAP7_75t_L g989 ( 
.A(n_844),
.B(n_768),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_848),
.B(n_727),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_834),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_821),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_848),
.B(n_768),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_891),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_858),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_888),
.B(n_464),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_888),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_843),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_898),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_892),
.B(n_901),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_843),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_905),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_916),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_983),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_943),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_933),
.B(n_892),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_911),
.B(n_900),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_907),
.B(n_897),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_936),
.B(n_824),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_951),
.B(n_828),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_915),
.B(n_913),
.Y(n_1011)
);

INVxp33_ASAP7_75t_L g1012 ( 
.A(n_909),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_938),
.A2(n_823),
.B1(n_812),
.B2(n_819),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_948),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_947),
.B(n_815),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_966),
.Y(n_1016)
);

OR2x6_ASAP7_75t_L g1017 ( 
.A(n_989),
.B(n_816),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_908),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_955),
.B(n_822),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_956),
.B(n_829),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_971),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_978),
.B(n_819),
.Y(n_1022)
);

AND2x4_ASAP7_75t_SL g1023 ( 
.A(n_966),
.B(n_854),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_933),
.B(n_854),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_986),
.Y(n_1025)
);

AND2x6_ASAP7_75t_L g1026 ( 
.A(n_1000),
.B(n_861),
.Y(n_1026)
);

NAND2xp33_ASAP7_75t_L g1027 ( 
.A(n_933),
.B(n_865),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_942),
.B(n_861),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_994),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_983),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_939),
.B(n_854),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_999),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_959),
.B(n_856),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_904),
.Y(n_1034)
);

NOR3xp33_ASAP7_75t_L g1035 ( 
.A(n_928),
.B(n_870),
.C(n_868),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_912),
.B(n_872),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_920),
.B(n_876),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_923),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_903),
.B(n_884),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_952),
.B(n_838),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_982),
.A2(n_884),
.B(n_845),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_960),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_924),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_906),
.B(n_847),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_937),
.B(n_851),
.Y(n_1045)
);

NOR3xp33_ASAP7_75t_L g1046 ( 
.A(n_922),
.B(n_467),
.C(n_466),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_945),
.A2(n_857),
.B1(n_859),
.B2(n_856),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_959),
.B(n_856),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_960),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_926),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_953),
.B(n_930),
.Y(n_1051)
);

OR2x2_ASAP7_75t_SL g1052 ( 
.A(n_957),
.B(n_944),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_946),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_960),
.B(n_859),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_917),
.Y(n_1055)
);

NOR2xp67_ASAP7_75t_L g1056 ( 
.A(n_941),
.B(n_859),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_918),
.B(n_845),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_919),
.B(n_921),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_962),
.B(n_1),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_927),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_929),
.B(n_469),
.Y(n_1061)
);

INVxp67_ASAP7_75t_SL g1062 ( 
.A(n_984),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_932),
.B(n_470),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_935),
.B(n_471),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_976),
.A2(n_477),
.B1(n_478),
.B2(n_472),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_965),
.A2(n_482),
.B1(n_484),
.B2(n_480),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_949),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_958),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_985),
.B(n_950),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_910),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_985),
.B(n_485),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_993),
.B(n_2),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_967),
.A2(n_498),
.B1(n_505),
.B2(n_487),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_964),
.B(n_506),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_981),
.B(n_512),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_962),
.B(n_3),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_996),
.A2(n_514),
.B1(n_516),
.B2(n_515),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_961),
.B(n_997),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_969),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1011),
.B(n_972),
.Y(n_1080)
);

OR2x6_ASAP7_75t_L g1081 ( 
.A(n_1017),
.B(n_989),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1025),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1029),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_1012),
.B(n_931),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1032),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_1007),
.B(n_979),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1055),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_1008),
.B(n_1001),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_1003),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_1052),
.B(n_940),
.Y(n_1090)
);

AND2x6_ASAP7_75t_L g1091 ( 
.A(n_1004),
.B(n_1030),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1076),
.B(n_934),
.Y(n_1092)
);

AND2x2_ASAP7_75t_SL g1093 ( 
.A(n_1027),
.B(n_1059),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_1023),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_1016),
.B(n_964),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1009),
.B(n_973),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1079),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_1043),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1010),
.B(n_1058),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_1034),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1002),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_1070),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_1069),
.B(n_991),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1060),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1062),
.B(n_975),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1049),
.B(n_964),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_SL g1107 ( 
.A(n_1074),
.B(n_1063),
.C(n_1061),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1018),
.A2(n_995),
.B1(n_963),
.B2(n_988),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_1017),
.B(n_1004),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_SL g1110 ( 
.A1(n_1072),
.A2(n_914),
.B1(n_992),
.B2(n_954),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1038),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_1049),
.B(n_970),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_1036),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_1019),
.B(n_941),
.Y(n_1114)
);

BUFx2_ASAP7_75t_SL g1115 ( 
.A(n_1056),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_1049),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1057),
.A2(n_977),
.B(n_925),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1040),
.B(n_968),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1005),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1014),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_1051),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1064),
.A2(n_925),
.B(n_998),
.C(n_990),
.Y(n_1122)
);

NAND2xp33_ASAP7_75t_L g1123 ( 
.A(n_1021),
.B(n_970),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_1042),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1042),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1050),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_1035),
.B(n_970),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1044),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_1015),
.Y(n_1129)
);

BUFx8_ASAP7_75t_L g1130 ( 
.A(n_1026),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1013),
.B(n_968),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1053),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_1067),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1020),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_1068),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1030),
.B(n_974),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1078),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1026),
.Y(n_1138)
);

XOR2x2_ASAP7_75t_L g1139 ( 
.A(n_1046),
.B(n_987),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1037),
.B(n_974),
.Y(n_1140)
);

O2A1O1Ixp5_ASAP7_75t_L g1141 ( 
.A1(n_1031),
.A2(n_1054),
.B(n_1075),
.C(n_1066),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1026),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1045),
.B(n_980),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1039),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1022),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_1026),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1071),
.B(n_980),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1077),
.B(n_980),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1109),
.B(n_1033),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1086),
.B(n_987),
.Y(n_1150)
);

AND3x1_ASAP7_75t_SL g1151 ( 
.A(n_1119),
.B(n_4),
.C(n_5),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1080),
.B(n_1065),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1099),
.B(n_990),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1113),
.B(n_4),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_1146),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1082),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1138),
.Y(n_1157)
);

NOR2x1p5_ASAP7_75t_L g1158 ( 
.A(n_1098),
.B(n_1028),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1137),
.B(n_1047),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1083),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1109),
.B(n_1048),
.Y(n_1161)
);

OR2x2_ASAP7_75t_SL g1162 ( 
.A(n_1090),
.B(n_493),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1145),
.A2(n_1096),
.B1(n_1118),
.B2(n_1107),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1102),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1085),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1088),
.B(n_1073),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1097),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1087),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1104),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1101),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1111),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1146),
.B(n_1006),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1146),
.B(n_1024),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1129),
.B(n_1041),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1120),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1093),
.B(n_521),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1084),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1138),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1126),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1128),
.B(n_5),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1138),
.B(n_727),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1132),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1081),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1133),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1125),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_1081),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1144),
.B(n_6),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1125),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1130),
.Y(n_1189)
);

NOR2x1p5_ASAP7_75t_L g1190 ( 
.A(n_1094),
.B(n_524),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1134),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1135),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1121),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1135),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1092),
.B(n_7),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1103),
.B(n_8),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1130),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1125),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1141),
.A2(n_531),
.B(n_533),
.C(n_528),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1110),
.A2(n_537),
.B1(n_538),
.B2(n_534),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1114),
.B(n_8),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1139),
.A2(n_1142),
.B1(n_1123),
.B2(n_1140),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1105),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1100),
.B(n_9),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_1089),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1124),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1143),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1095),
.B(n_549),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1116),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_1115),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1108),
.B(n_9),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1136),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1147),
.Y(n_1213)
);

OAI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1196),
.A2(n_1142),
.B1(n_1131),
.B2(n_1148),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_SL g1215 ( 
.A1(n_1201),
.A2(n_1122),
.B(n_1117),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1199),
.A2(n_1163),
.B(n_1174),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1153),
.B(n_1091),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1156),
.B(n_1127),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1213),
.A2(n_1112),
.B(n_1106),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1207),
.A2(n_1091),
.A3(n_1136),
.B(n_62),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1191),
.A2(n_1091),
.B(n_66),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1160),
.A2(n_70),
.B(n_58),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1152),
.B(n_10),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1170),
.A2(n_72),
.A3(n_73),
.B(n_71),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1165),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1164),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1193),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1168),
.A2(n_1175),
.B(n_1169),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1176),
.A2(n_740),
.B(n_731),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1203),
.B(n_10),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1167),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1166),
.A2(n_552),
.B(n_550),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1150),
.B(n_11),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1202),
.A2(n_555),
.B1(n_558),
.B2(n_553),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1177),
.B(n_11),
.Y(n_1235)
);

AOI211x1_ASAP7_75t_L g1236 ( 
.A1(n_1180),
.A2(n_14),
.B(n_12),
.C(n_13),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1198),
.A2(n_75),
.B(n_74),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1171),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1159),
.A2(n_561),
.B(n_559),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_1210),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1179),
.Y(n_1241)
);

OR2x6_ASAP7_75t_L g1242 ( 
.A(n_1189),
.B(n_77),
.Y(n_1242)
);

OAI22x1_ASAP7_75t_L g1243 ( 
.A1(n_1158),
.A2(n_565),
.B1(n_567),
.B2(n_564),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1211),
.A2(n_1187),
.B(n_1208),
.C(n_1200),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1155),
.A2(n_570),
.B(n_568),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1172),
.A2(n_573),
.B(n_574),
.C(n_571),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1204),
.A2(n_577),
.B(n_576),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1205),
.Y(n_1248)
);

NOR4xp25_ASAP7_75t_L g1249 ( 
.A(n_1154),
.B(n_15),
.C(n_13),
.D(n_14),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1206),
.B(n_1195),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1212),
.B(n_16),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1185),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1149),
.B(n_16),
.Y(n_1253)
);

AOI221x1_ASAP7_75t_L g1254 ( 
.A1(n_1184),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.C(n_22),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1189),
.A2(n_1197),
.B(n_1182),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1197),
.A2(n_79),
.B(n_78),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1209),
.B(n_20),
.Y(n_1257)
);

INVx5_ASAP7_75t_L g1258 ( 
.A(n_1157),
.Y(n_1258)
);

NAND2x1_ASAP7_75t_L g1259 ( 
.A(n_1155),
.B(n_80),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1185),
.B(n_579),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1173),
.A2(n_590),
.B(n_584),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1192),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1194),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1190),
.A2(n_83),
.B(n_82),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1149),
.B(n_21),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1162),
.A2(n_603),
.B1(n_607),
.B2(n_596),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1172),
.A2(n_1161),
.B(n_1173),
.C(n_1151),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1161),
.A2(n_610),
.B(n_609),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1188),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1181),
.A2(n_612),
.B(n_611),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1185),
.A2(n_616),
.B(n_614),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1157),
.A2(n_620),
.B(n_619),
.C(n_731),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1157),
.A2(n_85),
.A3(n_87),
.B(n_84),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1186),
.B(n_23),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1183),
.B(n_23),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1188),
.Y(n_1276)
);

INVxp67_ASAP7_75t_SL g1277 ( 
.A(n_1188),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1178),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1178),
.A2(n_90),
.B(n_89),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1178),
.A2(n_1181),
.B(n_95),
.Y(n_1280)
);

OAI222xp33_ASAP7_75t_L g1281 ( 
.A1(n_1211),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.C1(n_27),
.C2(n_28),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1152),
.A2(n_740),
.B1(n_731),
.B2(n_29),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1177),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1177),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1167),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1153),
.B(n_26),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1174),
.A2(n_96),
.B(n_91),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1153),
.B(n_28),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1152),
.B(n_29),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1199),
.A2(n_98),
.A3(n_99),
.B(n_97),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1152),
.B(n_30),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1199),
.A2(n_740),
.B(n_30),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1199),
.A2(n_31),
.B(n_33),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1156),
.Y(n_1294)
);

OAI21xp33_ASAP7_75t_L g1295 ( 
.A1(n_1201),
.A2(n_31),
.B(n_33),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1283),
.B(n_34),
.Y(n_1296)
);

CKINVDCx9p33_ASAP7_75t_R g1297 ( 
.A(n_1223),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1225),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1294),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1284),
.B(n_34),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1289),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1228),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1231),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1291),
.B(n_35),
.Y(n_1304)
);

CKINVDCx16_ASAP7_75t_R g1305 ( 
.A(n_1226),
.Y(n_1305)
);

CKINVDCx8_ASAP7_75t_R g1306 ( 
.A(n_1227),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1248),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1216),
.A2(n_36),
.B(n_38),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1221),
.A2(n_101),
.B(n_100),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1258),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1250),
.B(n_38),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_SL g1312 ( 
.A(n_1240),
.B(n_1267),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1258),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1242),
.B(n_102),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1269),
.B(n_40),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1252),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1218),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1215),
.A2(n_1217),
.B(n_1214),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1285),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1238),
.Y(n_1320)
);

OR2x6_ASAP7_75t_SL g1321 ( 
.A(n_1235),
.B(n_41),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1276),
.Y(n_1322)
);

CKINVDCx11_ASAP7_75t_R g1323 ( 
.A(n_1242),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1258),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1277),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1278),
.B(n_103),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1241),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1282),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1255),
.B(n_105),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1262),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1263),
.Y(n_1331)
);

O2A1O1Ixp5_ASAP7_75t_SL g1332 ( 
.A1(n_1230),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1233),
.B(n_45),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1275),
.Y(n_1334)
);

INVx5_ASAP7_75t_L g1335 ( 
.A(n_1243),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1292),
.A2(n_46),
.B(n_47),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1293),
.A2(n_1295),
.B(n_1244),
.Y(n_1337)
);

NOR2xp67_ASAP7_75t_SL g1338 ( 
.A(n_1268),
.B(n_47),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1257),
.B(n_48),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1274),
.Y(n_1340)
);

CKINVDCx6p67_ASAP7_75t_R g1341 ( 
.A(n_1253),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1286),
.B(n_48),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1219),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1288),
.B(n_49),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1249),
.B(n_50),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1265),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1236),
.B(n_50),
.Y(n_1347)
);

AND2x2_ASAP7_75t_SL g1348 ( 
.A(n_1251),
.B(n_51),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1220),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1261),
.B(n_52),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1232),
.A2(n_1259),
.B(n_1247),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1264),
.B(n_106),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1220),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1280),
.B(n_107),
.Y(n_1354)
);

INVx5_ASAP7_75t_L g1355 ( 
.A(n_1281),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1234),
.B(n_1270),
.Y(n_1356)
);

BUFx12f_ASAP7_75t_L g1357 ( 
.A(n_1260),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1287),
.A2(n_52),
.B(n_53),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1273),
.B(n_108),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1256),
.A2(n_53),
.B(n_54),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1224),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1290),
.Y(n_1362)
);

INVx5_ASAP7_75t_L g1363 ( 
.A(n_1273),
.Y(n_1363)
);

O2A1O1Ixp5_ASAP7_75t_SL g1364 ( 
.A1(n_1266),
.A2(n_56),
.B(n_57),
.C(n_113),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_1271),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1254),
.B(n_56),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1222),
.A2(n_57),
.B(n_114),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1224),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1229),
.B(n_115),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1290),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1246),
.B(n_118),
.Y(n_1371)
);

A2O1A1Ixp33_ASAP7_75t_SL g1372 ( 
.A1(n_1239),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1272),
.B(n_123),
.Y(n_1373)
);

OR2x6_ASAP7_75t_L g1374 ( 
.A(n_1279),
.B(n_124),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1317),
.B(n_1237),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1337),
.A2(n_1245),
.B(n_125),
.Y(n_1376)
);

OA22x2_ASAP7_75t_L g1377 ( 
.A1(n_1314),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1306),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1322),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1325),
.B(n_129),
.Y(n_1380)
);

NOR2xp67_ASAP7_75t_L g1381 ( 
.A(n_1335),
.B(n_131),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1298),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1305),
.B(n_447),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1351),
.A2(n_132),
.B(n_133),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1341),
.B(n_134),
.Y(n_1385)
);

AND2x2_ASAP7_75t_SL g1386 ( 
.A(n_1312),
.B(n_135),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1318),
.B(n_137),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1299),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1308),
.A2(n_138),
.B(n_139),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1330),
.B(n_140),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1331),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1303),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1316),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1346),
.B(n_141),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1320),
.B(n_143),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1313),
.B(n_144),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1314),
.A2(n_145),
.B(n_148),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1304),
.A2(n_153),
.B(n_149),
.C(n_151),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1296),
.B(n_154),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1307),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_SL g1401 ( 
.A1(n_1344),
.A2(n_161),
.B(n_156),
.C(n_158),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1356),
.A2(n_166),
.B1(n_163),
.B2(n_164),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1319),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1302),
.B(n_169),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1327),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1370),
.A2(n_171),
.B(n_173),
.Y(n_1406)
);

INVxp67_ASAP7_75t_SL g1407 ( 
.A(n_1343),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1311),
.B(n_175),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1334),
.B(n_445),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1300),
.B(n_177),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1362),
.A2(n_178),
.B(n_179),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1349),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1333),
.B(n_180),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1339),
.B(n_181),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1342),
.B(n_183),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1353),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1348),
.B(n_185),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1340),
.B(n_444),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1323),
.B(n_187),
.Y(n_1419)
);

O2A1O1Ixp5_ASAP7_75t_L g1420 ( 
.A1(n_1345),
.A2(n_191),
.B(n_189),
.C(n_190),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1315),
.B(n_192),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1310),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1361),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1368),
.Y(n_1424)
);

BUFx5_ASAP7_75t_L g1425 ( 
.A(n_1359),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1310),
.B(n_193),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1347),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1363),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1363),
.Y(n_1429)
);

O2A1O1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1301),
.A2(n_195),
.B(n_200),
.C(n_201),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1357),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1355),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1324),
.B(n_206),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1366),
.B(n_207),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1321),
.B(n_208),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1350),
.B(n_443),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1324),
.B(n_209),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1326),
.B(n_210),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1329),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1328),
.A2(n_213),
.B(n_214),
.C(n_215),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1297),
.A2(n_442),
.B1(n_218),
.B2(n_219),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1369),
.A2(n_216),
.B(n_220),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1335),
.Y(n_1443)
);

OR2x6_ASAP7_75t_SL g1444 ( 
.A(n_1371),
.B(n_221),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1367),
.A2(n_222),
.B(n_223),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_SL g1446 ( 
.A(n_1355),
.B(n_224),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1365),
.Y(n_1447)
);

NOR2xp67_ASAP7_75t_L g1448 ( 
.A(n_1360),
.B(n_226),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1354),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1352),
.B(n_441),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1338),
.B(n_227),
.Y(n_1451)
);

AOI21x1_ASAP7_75t_SL g1452 ( 
.A1(n_1373),
.A2(n_228),
.B(n_229),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1374),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1382),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1388),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1447),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1391),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1379),
.B(n_1374),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1392),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1416),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_1375),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1403),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1411),
.A2(n_1358),
.B(n_1332),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1453),
.B(n_1309),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1386),
.A2(n_1446),
.B1(n_1427),
.B2(n_1377),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1443),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1412),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1422),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1405),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1439),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1407),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1411),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1423),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1424),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1422),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1449),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1428),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1429),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1425),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1425),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1400),
.B(n_1336),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1425),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1425),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1395),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1395),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1378),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1404),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1397),
.B(n_1380),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1452),
.A2(n_1384),
.B(n_1420),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1404),
.Y(n_1490)
);

OA21x2_ASAP7_75t_L g1491 ( 
.A1(n_1409),
.A2(n_1364),
.B(n_1372),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1434),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1394),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1396),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1390),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1413),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1393),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1444),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1432),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1387),
.A2(n_234),
.B(n_235),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1431),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1435),
.B(n_236),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1415),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1396),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1383),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1406),
.A2(n_238),
.B(n_239),
.Y(n_1506)
);

AO21x2_ASAP7_75t_L g1507 ( 
.A1(n_1448),
.A2(n_240),
.B(n_241),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1385),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1471),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1460),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1488),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1456),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1456),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1454),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1461),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1461),
.B(n_1418),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1492),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1467),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1465),
.A2(n_1441),
.B1(n_1414),
.B2(n_1436),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1455),
.Y(n_1520)
);

AO31x2_ASAP7_75t_L g1521 ( 
.A1(n_1477),
.A2(n_1493),
.A3(n_1473),
.B(n_1474),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1458),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1498),
.B(n_1417),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1458),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1476),
.B(n_1419),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1457),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1470),
.B(n_1408),
.Y(n_1527)
);

AOI221xp5_ASAP7_75t_L g1528 ( 
.A1(n_1472),
.A2(n_1410),
.B1(n_1398),
.B2(n_1430),
.C(n_1399),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1476),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1459),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1462),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1478),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1492),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1466),
.B(n_1421),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1469),
.Y(n_1535)
);

BUFx12f_ASAP7_75t_L g1536 ( 
.A(n_1501),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1496),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1466),
.B(n_1450),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1503),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1505),
.B(n_1437),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1488),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1472),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1505),
.B(n_1451),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1464),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1497),
.B(n_1426),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1464),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1488),
.A2(n_1376),
.B1(n_1440),
.B2(n_1389),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1479),
.B(n_1401),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_1486),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1480),
.B(n_1426),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1468),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1482),
.B(n_1438),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1468),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1517),
.B(n_1487),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1522),
.B(n_1475),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1533),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1517),
.B(n_1490),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1522),
.B(n_1475),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1521),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1523),
.B(n_1502),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1512),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1524),
.B(n_1483),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1536),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1513),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1511),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1521),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1524),
.B(n_1525),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1551),
.B(n_1508),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1511),
.B(n_1541),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1553),
.B(n_1484),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1510),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1514),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1542),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1548),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1529),
.B(n_1485),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1529),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1542),
.B(n_1481),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1519),
.A2(n_1491),
.B1(n_1463),
.B2(n_1502),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1543),
.B(n_1494),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1532),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1532),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1521),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1521),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1577),
.B(n_1539),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1571),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1567),
.B(n_1534),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1554),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1577),
.B(n_1515),
.Y(n_1588)
);

INVxp67_ASAP7_75t_SL g1589 ( 
.A(n_1574),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1556),
.B(n_1511),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1574),
.B(n_1531),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1565),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1561),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1572),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1573),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1580),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1573),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1565),
.Y(n_1598)
);

BUFx2_ASAP7_75t_SL g1599 ( 
.A(n_1563),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1557),
.B(n_1564),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1578),
.B(n_1520),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1555),
.B(n_1538),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1580),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1557),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1565),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1563),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1578),
.B(n_1581),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1581),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1568),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1589),
.B(n_1560),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1586),
.B(n_1558),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1602),
.B(n_1549),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1593),
.Y(n_1613)
);

NAND4xp25_ASAP7_75t_L g1614 ( 
.A(n_1606),
.B(n_1519),
.C(n_1523),
.D(n_1528),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1592),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1609),
.B(n_1562),
.Y(n_1616)
);

NAND4xp25_ASAP7_75t_L g1617 ( 
.A(n_1607),
.B(n_1528),
.C(n_1548),
.D(n_1560),
.Y(n_1617)
);

INVx4_ASAP7_75t_L g1618 ( 
.A(n_1599),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1585),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1584),
.B(n_1527),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1607),
.A2(n_1601),
.B1(n_1547),
.B2(n_1587),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1598),
.Y(n_1622)
);

AO21x2_ASAP7_75t_L g1623 ( 
.A1(n_1601),
.A2(n_1566),
.B(n_1559),
.Y(n_1623)
);

OAI222xp33_ASAP7_75t_SL g1624 ( 
.A1(n_1591),
.A2(n_1541),
.B1(n_1511),
.B2(n_1565),
.C1(n_1530),
.C2(n_1526),
.Y(n_1624)
);

OAI33xp33_ASAP7_75t_L g1625 ( 
.A1(n_1596),
.A2(n_1516),
.A3(n_1547),
.B1(n_1515),
.B2(n_1509),
.B3(n_1535),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1610),
.B(n_1591),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1619),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1611),
.B(n_1605),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1615),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1619),
.Y(n_1630)
);

NAND2x1_ASAP7_75t_L g1631 ( 
.A(n_1612),
.B(n_1576),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1612),
.B(n_1604),
.Y(n_1632)
);

AND2x4_ASAP7_75t_SL g1633 ( 
.A(n_1618),
.B(n_1545),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1613),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1620),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1622),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1635),
.B(n_1617),
.Y(n_1637)
);

NOR2x1_ASAP7_75t_L g1638 ( 
.A(n_1631),
.B(n_1618),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1626),
.B(n_1614),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1629),
.B(n_1621),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1628),
.B(n_1616),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1627),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1632),
.B(n_1594),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1636),
.B(n_1595),
.Y(n_1644)
);

AND2x2_ASAP7_75t_SL g1645 ( 
.A(n_1633),
.B(n_1541),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1636),
.B(n_1595),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1630),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1634),
.Y(n_1648)
);

NOR2x1p5_ASAP7_75t_L g1649 ( 
.A(n_1637),
.B(n_1603),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1643),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1644),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1641),
.B(n_1600),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1646),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1645),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1648),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1638),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1648),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1642),
.B(n_1597),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1639),
.B(n_1597),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1659),
.B(n_1647),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1652),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1650),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1658),
.B(n_1640),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1656),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1649),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1655),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1657),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1651),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1649),
.B(n_1608),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1654),
.B(n_1590),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1662),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1663),
.A2(n_1625),
.B1(n_1653),
.B2(n_1623),
.Y(n_1672)
);

AOI32xp33_ASAP7_75t_L g1673 ( 
.A1(n_1665),
.A2(n_1590),
.A3(n_1624),
.B1(n_1588),
.B2(n_1489),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1661),
.A2(n_1541),
.B(n_1569),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1660),
.Y(n_1675)
);

NAND4xp25_ASAP7_75t_L g1676 ( 
.A(n_1664),
.B(n_1381),
.C(n_1500),
.D(n_1569),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1665),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_SL g1678 ( 
.A(n_1668),
.B(n_1500),
.C(n_1499),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1670),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_SL g1680 ( 
.A1(n_1666),
.A2(n_1509),
.B(n_1402),
.C(n_1546),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1679),
.B(n_1669),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1674),
.B(n_1667),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1675),
.B(n_1579),
.Y(n_1683)
);

CKINVDCx16_ASAP7_75t_R g1684 ( 
.A(n_1671),
.Y(n_1684)
);

AOI21xp33_ASAP7_75t_L g1685 ( 
.A1(n_1677),
.A2(n_1583),
.B(n_1582),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1672),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1678),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_SL g1688 ( 
.A1(n_1673),
.A2(n_1552),
.B(n_1570),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1680),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1676),
.B(n_1575),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1679),
.B(n_1540),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1675),
.Y(n_1692)
);

OAI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1672),
.A2(n_1546),
.B1(n_1504),
.B2(n_1494),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1679),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1681),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1684),
.B(n_1494),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1694),
.B(n_1550),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1691),
.B(n_1692),
.Y(n_1698)
);

NAND2xp33_ASAP7_75t_L g1699 ( 
.A(n_1689),
.B(n_1504),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1683),
.B(n_1518),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1687),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1682),
.B(n_1504),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1693),
.A2(n_1445),
.B(n_1442),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1690),
.B(n_1544),
.Y(n_1704)
);

INVxp67_ASAP7_75t_L g1705 ( 
.A(n_1686),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1685),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1698),
.B(n_1688),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1701),
.Y(n_1708)
);

NOR2x1_ASAP7_75t_L g1709 ( 
.A(n_1695),
.B(n_1433),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1697),
.B(n_1518),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_L g1711 ( 
.A(n_1699),
.B(n_1491),
.C(n_1537),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1696),
.B(n_1507),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1700),
.Y(n_1713)
);

NAND3xp33_ASAP7_75t_L g1714 ( 
.A(n_1705),
.B(n_1495),
.C(n_1506),
.Y(n_1714)
);

AOI222xp33_ASAP7_75t_L g1715 ( 
.A1(n_1706),
.A2(n_1507),
.B1(n_244),
.B2(n_247),
.C1(n_248),
.C2(n_249),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1708),
.A2(n_1707),
.B(n_1702),
.Y(n_1716)
);

OAI211xp5_ASAP7_75t_L g1717 ( 
.A1(n_1713),
.A2(n_1704),
.B(n_1703),
.C(n_252),
.Y(n_1717)
);

AOI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1711),
.A2(n_242),
.B(n_250),
.C(n_253),
.Y(n_1718)
);

O2A1O1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1712),
.A2(n_254),
.B(n_255),
.C(n_256),
.Y(n_1719)
);

OAI22xp33_ASAP7_75t_SL g1720 ( 
.A1(n_1709),
.A2(n_257),
.B1(n_259),
.B2(n_262),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1715),
.B(n_263),
.Y(n_1721)
);

NAND3xp33_ASAP7_75t_L g1722 ( 
.A(n_1714),
.B(n_265),
.C(n_266),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1710),
.A2(n_268),
.B(n_269),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1713),
.B(n_274),
.Y(n_1724)
);

NAND5xp2_ASAP7_75t_L g1725 ( 
.A(n_1707),
.B(n_275),
.C(n_276),
.D(n_278),
.E(n_282),
.Y(n_1725)
);

OAI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1708),
.A2(n_283),
.B1(n_285),
.B2(n_287),
.C(n_288),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1708),
.A2(n_290),
.B1(n_292),
.B2(n_296),
.Y(n_1727)
);

NOR2x1_ASAP7_75t_L g1728 ( 
.A(n_1708),
.B(n_297),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1724),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1728),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1716),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1717),
.Y(n_1732)
);

AOI211xp5_ASAP7_75t_L g1733 ( 
.A1(n_1720),
.A2(n_298),
.B(n_301),
.C(n_302),
.Y(n_1733)
);

OAI32xp33_ASAP7_75t_L g1734 ( 
.A1(n_1722),
.A2(n_303),
.A3(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1721),
.A2(n_310),
.B1(n_312),
.B2(n_313),
.Y(n_1735)
);

NAND4xp25_ASAP7_75t_L g1736 ( 
.A(n_1718),
.B(n_314),
.C(n_315),
.D(n_316),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1725),
.B(n_317),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1723),
.B(n_318),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1719),
.Y(n_1739)
);

OAI21xp33_ASAP7_75t_L g1740 ( 
.A1(n_1726),
.A2(n_320),
.B(n_321),
.Y(n_1740)
);

O2A1O1Ixp33_ASAP7_75t_L g1741 ( 
.A1(n_1727),
.A2(n_322),
.B(n_326),
.C(n_327),
.Y(n_1741)
);

NAND3xp33_ASAP7_75t_L g1742 ( 
.A(n_1728),
.B(n_328),
.C(n_329),
.Y(n_1742)
);

AOI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1722),
.A2(n_331),
.B1(n_334),
.B2(n_335),
.C(n_336),
.Y(n_1743)
);

NOR3xp33_ASAP7_75t_L g1744 ( 
.A(n_1731),
.B(n_337),
.C(n_338),
.Y(n_1744)
);

NOR3xp33_ASAP7_75t_L g1745 ( 
.A(n_1729),
.B(n_339),
.C(n_340),
.Y(n_1745)
);

NAND3xp33_ASAP7_75t_L g1746 ( 
.A(n_1730),
.B(n_342),
.C(n_344),
.Y(n_1746)
);

OAI21xp33_ASAP7_75t_L g1747 ( 
.A1(n_1732),
.A2(n_346),
.B(n_347),
.Y(n_1747)
);

NOR2x1_ASAP7_75t_L g1748 ( 
.A(n_1742),
.B(n_348),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1737),
.Y(n_1749)
);

NAND4xp75_ASAP7_75t_L g1750 ( 
.A(n_1739),
.B(n_349),
.C(n_350),
.D(n_351),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1738),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1735),
.B(n_352),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1743),
.B(n_356),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1740),
.B(n_358),
.Y(n_1754)
);

NOR2x1_ASAP7_75t_L g1755 ( 
.A(n_1736),
.B(n_359),
.Y(n_1755)
);

NAND4xp75_ASAP7_75t_L g1756 ( 
.A(n_1733),
.B(n_360),
.C(n_361),
.D(n_362),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1741),
.B(n_363),
.Y(n_1757)
);

NAND3xp33_ASAP7_75t_L g1758 ( 
.A(n_1734),
.B(n_365),
.C(n_366),
.Y(n_1758)
);

NOR2x1_ASAP7_75t_L g1759 ( 
.A(n_1731),
.B(n_367),
.Y(n_1759)
);

OAI211xp5_ASAP7_75t_L g1760 ( 
.A1(n_1731),
.A2(n_369),
.B(n_370),
.C(n_371),
.Y(n_1760)
);

NOR2x1_ASAP7_75t_L g1761 ( 
.A(n_1731),
.B(n_372),
.Y(n_1761)
);

AOI21xp33_ASAP7_75t_SL g1762 ( 
.A1(n_1731),
.A2(n_373),
.B(n_374),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1737),
.Y(n_1763)
);

NOR2x1_ASAP7_75t_L g1764 ( 
.A(n_1749),
.B(n_376),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1763),
.B(n_378),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1751),
.Y(n_1766)
);

XNOR2x1_ASAP7_75t_L g1767 ( 
.A(n_1759),
.B(n_380),
.Y(n_1767)
);

NOR3xp33_ASAP7_75t_L g1768 ( 
.A(n_1761),
.B(n_384),
.C(n_385),
.Y(n_1768)
);

OAI211xp5_ASAP7_75t_SL g1769 ( 
.A1(n_1753),
.A2(n_386),
.B(n_389),
.C(n_390),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1755),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1757),
.B(n_393),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1754),
.B(n_394),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1748),
.Y(n_1773)
);

INVx2_ASAP7_75t_SL g1774 ( 
.A(n_1752),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1770),
.B(n_1762),
.Y(n_1775)
);

XNOR2xp5_ASAP7_75t_L g1776 ( 
.A(n_1767),
.B(n_1756),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1773),
.B(n_1747),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1764),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1765),
.B(n_1774),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1766),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1771),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1772),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1779),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1778),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1781),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1782),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_1783),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1784),
.A2(n_1780),
.B1(n_1775),
.B2(n_1777),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1788),
.A2(n_1785),
.B1(n_1786),
.B2(n_1776),
.Y(n_1789)
);

BUFx6f_ASAP7_75t_L g1790 ( 
.A(n_1787),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_SL g1791 ( 
.A1(n_1790),
.A2(n_1746),
.B1(n_1758),
.B2(n_1768),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1789),
.A2(n_1769),
.B(n_1744),
.Y(n_1792)
);

AOI21xp33_ASAP7_75t_L g1793 ( 
.A1(n_1792),
.A2(n_1791),
.B(n_1760),
.Y(n_1793)
);

NOR3xp33_ASAP7_75t_SL g1794 ( 
.A(n_1792),
.B(n_1750),
.C(n_1745),
.Y(n_1794)
);

NOR2x1_ASAP7_75t_L g1795 ( 
.A(n_1793),
.B(n_1794),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1794),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1795),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1796),
.A2(n_395),
.B1(n_396),
.B2(n_397),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_L g1799 ( 
.A(n_1797),
.B(n_399),
.C(n_400),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_SL g1800 ( 
.A1(n_1798),
.A2(n_402),
.B1(n_407),
.B2(n_408),
.Y(n_1800)
);

OAI21xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1797),
.A2(n_410),
.B(n_411),
.Y(n_1801)
);

NAND3xp33_ASAP7_75t_L g1802 ( 
.A(n_1797),
.B(n_412),
.C(n_414),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1800),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1801),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1799),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1803),
.B(n_1802),
.Y(n_1806)
);

OR2x6_ASAP7_75t_L g1807 ( 
.A(n_1804),
.B(n_1805),
.Y(n_1807)
);

OR2x6_ASAP7_75t_L g1808 ( 
.A(n_1804),
.B(n_415),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1807),
.A2(n_416),
.B(n_418),
.Y(n_1809)
);

AOI211xp5_ASAP7_75t_L g1810 ( 
.A1(n_1809),
.A2(n_1806),
.B(n_1808),
.C(n_425),
.Y(n_1810)
);


endmodule