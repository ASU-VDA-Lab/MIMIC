module fake_netlist_6_3144_n_1925 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1925);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1925;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_873;
wire n_461;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_102),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_54),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_164),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_96),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_81),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_120),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_79),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_44),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_142),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_130),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_155),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_134),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_62),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_100),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_49),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_9),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_27),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_131),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_119),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_34),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_77),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_18),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_68),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_129),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_140),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_82),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_86),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_128),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_50),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_136),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_168),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_87),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_45),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_71),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_135),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_112),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_64),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_196),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_169),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_10),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_111),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_183),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_9),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_32),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_69),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_144),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_181),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_176),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_48),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_182),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_137),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_84),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_159),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_5),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_171),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_72),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_39),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_19),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_114),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_113),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_122),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_174),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_66),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_23),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_150),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_192),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_166),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_51),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_165),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_170),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_21),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_51),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_78),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_123),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_90),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_97),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_158),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_19),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_65),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_58),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_127),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_55),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_110),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_58),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_99),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_12),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_61),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_74),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_24),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_46),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_115),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_40),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_59),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_21),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_188),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_197),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_64),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_46),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_107),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_5),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_7),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_2),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_13),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_14),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_163),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_76),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_57),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_152),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_56),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_13),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_67),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_72),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_186),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_60),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_26),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_6),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_121),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_173),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_67),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_156),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_179),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_194),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_141),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_23),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_91),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_178),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_125),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_55),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_195),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_75),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_109),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_50),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_66),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_7),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_172),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_124),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_34),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_63),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_63),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_153),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_49),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_39),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_69),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_47),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_40),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_185),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_60),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_68),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_28),
.Y(n_351)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_151),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_6),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_24),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_154),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_108),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_3),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_117),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_94),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_145),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_106),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_27),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_139),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_15),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_95),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_143),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_161),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_167),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_31),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_41),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_61),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_88),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_15),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_36),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_104),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_193),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_53),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_18),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_162),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_157),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_4),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_41),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_16),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_80),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_160),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_56),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_126),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_118),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_93),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_146),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_98),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_38),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_52),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_294),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_294),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_202),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_294),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_294),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_294),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_201),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_311),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_204),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_311),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_311),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_311),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_311),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_217),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_217),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_357),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_349),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_357),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_205),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_200),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_318),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_226),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_200),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_206),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_207),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_208),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_207),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_283),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_227),
.Y(n_423)
);

INVxp33_ASAP7_75t_SL g424 ( 
.A(n_347),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_209),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_231),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_210),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_213),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_239),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_218),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_213),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_223),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_223),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_283),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_224),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_228),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_230),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_262),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_377),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_198),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_232),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_243),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_235),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_341),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_370),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_264),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_238),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_283),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_243),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_246),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_242),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_246),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_268),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_266),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_331),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_247),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_283),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_266),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_282),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_356),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_273),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_273),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_274),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_274),
.Y(n_464)
);

INVxp33_ASAP7_75t_SL g465 ( 
.A(n_215),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_214),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_211),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_225),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_289),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_289),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_236),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_198),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_216),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_240),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_292),
.Y(n_475)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_211),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_292),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_306),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_306),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_240),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_313),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_326),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_326),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_283),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_229),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_335),
.Y(n_486)
);

INVxp33_ASAP7_75t_L g487 ( 
.A(n_335),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_220),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_283),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_350),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_350),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_353),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_250),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_353),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_236),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_396),
.B(n_380),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_404),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_404),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_402),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_394),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_459),
.A2(n_346),
.B1(n_362),
.B2(n_354),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_395),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_395),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_397),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_398),
.B(n_221),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_398),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_354),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_445),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_399),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_418),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_485),
.Y(n_514)
);

AO22x1_ASAP7_75t_L g515 ( 
.A1(n_467),
.A2(n_364),
.B1(n_369),
.B2(n_362),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_399),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_401),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_401),
.Y(n_518)
);

INVx6_ASAP7_75t_L g519 ( 
.A(n_471),
.Y(n_519)
);

AND2x2_ASAP7_75t_SL g520 ( 
.A(n_468),
.B(n_221),
.Y(n_520)
);

BUFx10_ASAP7_75t_L g521 ( 
.A(n_420),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_471),
.B(n_364),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_403),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_425),
.B(n_245),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_422),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_466),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_422),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_427),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_430),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_403),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_405),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_465),
.B(n_252),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_476),
.B(n_369),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_434),
.A2(n_261),
.B(n_245),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_487),
.B(n_371),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_405),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_435),
.B(n_320),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_424),
.A2(n_336),
.B1(n_234),
.B2(n_233),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_436),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_406),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_406),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_437),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_434),
.Y(n_543)
);

CKINVDCx6p67_ASAP7_75t_R g544 ( 
.A(n_415),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_448),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_414),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_448),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_457),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_457),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_440),
.B(n_261),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_438),
.B(n_371),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_441),
.B(n_333),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_444),
.B(n_372),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_417),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_484),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_472),
.B(n_333),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_484),
.B(n_363),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_417),
.Y(n_558)
);

INVx6_ASAP7_75t_L g559 ( 
.A(n_474),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_419),
.Y(n_560)
);

NOR2x1_ASAP7_75t_L g561 ( 
.A(n_493),
.B(n_363),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_419),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_421),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_410),
.A2(n_393),
.B1(n_392),
.B2(n_256),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_489),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_421),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_443),
.B(n_376),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_400),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_428),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_413),
.A2(n_383),
.B1(n_258),
.B2(n_259),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_428),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_489),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_407),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_416),
.A2(n_383),
.B1(n_251),
.B2(n_244),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_447),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_431),
.B(n_376),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_431),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_423),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_432),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_527),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_532),
.B(n_451),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_496),
.B(n_456),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_502),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_502),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_547),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_514),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_547),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_537),
.B(n_460),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_504),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_524),
.B(n_473),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_543),
.Y(n_591)
);

AO21x2_ASAP7_75t_L g592 ( 
.A1(n_552),
.A2(n_348),
.B(n_199),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_543),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_544),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_545),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_L g596 ( 
.A(n_567),
.B(n_283),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_545),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_504),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_547),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_547),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_507),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g602 ( 
.A(n_564),
.B(n_488),
.C(n_412),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_507),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_520),
.B(n_480),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_520),
.B(n_439),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_501),
.B(n_253),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_548),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_527),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_497),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_559),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_544),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_501),
.B(n_254),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_519),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_511),
.Y(n_614)
);

BUFx6f_ASAP7_75t_SL g615 ( 
.A(n_521),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_548),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_501),
.B(n_255),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_501),
.B(n_257),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_510),
.B(n_263),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_510),
.B(n_407),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_515),
.B(n_203),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_520),
.B(n_267),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_549),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_512),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_521),
.B(n_276),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_533),
.B(n_277),
.Y(n_626)
);

INVxp33_ASAP7_75t_L g627 ( 
.A(n_511),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_547),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_512),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_518),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_559),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_518),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_541),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_549),
.Y(n_634)
);

NAND2xp33_ASAP7_75t_L g635 ( 
.A(n_561),
.B(n_283),
.Y(n_635)
);

INVxp33_ASAP7_75t_SL g636 ( 
.A(n_570),
.Y(n_636)
);

INVxp33_ASAP7_75t_L g637 ( 
.A(n_535),
.Y(n_637)
);

BUFx10_ASAP7_75t_L g638 ( 
.A(n_559),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_546),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_541),
.Y(n_640)
);

BUFx10_ASAP7_75t_L g641 ( 
.A(n_559),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_561),
.A2(n_429),
.B1(n_446),
.B2(n_426),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_546),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_497),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_554),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_535),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_521),
.B(n_278),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_555),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_521),
.B(n_287),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_553),
.A2(n_455),
.B1(n_453),
.B2(n_297),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_564),
.B(n_237),
.C(n_222),
.Y(n_651)
);

INVxp67_ASAP7_75t_SL g652 ( 
.A(n_547),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_522),
.B(n_408),
.Y(n_653)
);

AOI21x1_ASAP7_75t_L g654 ( 
.A1(n_557),
.A2(n_212),
.B(n_203),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_568),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_578),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_555),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_575),
.A2(n_304),
.B1(n_300),
.B2(n_299),
.Y(n_658)
);

CKINVDCx16_ASAP7_75t_R g659 ( 
.A(n_526),
.Y(n_659)
);

CKINVDCx6p67_ASAP7_75t_R g660 ( 
.A(n_575),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_565),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_497),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_519),
.B(n_260),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_L g664 ( 
.A(n_572),
.B(n_283),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_565),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_499),
.B(n_293),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_L g667 ( 
.A(n_538),
.B(n_270),
.C(n_265),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_557),
.Y(n_668)
);

AO21x2_ASAP7_75t_L g669 ( 
.A1(n_534),
.A2(n_219),
.B(n_212),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_515),
.B(n_219),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_557),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_572),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_573),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_557),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_519),
.B(n_280),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_519),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_522),
.B(n_576),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_572),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_533),
.B(n_298),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_572),
.B(n_301),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_551),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_573),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_554),
.Y(n_683)
);

NAND3xp33_ASAP7_75t_L g684 ( 
.A(n_551),
.B(n_284),
.C(n_281),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_573),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_558),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_573),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_573),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_500),
.Y(n_689)
);

INVx5_ASAP7_75t_L g690 ( 
.A(n_572),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_513),
.B(n_286),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_500),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_505),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_528),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_572),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_529),
.B(n_288),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_497),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_558),
.B(n_408),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_L g699 ( 
.A(n_539),
.B(n_295),
.C(n_291),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_573),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_497),
.B(n_308),
.Y(n_701)
);

CKINVDCx6p67_ASAP7_75t_R g702 ( 
.A(n_526),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_505),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_542),
.A2(n_296),
.B1(n_302),
.B2(n_303),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_509),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_525),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_570),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_497),
.B(n_315),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_525),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_574),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_525),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_525),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_527),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_509),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_516),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_498),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_498),
.B(n_319),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_516),
.Y(n_718)
);

AND3x2_ASAP7_75t_L g719 ( 
.A(n_576),
.B(n_379),
.C(n_248),
.Y(n_719)
);

BUFx4f_ASAP7_75t_L g720 ( 
.A(n_498),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_574),
.B(n_241),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_517),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_560),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_498),
.B(n_324),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_R g725 ( 
.A(n_579),
.B(n_325),
.Y(n_725)
);

XOR2xp5_ASAP7_75t_L g726 ( 
.A(n_503),
.B(n_305),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_498),
.B(n_352),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_668),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_582),
.B(n_508),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_668),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_671),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_681),
.A2(n_503),
.B1(n_550),
.B2(n_556),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_684),
.B(n_312),
.C(n_309),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_681),
.B(n_338),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_671),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_674),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_674),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_588),
.B(n_508),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_698),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_637),
.B(n_314),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_590),
.B(n_316),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_677),
.B(n_338),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_677),
.B(n_550),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_715),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_698),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_638),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_622),
.B(n_338),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_639),
.B(n_556),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_592),
.A2(n_556),
.B1(n_576),
.B2(n_241),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_643),
.B(n_517),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_586),
.B(n_560),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_638),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_715),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_653),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_646),
.B(n_338),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_L g756 ( 
.A(n_699),
.B(n_562),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_645),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_614),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_712),
.B(n_683),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_613),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_691),
.B(n_562),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_686),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_620),
.B(n_563),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_718),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_723),
.B(n_530),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_620),
.B(n_530),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_689),
.B(n_531),
.Y(n_767)
);

BUFx12f_ASAP7_75t_L g768 ( 
.A(n_594),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_718),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_689),
.Y(n_770)
);

INVx8_ASAP7_75t_L g771 ( 
.A(n_615),
.Y(n_771)
);

AND2x6_ASAP7_75t_L g772 ( 
.A(n_631),
.B(n_248),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_614),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_696),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_722),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_605),
.B(n_317),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_692),
.B(n_531),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_581),
.B(n_321),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_722),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_712),
.B(n_352),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_692),
.B(n_536),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_725),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_648),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_SL g784 ( 
.A(n_615),
.B(n_327),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_604),
.B(n_330),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_627),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_592),
.A2(n_576),
.B1(n_332),
.B2(n_323),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_712),
.B(n_352),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_626),
.B(n_352),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_638),
.B(n_641),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_693),
.B(n_703),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_679),
.B(n_352),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_619),
.B(n_352),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_602),
.B(n_334),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_693),
.B(n_536),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_694),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_703),
.B(n_540),
.Y(n_797)
);

O2A1O1Ixp5_ASAP7_75t_L g798 ( 
.A1(n_654),
.A2(n_705),
.B(n_714),
.C(n_680),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_613),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_641),
.B(n_352),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_705),
.B(n_540),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_704),
.B(n_339),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_641),
.B(n_563),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_714),
.B(n_498),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_591),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_591),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_593),
.Y(n_807)
);

AND2x2_ASAP7_75t_SL g808 ( 
.A(n_635),
.B(n_596),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_610),
.B(n_352),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_648),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_592),
.B(n_506),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_610),
.B(n_352),
.Y(n_812)
);

NOR2xp67_ASAP7_75t_L g813 ( 
.A(n_694),
.B(n_566),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_658),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_719),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_673),
.B(n_342),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_583),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_595),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_595),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_676),
.Y(n_820)
);

NOR2xp67_ASAP7_75t_L g821 ( 
.A(n_650),
.B(n_566),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_621),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_583),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_676),
.B(n_506),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_584),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_621),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_597),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_652),
.B(n_506),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_SL g829 ( 
.A1(n_636),
.A2(n_340),
.B1(n_382),
.B2(n_378),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_673),
.B(n_358),
.Y(n_830)
);

NOR2xp67_ASAP7_75t_L g831 ( 
.A(n_642),
.B(n_594),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_584),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_663),
.B(n_506),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_609),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_682),
.B(n_359),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_716),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_675),
.B(n_506),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_606),
.B(n_506),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_660),
.B(n_569),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_612),
.B(n_523),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_651),
.B(n_343),
.Y(n_841)
);

BUFx5_ASAP7_75t_L g842 ( 
.A(n_716),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_607),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_589),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_617),
.B(n_523),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_618),
.B(n_523),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_598),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_660),
.Y(n_848)
);

O2A1O1Ixp5_ASAP7_75t_L g849 ( 
.A1(n_654),
.A2(n_285),
.B(n_391),
.C(n_390),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_621),
.A2(n_285),
.B1(n_391),
.B2(n_390),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_596),
.A2(n_360),
.B1(n_361),
.B2(n_388),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_621),
.Y(n_852)
);

BUFx8_ASAP7_75t_L g853 ( 
.A(n_615),
.Y(n_853)
);

INVx5_ASAP7_75t_L g854 ( 
.A(n_580),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_585),
.B(n_523),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_585),
.B(n_523),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_585),
.B(n_523),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_682),
.B(n_365),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_685),
.B(n_366),
.Y(n_859)
);

NOR3xp33_ASAP7_75t_L g860 ( 
.A(n_659),
.B(n_345),
.C(n_344),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_685),
.B(n_367),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_655),
.Y(n_862)
);

BUFx12f_ASAP7_75t_SL g863 ( 
.A(n_670),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_687),
.B(n_368),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_687),
.B(n_375),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_598),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_601),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_601),
.Y(n_868)
);

OA21x2_ASAP7_75t_L g869 ( 
.A1(n_706),
.A2(n_534),
.B(n_577),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_587),
.B(n_249),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_670),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_603),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_587),
.B(n_269),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_599),
.B(n_269),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_599),
.B(n_271),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_667),
.B(n_351),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_599),
.B(n_271),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_600),
.B(n_272),
.Y(n_878)
);

INVx8_ASAP7_75t_L g879 ( 
.A(n_611),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_670),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_600),
.B(n_272),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_600),
.B(n_628),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_688),
.B(n_384),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_628),
.B(n_672),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_616),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_623),
.Y(n_886)
);

NOR3xp33_ASAP7_75t_L g887 ( 
.A(n_625),
.B(n_373),
.C(n_381),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_728),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_808),
.B(n_628),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_808),
.B(n_672),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_773),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_728),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_746),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_760),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_738),
.B(n_670),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_737),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_758),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_746),
.B(n_752),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_729),
.B(n_672),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_751),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_763),
.A2(n_721),
.B1(n_636),
.B2(n_726),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_737),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_730),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_774),
.B(n_666),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_741),
.B(n_647),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_731),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_786),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_735),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_869),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_761),
.B(n_678),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_814),
.A2(n_649),
.B1(n_708),
.B2(n_724),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_736),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_741),
.B(n_770),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_841),
.A2(n_701),
.B1(n_717),
.B2(n_721),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_833),
.A2(n_720),
.B(n_690),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_791),
.B(n_678),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_834),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_862),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_863),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_766),
.B(n_695),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_826),
.B(n_695),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_852),
.B(n_871),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_837),
.A2(n_840),
.B(n_838),
.Y(n_923)
);

NOR2x1p5_ASAP7_75t_L g924 ( 
.A(n_848),
.B(n_611),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_739),
.B(n_695),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_744),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_822),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_744),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_753),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_752),
.B(n_656),
.Y(n_930)
);

AO22x1_ASAP7_75t_L g931 ( 
.A1(n_802),
.A2(n_710),
.B1(n_707),
.B2(n_386),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_745),
.B(n_623),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_841),
.A2(n_880),
.B1(n_778),
.B2(n_876),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_869),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_834),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_869),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_764),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_764),
.Y(n_938)
);

INVx4_ASAP7_75t_L g939 ( 
.A(n_760),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_769),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_769),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_796),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_848),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_740),
.B(n_702),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_776),
.B(n_726),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_SL g946 ( 
.A1(n_778),
.A2(n_710),
.B1(n_707),
.B2(n_721),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_SL g947 ( 
.A1(n_829),
.A2(n_655),
.B1(n_721),
.B2(n_374),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_757),
.B(n_634),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_775),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_879),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_762),
.B(n_634),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_775),
.Y(n_952)
);

OR2x4_ASAP7_75t_L g953 ( 
.A(n_802),
.B(n_432),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_803),
.B(n_657),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_754),
.B(n_657),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_743),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_779),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_779),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_790),
.B(n_815),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_805),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_776),
.B(n_661),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_740),
.B(n_702),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_813),
.B(n_688),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_783),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_806),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_783),
.Y(n_966)
);

INVx1_ASAP7_75t_SL g967 ( 
.A(n_839),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_756),
.B(n_700),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_748),
.B(n_665),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_807),
.B(n_706),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_794),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_SL g972 ( 
.A1(n_794),
.A2(n_458),
.B1(n_433),
.B2(n_442),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_818),
.B(n_709),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_821),
.B(n_700),
.Y(n_974)
);

CKINVDCx11_ASAP7_75t_R g975 ( 
.A(n_768),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_819),
.B(n_709),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_827),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_768),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_810),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_785),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_843),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_810),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_787),
.A2(n_669),
.B1(n_279),
.B2(n_387),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_820),
.B(n_571),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_785),
.B(n_711),
.Y(n_985)
);

INVx5_ASAP7_75t_L g986 ( 
.A(n_834),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_782),
.B(n_571),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_885),
.B(n_711),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_886),
.B(n_603),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_732),
.B(n_577),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_876),
.A2(n_275),
.B(n_290),
.C(n_307),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_SL g992 ( 
.A1(n_733),
.A2(n_469),
.B1(n_464),
.B2(n_463),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_820),
.B(n_624),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_879),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_817),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_760),
.B(n_579),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_750),
.B(n_624),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_817),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_SL g999 ( 
.A1(n_772),
.A2(n_385),
.B1(n_290),
.B2(n_307),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_842),
.B(n_609),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_SL g1001 ( 
.A(n_850),
.B(n_755),
.C(n_734),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_772),
.Y(n_1002)
);

NAND2xp33_ASAP7_75t_L g1003 ( 
.A(n_799),
.B(n_609),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_853),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_834),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_772),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_747),
.A2(n_669),
.B1(n_310),
.B2(n_322),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_772),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_823),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_816),
.A2(n_669),
.B1(n_664),
.B2(n_727),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_765),
.B(n_629),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_842),
.B(n_609),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_836),
.B(n_629),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_825),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_799),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_825),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_832),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_836),
.B(n_630),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_799),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_832),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_831),
.Y(n_1021)
);

NAND2x1p5_ASAP7_75t_L g1022 ( 
.A(n_799),
.B(n_720),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_844),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_771),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_784),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_844),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_759),
.B(n_767),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_847),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_860),
.B(n_433),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_847),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_866),
.Y(n_1031)
);

NAND2x1p5_ASAP7_75t_L g1032 ( 
.A(n_759),
.B(n_720),
.Y(n_1032)
);

NAND2x1p5_ASAP7_75t_L g1033 ( 
.A(n_742),
.B(n_609),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_771),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_777),
.B(n_630),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_781),
.B(n_632),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_842),
.B(n_644),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_795),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_866),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_771),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_797),
.B(n_632),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_801),
.B(n_633),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_867),
.Y(n_1043)
);

INVx5_ASAP7_75t_L g1044 ( 
.A(n_854),
.Y(n_1044)
);

BUFx12f_ASAP7_75t_L g1045 ( 
.A(n_853),
.Y(n_1045)
);

OR2x6_ASAP7_75t_L g1046 ( 
.A(n_742),
.B(n_275),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_867),
.Y(n_1047)
);

INVx4_ASAP7_75t_L g1048 ( 
.A(n_842),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_816),
.A2(n_633),
.B1(n_640),
.B2(n_323),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_868),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_868),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_747),
.A2(n_310),
.B1(n_322),
.B2(n_328),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_887),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_872),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_830),
.Y(n_1055)
);

AOI21xp33_ASAP7_75t_L g1056 ( 
.A1(n_835),
.A2(n_328),
.B(n_329),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_804),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_882),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_888),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_888),
.Y(n_1060)
);

OR2x6_ASAP7_75t_L g1061 ( 
.A(n_950),
.B(n_809),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1038),
.B(n_749),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1028),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_945),
.B(n_789),
.Y(n_1064)
);

NAND2x1p5_ASAP7_75t_L g1065 ( 
.A(n_986),
.B(n_809),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_933),
.A2(n_811),
.B1(n_734),
.B2(n_884),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1048),
.A2(n_1044),
.B(n_923),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1038),
.B(n_913),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1048),
.A2(n_1044),
.B(n_986),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_891),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_907),
.B(n_789),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_945),
.B(n_792),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_892),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_905),
.A2(n_798),
.B(n_793),
.C(n_792),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_975),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1044),
.A2(n_846),
.B(n_845),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_971),
.B(n_851),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_900),
.B(n_967),
.Y(n_1078)
);

O2A1O1Ixp5_ASAP7_75t_SL g1079 ( 
.A1(n_974),
.A2(n_793),
.B(n_864),
.C(n_861),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_896),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1028),
.Y(n_1081)
);

OAI21xp33_ASAP7_75t_L g1082 ( 
.A1(n_905),
.A2(n_858),
.B(n_835),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_897),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_991),
.A2(n_812),
.B(n_865),
.C(n_864),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_991),
.A2(n_812),
.B(n_865),
.C(n_861),
.Y(n_1085)
);

OAI21xp33_ASAP7_75t_SL g1086 ( 
.A1(n_983),
.A2(n_883),
.B(n_858),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1044),
.A2(n_854),
.B(n_828),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_986),
.A2(n_854),
.B(n_824),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_943),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_895),
.A2(n_870),
.B1(n_881),
.B2(n_878),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_986),
.A2(n_854),
.B(n_856),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_904),
.B(n_859),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_902),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_917),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_904),
.B(n_859),
.Y(n_1095)
);

INVx6_ASAP7_75t_L g1096 ( 
.A(n_1024),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_942),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_956),
.B(n_883),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_943),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_930),
.Y(n_1100)
);

INVxp67_ASAP7_75t_SL g1101 ( 
.A(n_917),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_SL g1102 ( 
.A(n_978),
.B(n_337),
.Y(n_1102)
);

OAI22x1_ASAP7_75t_L g1103 ( 
.A1(n_962),
.A2(n_1053),
.B1(n_1025),
.B2(n_927),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_914),
.A2(n_877),
.B1(n_875),
.B2(n_874),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_944),
.B(n_987),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1050),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_1034),
.Y(n_1107)
);

NOR2xp67_ASAP7_75t_L g1108 ( 
.A(n_1021),
.B(n_800),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1056),
.A2(n_780),
.B(n_788),
.C(n_873),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1003),
.A2(n_857),
.B(n_855),
.Y(n_1110)
);

NOR2xp67_ASAP7_75t_SL g1111 ( 
.A(n_950),
.B(n_800),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1027),
.A2(n_849),
.B(n_780),
.C(n_788),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1050),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_961),
.A2(n_337),
.B1(n_355),
.B2(n_387),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1034),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1027),
.A2(n_355),
.B(n_389),
.C(n_477),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1054),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_901),
.B(n_442),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_962),
.B(n_842),
.Y(n_1119)
);

AOI221xp5_ASAP7_75t_L g1120 ( 
.A1(n_931),
.A2(n_452),
.B1(n_450),
.B2(n_449),
.C(n_494),
.Y(n_1120)
);

NOR2xp67_ASAP7_75t_L g1121 ( 
.A(n_1024),
.B(n_73),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1040),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_918),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_899),
.A2(n_690),
.B(n_527),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_927),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_946),
.A2(n_458),
.B1(n_454),
.B2(n_452),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_990),
.B(n_644),
.Y(n_1127)
);

OAI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_953),
.A2(n_454),
.B1(n_450),
.B2(n_449),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_964),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1029),
.B(n_461),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_903),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_SL g1132 ( 
.A1(n_972),
.A2(n_479),
.B1(n_492),
.B2(n_462),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_954),
.B(n_644),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_955),
.A2(n_478),
.B(n_491),
.C(n_462),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_906),
.B(n_644),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_983),
.A2(n_662),
.B1(n_697),
.B2(n_690),
.Y(n_1136)
);

INVxp33_ASAP7_75t_L g1137 ( 
.A(n_947),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_908),
.B(n_662),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_975),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_932),
.A2(n_479),
.B(n_490),
.C(n_464),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_985),
.A2(n_662),
.B1(n_697),
.B2(n_690),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_912),
.B(n_662),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_919),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1057),
.B(n_697),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1055),
.A2(n_697),
.B1(n_482),
.B2(n_469),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_984),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1000),
.A2(n_527),
.B(n_608),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_985),
.B(n_960),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1001),
.A2(n_481),
.B(n_490),
.C(n_470),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1001),
.A2(n_491),
.B(n_486),
.C(n_483),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_893),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_984),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_911),
.A2(n_486),
.B(n_483),
.C(n_482),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1045),
.Y(n_1154)
);

AND2x6_ASAP7_75t_SL g1155 ( 
.A(n_959),
.B(n_898),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1040),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_SL g1157 ( 
.A(n_1045),
.B(n_475),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_965),
.B(n_475),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_917),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_SL g1160 ( 
.A1(n_1002),
.A2(n_411),
.B(n_409),
.C(n_191),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_1019),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_893),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_901),
.B(n_411),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_977),
.B(n_0),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_926),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_959),
.B(n_608),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1004),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1012),
.A2(n_1037),
.B(n_916),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1010),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_981),
.B(n_4),
.Y(n_1170)
);

OR2x6_ASAP7_75t_L g1171 ( 
.A(n_994),
.B(n_713),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1012),
.A2(n_713),
.B(n_189),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_889),
.B(n_8),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_889),
.B(n_8),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_890),
.B(n_10),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1006),
.A2(n_11),
.B(n_14),
.C(n_16),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_996),
.B(n_17),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1033),
.A2(n_184),
.B1(n_177),
.B2(n_175),
.Y(n_1178)
);

INVx4_ASAP7_75t_L g1179 ( 
.A(n_1019),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_997),
.B(n_17),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_999),
.B(n_20),
.C(n_22),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_928),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1011),
.B(n_20),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_948),
.A2(n_22),
.B(n_25),
.C(n_26),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_1019),
.B(n_148),
.Y(n_1185)
);

AOI21x1_ASAP7_75t_L g1186 ( 
.A1(n_890),
.A2(n_147),
.B(n_138),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1035),
.B(n_1036),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1007),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1041),
.B(n_29),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1058),
.B(n_132),
.Y(n_1190)
);

AO32x2_ASAP7_75t_L g1191 ( 
.A1(n_1008),
.A2(n_30),
.A3(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_929),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_924),
.B(n_35),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1074),
.A2(n_915),
.A3(n_909),
.B(n_936),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1068),
.B(n_1042),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1060),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1148),
.B(n_920),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1129),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1086),
.A2(n_1007),
.B(n_969),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1067),
.A2(n_1013),
.B(n_1018),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1110),
.A2(n_1032),
.B(n_974),
.Y(n_1201)
);

NAND2x1p5_ASAP7_75t_L g1202 ( 
.A(n_1161),
.B(n_939),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1168),
.A2(n_1032),
.B(n_936),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1076),
.A2(n_968),
.B(n_963),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1131),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1079),
.A2(n_1049),
.B(n_968),
.Y(n_1206)
);

AOI221x1_ASAP7_75t_L g1207 ( 
.A1(n_1169),
.A2(n_992),
.B1(n_1058),
.B2(n_993),
.C(n_949),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1092),
.A2(n_1095),
.B(n_1072),
.C(n_1064),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1187),
.A2(n_1104),
.B(n_1119),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1066),
.A2(n_909),
.A3(n_934),
.B(n_937),
.Y(n_1210)
);

INVx5_ASAP7_75t_L g1211 ( 
.A(n_1094),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1095),
.B(n_951),
.Y(n_1212)
);

OAI22x1_ASAP7_75t_L g1213 ( 
.A1(n_1064),
.A2(n_922),
.B1(n_921),
.B2(n_1033),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1119),
.A2(n_1022),
.B(n_910),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1069),
.A2(n_934),
.B(n_937),
.Y(n_1215)
);

INVx3_ASAP7_75t_SL g1216 ( 
.A(n_1154),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1091),
.A2(n_952),
.B(n_970),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1072),
.B(n_952),
.Y(n_1218)
);

AO21x1_ASAP7_75t_L g1219 ( 
.A1(n_1173),
.A2(n_910),
.B(n_963),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1165),
.Y(n_1220)
);

AOI221xp5_ASAP7_75t_L g1221 ( 
.A1(n_1126),
.A2(n_1052),
.B1(n_989),
.B2(n_925),
.C(n_921),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1112),
.A2(n_973),
.B(n_976),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1130),
.B(n_1058),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1090),
.A2(n_1022),
.B(n_1005),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1082),
.A2(n_1052),
.B(n_941),
.C(n_958),
.Y(n_1225)
);

O2A1O1Ixp5_ASAP7_75t_SL g1226 ( 
.A1(n_1114),
.A2(n_938),
.B(n_957),
.C(n_940),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1149),
.A2(n_1150),
.B(n_1085),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1062),
.B(n_1020),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1088),
.A2(n_988),
.B(n_1051),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1087),
.A2(n_1020),
.B(n_1051),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1186),
.A2(n_1017),
.B(n_1047),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1137),
.A2(n_1046),
.B1(n_894),
.B2(n_1015),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1078),
.B(n_1046),
.Y(n_1233)
);

INVx2_ASAP7_75t_SL g1234 ( 
.A(n_1070),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1116),
.A2(n_1047),
.A3(n_966),
.B(n_979),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1083),
.Y(n_1236)
);

AOI221xp5_ASAP7_75t_SL g1237 ( 
.A1(n_1188),
.A2(n_995),
.B1(n_1043),
.B2(n_998),
.C(n_1031),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1084),
.A2(n_1174),
.B(n_1173),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1126),
.B(n_982),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1189),
.A2(n_1014),
.B(n_1009),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1109),
.A2(n_917),
.B(n_935),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1124),
.A2(n_1016),
.B(n_1039),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_1139),
.Y(n_1243)
);

NOR2xp67_ASAP7_75t_SL g1244 ( 
.A(n_1075),
.B(n_1005),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1098),
.B(n_1016),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1174),
.B(n_982),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1127),
.A2(n_935),
.B(n_1005),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1133),
.A2(n_935),
.B(n_1005),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1146),
.B(n_1046),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1141),
.A2(n_935),
.B(n_939),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_1125),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1182),
.Y(n_1252)
);

NAND2x1p5_ASAP7_75t_L g1253 ( 
.A(n_1161),
.B(n_894),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1192),
.Y(n_1254)
);

AOI21xp33_ASAP7_75t_L g1255 ( 
.A1(n_1175),
.A2(n_1030),
.B(n_1026),
.Y(n_1255)
);

NAND2x1p5_ASAP7_75t_L g1256 ( 
.A(n_1179),
.B(n_1023),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1147),
.A2(n_1017),
.B(n_116),
.Y(n_1257)
);

AOI221xp5_ASAP7_75t_SL g1258 ( 
.A1(n_1128),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.C(n_42),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_SL g1259 ( 
.A1(n_1101),
.A2(n_105),
.B(n_103),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1146),
.B(n_37),
.Y(n_1260)
);

INVxp67_ASAP7_75t_SL g1261 ( 
.A(n_1101),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1175),
.B(n_42),
.Y(n_1262)
);

OAI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1118),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_1263)
);

AOI21x1_ASAP7_75t_SL g1264 ( 
.A1(n_1180),
.A2(n_1183),
.B(n_1164),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1172),
.A2(n_101),
.B(n_92),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1077),
.A2(n_89),
.B(n_85),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1071),
.B(n_48),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1136),
.A2(n_83),
.B(n_53),
.Y(n_1268)
);

NAND2x1_ASAP7_75t_L g1269 ( 
.A(n_1096),
.B(n_52),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1089),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1144),
.A2(n_54),
.B(n_57),
.Y(n_1271)
);

AND3x4_ASAP7_75t_L g1272 ( 
.A(n_1099),
.B(n_59),
.C(n_62),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1152),
.B(n_65),
.Y(n_1273)
);

NOR4xp25_ASAP7_75t_L g1274 ( 
.A(n_1184),
.B(n_70),
.C(n_71),
.D(n_1176),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1059),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1083),
.Y(n_1276)
);

NOR2x1_ASAP7_75t_SL g1277 ( 
.A(n_1171),
.B(n_1061),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1107),
.Y(n_1278)
);

O2A1O1Ixp5_ASAP7_75t_L g1279 ( 
.A1(n_1111),
.A2(n_1190),
.B(n_1163),
.C(n_1160),
.Y(n_1279)
);

O2A1O1Ixp5_ASAP7_75t_SL g1280 ( 
.A1(n_1185),
.A2(n_1080),
.B(n_1073),
.C(n_1093),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1135),
.A2(n_1142),
.B(n_1138),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1097),
.A2(n_1108),
.B1(n_1103),
.B2(n_1152),
.Y(n_1282)
);

INVx3_ASAP7_75t_SL g1283 ( 
.A(n_1167),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1065),
.A2(n_1117),
.B(n_1063),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1065),
.A2(n_1106),
.B(n_1081),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1113),
.Y(n_1286)
);

AO32x2_ASAP7_75t_L g1287 ( 
.A1(n_1178),
.A2(n_1191),
.A3(n_1179),
.B1(n_1160),
.B2(n_1123),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1166),
.A2(n_1061),
.B(n_1158),
.Y(n_1288)
);

XNOR2xp5_ASAP7_75t_L g1289 ( 
.A(n_1143),
.B(n_1100),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1177),
.B(n_1151),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1061),
.A2(n_1121),
.B(n_1159),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1094),
.A2(n_1159),
.B(n_1171),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1094),
.A2(n_1159),
.B(n_1171),
.Y(n_1293)
);

CKINVDCx14_ASAP7_75t_R g1294 ( 
.A(n_1162),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1155),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1132),
.A2(n_1170),
.B1(n_1181),
.B2(n_1145),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1132),
.A2(n_1170),
.B1(n_1153),
.B2(n_1096),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1159),
.A2(n_1140),
.B(n_1134),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1096),
.A2(n_1120),
.B1(n_1191),
.B2(n_1193),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1115),
.Y(n_1300)
);

AOI21xp33_ASAP7_75t_L g1301 ( 
.A1(n_1102),
.A2(n_1157),
.B(n_1191),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1122),
.A2(n_1156),
.B(n_1191),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1092),
.A2(n_905),
.B(n_1095),
.C(n_1072),
.Y(n_1303)
);

AO22x2_ASAP7_75t_L g1304 ( 
.A1(n_1181),
.A2(n_1118),
.B1(n_980),
.B2(n_971),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1068),
.B(n_1038),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1131),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1074),
.A2(n_1086),
.B(n_1079),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1068),
.B(n_1148),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1131),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1068),
.B(n_1148),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1068),
.B(n_1148),
.Y(n_1311)
);

BUFx10_ASAP7_75t_L g1312 ( 
.A(n_1167),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1064),
.A2(n_945),
.B1(n_905),
.B2(n_1072),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1068),
.B(n_1148),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1105),
.B(n_1130),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1064),
.A2(n_945),
.B1(n_905),
.B2(n_1072),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1060),
.Y(n_1317)
);

AO32x2_ASAP7_75t_L g1318 ( 
.A1(n_1066),
.A2(n_1114),
.A3(n_972),
.B1(n_850),
.B2(n_1104),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1074),
.A2(n_1086),
.B(n_1079),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1068),
.B(n_1148),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1131),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1152),
.B(n_1146),
.Y(n_1322)
);

AOI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1067),
.A2(n_1076),
.B(n_923),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1074),
.A2(n_1104),
.A3(n_1066),
.B(n_1149),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1064),
.B(n_945),
.Y(n_1325)
);

AO31x2_ASAP7_75t_L g1326 ( 
.A1(n_1074),
.A2(n_1104),
.A3(n_1066),
.B(n_1149),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1105),
.B(n_980),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_SL g1328 ( 
.A1(n_1137),
.A2(n_945),
.B(n_946),
.Y(n_1328)
);

O2A1O1Ixp5_ASAP7_75t_SL g1329 ( 
.A1(n_1114),
.A2(n_747),
.B(n_1190),
.C(n_792),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1068),
.B(n_586),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1105),
.B(n_980),
.Y(n_1331)
);

AO32x2_ASAP7_75t_L g1332 ( 
.A1(n_1066),
.A2(n_1114),
.A3(n_972),
.B1(n_850),
.B2(n_1104),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1313),
.B(n_1316),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1261),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1211),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1257),
.A2(n_1201),
.B(n_1323),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1328),
.B(n_1330),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1307),
.A2(n_1319),
.B(n_1238),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1262),
.A2(n_1296),
.B1(n_1304),
.B2(n_1263),
.Y(n_1339)
);

AO31x2_ASAP7_75t_L g1340 ( 
.A1(n_1219),
.A2(n_1207),
.A3(n_1213),
.B(n_1209),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1199),
.A2(n_1301),
.B(n_1266),
.C(n_1227),
.Y(n_1341)
);

AO21x2_ASAP7_75t_L g1342 ( 
.A1(n_1307),
.A2(n_1319),
.B(n_1199),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1315),
.B(n_1290),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1328),
.B(n_1327),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1308),
.A2(n_1311),
.B1(n_1320),
.B2(n_1310),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1211),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1331),
.B(n_1212),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1262),
.A2(n_1296),
.B1(n_1304),
.B2(n_1301),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1272),
.A2(n_1297),
.B1(n_1227),
.B2(n_1266),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1297),
.A2(n_1195),
.B1(n_1314),
.B2(n_1320),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1200),
.A2(n_1242),
.B(n_1217),
.Y(n_1351)
);

AO31x2_ASAP7_75t_L g1352 ( 
.A1(n_1214),
.A2(n_1241),
.A3(n_1299),
.B(n_1224),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1206),
.A2(n_1237),
.B(n_1222),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1211),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1322),
.B(n_1277),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1305),
.B(n_1195),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1229),
.A2(n_1204),
.B(n_1203),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1223),
.B(n_1197),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1306),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1206),
.A2(n_1237),
.B(n_1222),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1279),
.A2(n_1255),
.B(n_1271),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1309),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1233),
.B(n_1249),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1236),
.Y(n_1364)
);

NOR2xp67_ASAP7_75t_L g1365 ( 
.A(n_1234),
.B(n_1251),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1230),
.A2(n_1231),
.B(n_1215),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1299),
.A2(n_1282),
.B1(n_1197),
.B2(n_1269),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1321),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_SL g1369 ( 
.A(n_1283),
.B(n_1243),
.Y(n_1369)
);

AOI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1240),
.A2(n_1298),
.B(n_1281),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1276),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1196),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1329),
.A2(n_1265),
.B(n_1226),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1264),
.A2(n_1250),
.B(n_1248),
.Y(n_1374)
);

NOR2xp67_ASAP7_75t_L g1375 ( 
.A(n_1289),
.B(n_1300),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1280),
.A2(n_1247),
.B(n_1284),
.Y(n_1376)
);

A2O1A1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1268),
.A2(n_1258),
.B(n_1302),
.C(n_1221),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1198),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1267),
.B(n_1273),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1235),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1285),
.A2(n_1292),
.B(n_1293),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1274),
.A2(n_1246),
.B(n_1218),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1294),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1260),
.B(n_1286),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1295),
.A2(n_1216),
.B1(n_1232),
.B2(n_1278),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1220),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1228),
.A2(n_1245),
.B(n_1256),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1312),
.A2(n_1254),
.B1(n_1252),
.B2(n_1239),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1228),
.A2(n_1256),
.B(n_1253),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1317),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1270),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1253),
.A2(n_1202),
.B(n_1259),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1258),
.B(n_1225),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1318),
.A2(n_1332),
.B(n_1326),
.Y(n_1394)
);

BUFx12f_ASAP7_75t_L g1395 ( 
.A(n_1312),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1332),
.A2(n_1324),
.B1(n_1326),
.B2(n_1287),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1235),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1210),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1194),
.A2(n_1210),
.B(n_1324),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1324),
.B(n_1326),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1332),
.A2(n_1287),
.B(n_1210),
.C(n_1194),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1287),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_1289),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1257),
.A2(n_1201),
.B(n_1323),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_1289),
.Y(n_1405)
);

BUFx5_ASAP7_75t_L g1406 ( 
.A(n_1220),
.Y(n_1406)
);

OR2x6_ASAP7_75t_L g1407 ( 
.A(n_1291),
.B(n_1288),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1307),
.A2(n_1319),
.B(n_1238),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1257),
.A2(n_1201),
.B(n_1323),
.Y(n_1409)
);

INVxp67_ASAP7_75t_L g1410 ( 
.A(n_1236),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1315),
.B(n_1290),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1275),
.Y(n_1412)
);

OAI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1313),
.A2(n_1316),
.B1(n_945),
.B2(n_1325),
.Y(n_1413)
);

AOI221xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1303),
.A2(n_945),
.B1(n_1208),
.B2(n_1325),
.C(n_1296),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1307),
.A2(n_1319),
.B(n_1238),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1205),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1303),
.A2(n_945),
.B(n_1325),
.C(n_905),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1313),
.A2(n_1316),
.B1(n_945),
.B2(n_1325),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_SL g1419 ( 
.A1(n_1277),
.A2(n_1227),
.B(n_1291),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1205),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1315),
.B(n_1290),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1257),
.A2(n_1201),
.B(n_1323),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1257),
.A2(n_1201),
.B(n_1323),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1315),
.B(n_1290),
.Y(n_1424)
);

NAND2x1p5_ASAP7_75t_L g1425 ( 
.A(n_1211),
.B(n_1244),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1313),
.B(n_945),
.C(n_905),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1243),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1205),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1257),
.A2(n_1201),
.B(n_1323),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1205),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1243),
.Y(n_1431)
);

OAI22x1_ASAP7_75t_L g1432 ( 
.A1(n_1313),
.A2(n_1316),
.B1(n_1325),
.B2(n_945),
.Y(n_1432)
);

OAI21xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1238),
.A2(n_933),
.B(n_1313),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1205),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1325),
.A2(n_945),
.B1(n_1316),
.B2(n_1313),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1307),
.A2(n_1319),
.B(n_1238),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1205),
.Y(n_1437)
);

OAI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1303),
.A2(n_1316),
.B(n_1313),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1313),
.A2(n_1316),
.B1(n_945),
.B2(n_1325),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1313),
.A2(n_1316),
.B1(n_945),
.B2(n_1325),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1307),
.A2(n_1319),
.B(n_1238),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1211),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1236),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1325),
.B(n_1313),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1325),
.B(n_1313),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1303),
.A2(n_1316),
.B(n_1313),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1205),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1305),
.B(n_1330),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1205),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1325),
.A2(n_945),
.B1(n_1316),
.B2(n_1313),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1257),
.A2(n_1201),
.B(n_1323),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1325),
.B(n_1313),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1211),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1257),
.A2(n_1201),
.B(n_1323),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1307),
.A2(n_1319),
.B(n_1199),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1313),
.A2(n_1316),
.B1(n_945),
.B2(n_1325),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1313),
.B(n_1316),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1322),
.B(n_1277),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1322),
.B(n_1277),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1315),
.B(n_1290),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1275),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1243),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1307),
.A2(n_1319),
.B(n_1238),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1313),
.A2(n_1316),
.B1(n_945),
.B2(n_1325),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1322),
.B(n_1277),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1315),
.B(n_1290),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1307),
.A2(n_1319),
.B(n_1238),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_SL g1468 ( 
.A1(n_1303),
.A2(n_1301),
.B(n_1169),
.C(n_1188),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1325),
.A2(n_945),
.B1(n_1316),
.B2(n_1313),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_1261),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1325),
.A2(n_945),
.B1(n_1316),
.B2(n_1313),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1257),
.A2(n_1201),
.B(n_1323),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1313),
.A2(n_1316),
.B1(n_945),
.B2(n_1325),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1313),
.A2(n_1316),
.B1(n_945),
.B2(n_1325),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1307),
.A2(n_1319),
.B(n_1238),
.Y(n_1475)
);

INVx8_ASAP7_75t_L g1476 ( 
.A(n_1211),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1363),
.B(n_1343),
.Y(n_1477)
);

BUFx2_ASAP7_75t_R g1478 ( 
.A(n_1427),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1355),
.B(n_1458),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1345),
.B(n_1350),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1448),
.B(n_1379),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1413),
.B(n_1473),
.Y(n_1482)
);

NOR2xp67_ASAP7_75t_R g1483 ( 
.A(n_1395),
.B(n_1383),
.Y(n_1483)
);

AOI21x1_ASAP7_75t_SL g1484 ( 
.A1(n_1444),
.A2(n_1452),
.B(n_1445),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1435),
.A2(n_1450),
.B1(n_1469),
.B2(n_1349),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1411),
.B(n_1421),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1364),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1350),
.B(n_1333),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1371),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1457),
.B(n_1438),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1446),
.B(n_1424),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1395),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1427),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1460),
.B(n_1466),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1435),
.A2(n_1450),
.B1(n_1469),
.B2(n_1349),
.Y(n_1495)
);

OR2x6_ASAP7_75t_L g1496 ( 
.A(n_1407),
.B(n_1419),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1426),
.B(n_1418),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1373),
.A2(n_1366),
.B(n_1377),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1471),
.A2(n_1439),
.B1(n_1474),
.B2(n_1440),
.Y(n_1499)
);

NOR2xp67_ASAP7_75t_L g1500 ( 
.A(n_1410),
.B(n_1443),
.Y(n_1500)
);

O2A1O1Ixp5_ASAP7_75t_L g1501 ( 
.A1(n_1393),
.A2(n_1341),
.B(n_1377),
.C(n_1456),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1358),
.B(n_1337),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1333),
.B(n_1356),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1347),
.B(n_1414),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1347),
.B(n_1382),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1334),
.A2(n_1470),
.B(n_1464),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1391),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1373),
.A2(n_1366),
.B(n_1351),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1337),
.B(n_1348),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1384),
.B(n_1344),
.Y(n_1510)
);

A2O1A1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1433),
.A2(n_1344),
.B(n_1341),
.C(n_1339),
.Y(n_1511)
);

O2A1O1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1468),
.A2(n_1393),
.B(n_1339),
.C(n_1367),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1348),
.B(n_1432),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_SL g1514 ( 
.A1(n_1425),
.A2(n_1335),
.B(n_1346),
.Y(n_1514)
);

BUFx4f_ASAP7_75t_SL g1515 ( 
.A(n_1431),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1385),
.A2(n_1388),
.B1(n_1365),
.B2(n_1403),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1394),
.B(n_1338),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1405),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1355),
.B(n_1458),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1375),
.A2(n_1459),
.B1(n_1465),
.B2(n_1425),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1431),
.A2(n_1462),
.B1(n_1407),
.B2(n_1459),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1335),
.A2(n_1346),
.B(n_1407),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1338),
.B(n_1408),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1462),
.A2(n_1465),
.B1(n_1449),
.B2(n_1386),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1359),
.A2(n_1437),
.B1(n_1416),
.B2(n_1420),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1362),
.A2(n_1430),
.B1(n_1434),
.B2(n_1368),
.Y(n_1526)
);

OR2x6_ASAP7_75t_L g1527 ( 
.A(n_1476),
.B(n_1381),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1338),
.B(n_1408),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1412),
.B(n_1461),
.Y(n_1529)
);

AOI211xp5_ASAP7_75t_L g1530 ( 
.A1(n_1428),
.A2(n_1447),
.B(n_1369),
.C(n_1401),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1372),
.B(n_1378),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1376),
.A2(n_1399),
.B(n_1357),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1408),
.B(n_1415),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1390),
.B(n_1406),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1415),
.B(n_1436),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1415),
.B(n_1436),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1389),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1400),
.B(n_1467),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1453),
.B(n_1354),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1335),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1342),
.A2(n_1455),
.B(n_1475),
.C(n_1467),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1436),
.B(n_1441),
.Y(n_1542)
);

OAI22x1_ASAP7_75t_L g1543 ( 
.A1(n_1441),
.A2(n_1467),
.B1(n_1463),
.B2(n_1402),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1441),
.B(n_1463),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1396),
.A2(n_1463),
.B1(n_1453),
.B2(n_1354),
.Y(n_1545)
);

O2A1O1Ixp5_ASAP7_75t_L g1546 ( 
.A1(n_1370),
.A2(n_1398),
.B(n_1380),
.C(n_1397),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1342),
.B(n_1455),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1442),
.B(n_1406),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1406),
.B(n_1396),
.Y(n_1549)
);

AOI211xp5_ASAP7_75t_L g1550 ( 
.A1(n_1374),
.A2(n_1402),
.B(n_1381),
.C(n_1389),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1346),
.A2(n_1476),
.B1(n_1360),
.B2(n_1353),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1387),
.B(n_1340),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1399),
.A2(n_1357),
.B(n_1422),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1476),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1352),
.B(n_1361),
.Y(n_1555)
);

O2A1O1Ixp33_ASAP7_75t_L g1556 ( 
.A1(n_1336),
.A2(n_1404),
.B(n_1409),
.C(n_1422),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1423),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1429),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1559)
);

O2A1O1Ixp33_ASAP7_75t_L g1560 ( 
.A1(n_1472),
.A2(n_1303),
.B(n_1417),
.C(n_1418),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1335),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1373),
.A2(n_1319),
.B(n_1307),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1435),
.A2(n_945),
.B1(n_1316),
.B2(n_1313),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1363),
.B(n_1343),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1435),
.A2(n_945),
.B1(n_1316),
.B2(n_1313),
.Y(n_1565)
);

NAND2x1p5_ASAP7_75t_L g1566 ( 
.A(n_1392),
.B(n_1389),
.Y(n_1566)
);

AOI211xp5_ASAP7_75t_L g1567 ( 
.A1(n_1426),
.A2(n_945),
.B(n_1325),
.C(n_1413),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1363),
.B(n_1343),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1427),
.Y(n_1569)
);

AOI21xp5_ASAP7_75t_SL g1570 ( 
.A1(n_1417),
.A2(n_1303),
.B(n_1208),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1364),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1448),
.B(n_1379),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1435),
.A2(n_945),
.B1(n_1316),
.B2(n_1313),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1364),
.Y(n_1574)
);

CKINVDCx20_ASAP7_75t_R g1575 ( 
.A(n_1515),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1538),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1544),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1510),
.B(n_1555),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1558),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1543),
.B(n_1517),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1517),
.B(n_1523),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1505),
.B(n_1503),
.Y(n_1582)
);

INVx4_ASAP7_75t_L g1583 ( 
.A(n_1496),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1557),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1537),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1496),
.B(n_1527),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1547),
.B(n_1523),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1528),
.B(n_1533),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1502),
.B(n_1503),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1527),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1552),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1549),
.B(n_1479),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1525),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1489),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1526),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1518),
.B(n_1481),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1528),
.B(n_1533),
.Y(n_1597)
);

OAI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1501),
.A2(n_1497),
.B(n_1482),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1527),
.B(n_1496),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1548),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1553),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1552),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1553),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1535),
.Y(n_1604)
);

NOR2x1_ASAP7_75t_SL g1605 ( 
.A(n_1551),
.B(n_1490),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1505),
.B(n_1480),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1480),
.B(n_1488),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1493),
.Y(n_1608)
);

CKINVDCx14_ASAP7_75t_R g1609 ( 
.A(n_1569),
.Y(n_1609)
);

XNOR2xp5_ASAP7_75t_L g1610 ( 
.A(n_1486),
.B(n_1477),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1571),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1541),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1536),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1519),
.B(n_1562),
.Y(n_1614)
);

OAI21xp33_ASAP7_75t_SL g1615 ( 
.A1(n_1488),
.A2(n_1570),
.B(n_1499),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1536),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1566),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1542),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1498),
.B(n_1550),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1532),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1507),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1534),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1559),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1532),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1545),
.Y(n_1625)
);

BUFx2_ASAP7_75t_SL g1626 ( 
.A(n_1500),
.Y(n_1626)
);

OA21x2_ASAP7_75t_L g1627 ( 
.A1(n_1546),
.A2(n_1511),
.B(n_1513),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1529),
.Y(n_1628)
);

AOI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1485),
.A2(n_1495),
.B1(n_1573),
.B2(n_1563),
.C(n_1565),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1572),
.B(n_1491),
.Y(n_1630)
);

AO21x2_ASAP7_75t_L g1631 ( 
.A1(n_1556),
.A2(n_1560),
.B(n_1513),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1509),
.A2(n_1504),
.B1(n_1521),
.B2(n_1516),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1574),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1508),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1581),
.B(n_1588),
.Y(n_1635)
);

NOR2xp67_ASAP7_75t_L g1636 ( 
.A(n_1616),
.B(n_1487),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1577),
.B(n_1588),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_1599),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1597),
.B(n_1560),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1587),
.B(n_1494),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_SL g1641 ( 
.A(n_1599),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1580),
.B(n_1614),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1580),
.B(n_1531),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1576),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1576),
.B(n_1616),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1613),
.B(n_1530),
.Y(n_1646)
);

OAI221xp5_ASAP7_75t_SL g1647 ( 
.A1(n_1629),
.A2(n_1567),
.B1(n_1512),
.B2(n_1506),
.C(n_1484),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1579),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1613),
.B(n_1512),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1601),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1585),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1585),
.Y(n_1652)
);

OAI21xp33_ASAP7_75t_L g1653 ( 
.A1(n_1598),
.A2(n_1478),
.B(n_1568),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1614),
.B(n_1564),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1618),
.B(n_1520),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1604),
.B(n_1524),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1623),
.B(n_1539),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1603),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_L g1659 ( 
.A(n_1583),
.B(n_1522),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1617),
.Y(n_1660)
);

NAND3xp33_ASAP7_75t_L g1661 ( 
.A(n_1647),
.B(n_1598),
.C(n_1629),
.Y(n_1661)
);

INVxp67_ASAP7_75t_SL g1662 ( 
.A(n_1636),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1646),
.A2(n_1632),
.B1(n_1609),
.B2(n_1627),
.Y(n_1663)
);

OAI211xp5_ASAP7_75t_L g1664 ( 
.A1(n_1647),
.A2(n_1615),
.B(n_1625),
.C(n_1606),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1649),
.A2(n_1610),
.B1(n_1607),
.B2(n_1589),
.Y(n_1665)
);

AND2x4_ASAP7_75t_SL g1666 ( 
.A(n_1657),
.B(n_1586),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1639),
.B(n_1591),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1642),
.B(n_1600),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1648),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1642),
.B(n_1600),
.Y(n_1670)
);

NAND2xp33_ASAP7_75t_SL g1671 ( 
.A(n_1641),
.B(n_1610),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1650),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1649),
.A2(n_1607),
.B1(n_1606),
.B2(n_1582),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1653),
.A2(n_1615),
.B1(n_1582),
.B2(n_1625),
.C(n_1630),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1639),
.B(n_1591),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1639),
.A2(n_1594),
.B1(n_1611),
.B2(n_1612),
.C(n_1633),
.Y(n_1676)
);

CKINVDCx16_ASAP7_75t_R g1677 ( 
.A(n_1641),
.Y(n_1677)
);

NAND4xp25_ASAP7_75t_SL g1678 ( 
.A(n_1646),
.B(n_1478),
.C(n_1575),
.D(n_1619),
.Y(n_1678)
);

OAI33xp33_ASAP7_75t_L g1679 ( 
.A1(n_1651),
.A2(n_1611),
.A3(n_1594),
.B1(n_1602),
.B2(n_1593),
.B3(n_1595),
.Y(n_1679)
);

AOI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1653),
.A2(n_1612),
.B1(n_1633),
.B2(n_1596),
.C(n_1622),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1660),
.Y(n_1681)
);

AOI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1655),
.A2(n_1622),
.B1(n_1593),
.B2(n_1595),
.C(n_1644),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1648),
.Y(n_1683)
);

INVxp67_ASAP7_75t_SL g1684 ( 
.A(n_1636),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1652),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1642),
.B(n_1592),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1652),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1635),
.B(n_1602),
.Y(n_1688)
);

OAI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1655),
.A2(n_1626),
.B1(n_1584),
.B2(n_1590),
.C(n_1621),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1640),
.B(n_1492),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1640),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1641),
.A2(n_1584),
.B1(n_1627),
.B2(n_1631),
.Y(n_1692)
);

AOI21x1_ASAP7_75t_L g1693 ( 
.A1(n_1658),
.A2(n_1603),
.B(n_1634),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1644),
.A2(n_1626),
.B1(n_1631),
.B2(n_1578),
.C(n_1592),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1637),
.B(n_1623),
.Y(n_1695)
);

NOR2x1_ASAP7_75t_L g1696 ( 
.A(n_1659),
.B(n_1583),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1660),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1637),
.B(n_1623),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1656),
.A2(n_1627),
.B1(n_1621),
.B2(n_1628),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1645),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1669),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1669),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1673),
.B(n_1643),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1693),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1696),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1700),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1673),
.B(n_1643),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1695),
.B(n_1654),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1683),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1681),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1685),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1681),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1687),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1667),
.B(n_1643),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1695),
.B(n_1654),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1698),
.B(n_1654),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1697),
.Y(n_1717)
);

OA21x2_ASAP7_75t_L g1718 ( 
.A1(n_1692),
.A2(n_1624),
.B(n_1620),
.Y(n_1718)
);

BUFx8_ASAP7_75t_L g1719 ( 
.A(n_1664),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1683),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1667),
.B(n_1645),
.Y(n_1721)
);

NAND3xp33_ASAP7_75t_L g1722 ( 
.A(n_1661),
.B(n_1627),
.C(n_1656),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1675),
.B(n_1645),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1672),
.Y(n_1724)
);

OA21x2_ASAP7_75t_L g1725 ( 
.A1(n_1694),
.A2(n_1624),
.B(n_1620),
.Y(n_1725)
);

NOR2x1p5_ASAP7_75t_L g1726 ( 
.A(n_1661),
.B(n_1638),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1717),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1717),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1713),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1710),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1708),
.B(n_1677),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1726),
.A2(n_1663),
.B1(n_1678),
.B2(n_1671),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1726),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1710),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1701),
.Y(n_1735)
);

INVx4_ASAP7_75t_L g1736 ( 
.A(n_1705),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_L g1737 ( 
.A(n_1722),
.B(n_1663),
.C(n_1678),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1701),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1717),
.B(n_1696),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1717),
.B(n_1666),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1701),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1710),
.B(n_1666),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1721),
.B(n_1675),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1703),
.B(n_1665),
.Y(n_1744)
);

NAND4xp75_ASAP7_75t_L g1745 ( 
.A(n_1725),
.B(n_1680),
.C(n_1676),
.D(n_1682),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1705),
.B(n_1666),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1708),
.B(n_1677),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1713),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1708),
.B(n_1668),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1703),
.B(n_1665),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1702),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1702),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1715),
.B(n_1668),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1715),
.B(n_1670),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1702),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1706),
.Y(n_1756)
);

NAND4xp25_ASAP7_75t_L g1757 ( 
.A(n_1722),
.B(n_1674),
.C(n_1699),
.D(n_1689),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1707),
.B(n_1690),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1721),
.B(n_1691),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1721),
.B(n_1688),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1724),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1706),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1715),
.B(n_1716),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_R g1764 ( 
.A(n_1719),
.B(n_1608),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1705),
.B(n_1638),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1709),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1709),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1707),
.B(n_1686),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1709),
.Y(n_1769)
);

OAI211xp5_ASAP7_75t_L g1770 ( 
.A1(n_1725),
.A2(n_1699),
.B(n_1684),
.C(n_1662),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1735),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1731),
.B(n_1716),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1731),
.B(n_1712),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1735),
.Y(n_1774)
);

AOI21xp33_ASAP7_75t_SL g1775 ( 
.A1(n_1737),
.A2(n_1732),
.B(n_1733),
.Y(n_1775)
);

AOI21xp33_ASAP7_75t_SL g1776 ( 
.A1(n_1744),
.A2(n_1725),
.B(n_1718),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1738),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1738),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1758),
.B(n_1719),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1763),
.Y(n_1780)
);

INVx2_ASAP7_75t_SL g1781 ( 
.A(n_1727),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1741),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1728),
.B(n_1712),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1750),
.B(n_1719),
.Y(n_1784)
);

INVxp33_ASAP7_75t_L g1785 ( 
.A(n_1764),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1745),
.B(n_1719),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1756),
.B(n_1723),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1741),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1763),
.Y(n_1789)
);

O2A1O1Ixp33_ASAP7_75t_L g1790 ( 
.A1(n_1757),
.A2(n_1711),
.B(n_1679),
.C(n_1725),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1751),
.Y(n_1791)
);

OR2x6_ASAP7_75t_L g1792 ( 
.A(n_1745),
.B(n_1514),
.Y(n_1792)
);

O2A1O1Ixp5_ASAP7_75t_L g1793 ( 
.A1(n_1770),
.A2(n_1711),
.B(n_1714),
.C(n_1723),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1729),
.B(n_1719),
.C(n_1718),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1748),
.B(n_1719),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1747),
.B(n_1723),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1747),
.B(n_1714),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1762),
.B(n_1686),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1742),
.B(n_1697),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1740),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1727),
.Y(n_1801)
);

NAND3xp33_ASAP7_75t_L g1802 ( 
.A(n_1736),
.B(n_1718),
.C(n_1725),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1742),
.B(n_1749),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1751),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1768),
.B(n_1640),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1752),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1728),
.B(n_1720),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1752),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1727),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1800),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1771),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1775),
.B(n_1749),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1771),
.Y(n_1813)
);

BUFx4f_ASAP7_75t_SL g1814 ( 
.A(n_1783),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1783),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1803),
.B(n_1740),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1774),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1807),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1785),
.B(n_1740),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1774),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1777),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1773),
.B(n_1753),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1777),
.Y(n_1823)
);

CKINVDCx14_ASAP7_75t_R g1824 ( 
.A(n_1792),
.Y(n_1824)
);

CKINVDCx16_ASAP7_75t_R g1825 ( 
.A(n_1792),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1778),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1778),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1803),
.B(n_1742),
.Y(n_1828)
);

INVx1_ASAP7_75t_SL g1829 ( 
.A(n_1773),
.Y(n_1829)
);

INVx4_ASAP7_75t_L g1830 ( 
.A(n_1783),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1782),
.Y(n_1831)
);

INVx1_ASAP7_75t_SL g1832 ( 
.A(n_1787),
.Y(n_1832)
);

AOI222xp33_ASAP7_75t_L g1833 ( 
.A1(n_1786),
.A2(n_1736),
.B1(n_1739),
.B2(n_1746),
.C1(n_1765),
.C2(n_1605),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1772),
.B(n_1753),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1782),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1788),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1788),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1807),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1828),
.B(n_1772),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1825),
.A2(n_1792),
.B1(n_1794),
.B2(n_1795),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1824),
.A2(n_1792),
.B1(n_1779),
.B2(n_1784),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1818),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1824),
.A2(n_1793),
.B(n_1790),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1829),
.B(n_1796),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1813),
.Y(n_1845)
);

NOR2xp67_ASAP7_75t_SL g1846 ( 
.A(n_1815),
.B(n_1736),
.Y(n_1846)
);

OAI222xp33_ASAP7_75t_L g1847 ( 
.A1(n_1812),
.A2(n_1814),
.B1(n_1832),
.B2(n_1810),
.C1(n_1830),
.C2(n_1815),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1819),
.B(n_1797),
.Y(n_1848)
);

AOI221xp5_ASAP7_75t_L g1849 ( 
.A1(n_1822),
.A2(n_1776),
.B1(n_1802),
.B2(n_1789),
.C(n_1780),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1813),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1817),
.Y(n_1851)
);

AO22x1_ASAP7_75t_L g1852 ( 
.A1(n_1815),
.A2(n_1739),
.B1(n_1781),
.B2(n_1801),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1817),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1816),
.A2(n_1789),
.B1(n_1780),
.B2(n_1796),
.Y(n_1854)
);

NOR3xp33_ASAP7_75t_L g1855 ( 
.A(n_1830),
.B(n_1781),
.C(n_1801),
.Y(n_1855)
);

AOI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1816),
.A2(n_1799),
.B1(n_1746),
.B2(n_1797),
.Y(n_1856)
);

A2O1A1Ixp33_ASAP7_75t_L g1857 ( 
.A1(n_1828),
.A2(n_1739),
.B(n_1787),
.C(n_1746),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1830),
.B(n_1834),
.Y(n_1858)
);

AOI21xp33_ASAP7_75t_SL g1859 ( 
.A1(n_1833),
.A2(n_1809),
.B(n_1798),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1835),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1839),
.B(n_1856),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1848),
.B(n_1838),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1842),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1842),
.B(n_1838),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1855),
.B(n_1838),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1858),
.B(n_1811),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1854),
.B(n_1799),
.Y(n_1867)
);

INVx1_ASAP7_75t_SL g1868 ( 
.A(n_1844),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1845),
.Y(n_1869)
);

INVx1_ASAP7_75t_SL g1870 ( 
.A(n_1852),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1850),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1859),
.B(n_1820),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1843),
.B(n_1809),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1864),
.Y(n_1874)
);

AOI221xp5_ASAP7_75t_L g1875 ( 
.A1(n_1872),
.A2(n_1847),
.B1(n_1849),
.B2(n_1841),
.C(n_1840),
.Y(n_1875)
);

A2O1A1Ixp33_ASAP7_75t_L g1876 ( 
.A1(n_1870),
.A2(n_1857),
.B(n_1846),
.C(n_1847),
.Y(n_1876)
);

AOI211xp5_ASAP7_75t_SL g1877 ( 
.A1(n_1865),
.A2(n_1860),
.B(n_1853),
.C(n_1851),
.Y(n_1877)
);

NAND3xp33_ASAP7_75t_L g1878 ( 
.A(n_1873),
.B(n_1823),
.C(n_1821),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1873),
.A2(n_1861),
.B1(n_1867),
.B2(n_1868),
.Y(n_1879)
);

NOR3xp33_ASAP7_75t_L g1880 ( 
.A(n_1862),
.B(n_1827),
.C(n_1826),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1861),
.A2(n_1863),
.B(n_1866),
.Y(n_1881)
);

O2A1O1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1869),
.A2(n_1831),
.B(n_1836),
.C(n_1835),
.Y(n_1882)
);

NAND4xp25_ASAP7_75t_L g1883 ( 
.A(n_1867),
.B(n_1871),
.C(n_1837),
.D(n_1836),
.Y(n_1883)
);

XOR2xp5_ASAP7_75t_L g1884 ( 
.A(n_1861),
.B(n_1837),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1874),
.B(n_1730),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1875),
.A2(n_1807),
.B1(n_1734),
.B2(n_1730),
.Y(n_1886)
);

O2A1O1Ixp5_ASAP7_75t_L g1887 ( 
.A1(n_1876),
.A2(n_1808),
.B(n_1806),
.C(n_1804),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1879),
.A2(n_1806),
.B1(n_1791),
.B2(n_1804),
.Y(n_1888)
);

A2O1A1Ixp33_ASAP7_75t_L g1889 ( 
.A1(n_1881),
.A2(n_1734),
.B(n_1765),
.C(n_1791),
.Y(n_1889)
);

AOI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1878),
.A2(n_1808),
.B1(n_1765),
.B2(n_1805),
.C(n_1767),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1884),
.A2(n_1759),
.B1(n_1743),
.B2(n_1760),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1887),
.Y(n_1892)
);

INVxp67_ASAP7_75t_SL g1893 ( 
.A(n_1885),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1886),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1891),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1889),
.B(n_1877),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1888),
.B(n_1883),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1890),
.B(n_1880),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1886),
.Y(n_1899)
);

BUFx3_ASAP7_75t_L g1900 ( 
.A(n_1895),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1893),
.Y(n_1901)
);

NOR2x1p5_ASAP7_75t_L g1902 ( 
.A(n_1896),
.B(n_1882),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1894),
.Y(n_1903)
);

NOR3xp33_ASAP7_75t_L g1904 ( 
.A(n_1897),
.B(n_1483),
.C(n_1759),
.Y(n_1904)
);

INVx3_ASAP7_75t_SL g1905 ( 
.A(n_1899),
.Y(n_1905)
);

NOR3x1_ASAP7_75t_L g1906 ( 
.A(n_1903),
.B(n_1898),
.C(n_1901),
.Y(n_1906)
);

NOR3xp33_ASAP7_75t_L g1907 ( 
.A(n_1900),
.B(n_1894),
.C(n_1892),
.Y(n_1907)
);

NOR3xp33_ASAP7_75t_L g1908 ( 
.A(n_1904),
.B(n_1743),
.C(n_1755),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1902),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1907),
.B(n_1902),
.Y(n_1910)
);

INVxp33_ASAP7_75t_SL g1911 ( 
.A(n_1906),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1910),
.B(n_1905),
.Y(n_1912)
);

AOI221xp5_ASAP7_75t_L g1913 ( 
.A1(n_1911),
.A2(n_1909),
.B1(n_1908),
.B2(n_1769),
.C(n_1755),
.Y(n_1913)
);

XNOR2xp5_ASAP7_75t_L g1914 ( 
.A(n_1912),
.B(n_1554),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1913),
.Y(n_1915)
);

AO21x2_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1914),
.B(n_1767),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1915),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_1917),
.Y(n_1918)
);

BUFx2_ASAP7_75t_L g1919 ( 
.A(n_1916),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1919),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1920),
.A2(n_1918),
.B1(n_1916),
.B2(n_1769),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1921),
.B(n_1761),
.Y(n_1922)
);

OAI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1922),
.A2(n_1760),
.B1(n_1761),
.B2(n_1766),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1923),
.A2(n_1766),
.B1(n_1761),
.B2(n_1754),
.Y(n_1924)
);

AOI211xp5_ASAP7_75t_L g1925 ( 
.A1(n_1924),
.A2(n_1540),
.B(n_1561),
.C(n_1704),
.Y(n_1925)
);


endmodule