module fake_jpeg_21623_n_297 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_17),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_45),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_41),
.B1(n_50),
.B2(n_17),
.Y(n_52)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_51),
.Y(n_69)
);

NAND2x1_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_2),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_30),
.Y(n_66)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_16),
.B1(n_45),
.B2(n_38),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_54),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_62),
.B(n_67),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_36),
.B1(n_20),
.B2(n_24),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_54),
.B1(n_49),
.B2(n_53),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_30),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_95),
.B1(n_102),
.B2(n_40),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_71),
.A2(n_93),
.B1(n_99),
.B2(n_100),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_29),
.B(n_23),
.C(n_27),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_98),
.A3(n_32),
.B1(n_35),
.B2(n_22),
.Y(n_113)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_74),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_76),
.A2(n_90),
.B1(n_101),
.B2(n_103),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_81),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_36),
.B1(n_51),
.B2(n_25),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_80),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_85),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_36),
.B1(n_51),
.B2(n_19),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_88),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_43),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_92),
.Y(n_118)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_42),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_19),
.B1(n_24),
.B2(n_28),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_60),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_94),
.B(n_104),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_40),
.B1(n_67),
.B2(n_62),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_96),
.Y(n_134)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_23),
.B(n_18),
.C(n_27),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_56),
.A2(n_59),
.B1(n_63),
.B2(n_42),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_28),
.B1(n_29),
.B2(n_18),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_39),
.B1(n_37),
.B2(n_35),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_60),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_34),
.B1(n_31),
.B2(n_26),
.Y(n_123)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_106),
.B(n_108),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_30),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_30),
.C(n_39),
.Y(n_109)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_108),
.C(n_80),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_125),
.B1(n_132),
.B2(n_87),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_113),
.B(n_121),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_78),
.A2(n_37),
.B(n_22),
.C(n_31),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_129),
.B(n_10),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_34),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_127),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_75),
.A2(n_34),
.B1(n_31),
.B2(n_26),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_3),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_3),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_8),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_84),
.A2(n_99),
.B(n_95),
.C(n_102),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_89),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_88),
.A2(n_4),
.B(n_6),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_98),
.B(n_72),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_146),
.B(n_152),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_70),
.B1(n_77),
.B2(n_95),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_154),
.B1(n_157),
.B2(n_121),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_88),
.B1(n_87),
.B2(n_95),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_140),
.A2(n_139),
.B1(n_115),
.B2(n_146),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_97),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_143),
.Y(n_167)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_76),
.B1(n_90),
.B2(n_85),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

AND2x4_ASAP7_75t_SL g146 ( 
.A(n_113),
.B(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_133),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_130),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_161),
.Y(n_164)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_96),
.B1(n_91),
.B2(n_73),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_155),
.B(n_118),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_9),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_158),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_105),
.B1(n_10),
.B2(n_11),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_9),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_9),
.B(n_10),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_118),
.B(n_132),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_155),
.B1(n_157),
.B2(n_159),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_130),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_117),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_160),
.A2(n_122),
.B(n_112),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_163),
.A2(n_169),
.B(n_190),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_166),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_112),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_168),
.B(n_185),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_120),
.B(n_111),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_174),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_127),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_174),
.B(n_142),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_120),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_119),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_179),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_181),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_119),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_137),
.B(n_156),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_134),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_154),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_152),
.A2(n_131),
.B1(n_125),
.B2(n_134),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

AOI22x1_ASAP7_75t_SL g190 ( 
.A1(n_138),
.A2(n_133),
.B1(n_116),
.B2(n_13),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_150),
.C(n_142),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_196),
.C(n_205),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_165),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_185),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_201),
.Y(n_228)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_177),
.Y(n_201)
);

OAI22x1_ASAP7_75t_SL g203 ( 
.A1(n_190),
.A2(n_140),
.B1(n_149),
.B2(n_139),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_166),
.B1(n_189),
.B2(n_171),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_150),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_173),
.B1(n_178),
.B2(n_190),
.Y(n_221)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_153),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_208),
.B(n_164),
.Y(n_225)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_176),
.C(n_167),
.Y(n_227)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_163),
.A2(n_147),
.B(n_158),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_183),
.B(n_164),
.Y(n_223)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_188),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_215),
.B(n_218),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_168),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_217),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_180),
.B1(n_163),
.B2(n_169),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_219),
.A2(n_197),
.B1(n_202),
.B2(n_213),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_209),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_220),
.B(n_212),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_191),
.C(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_223),
.A2(n_192),
.B1(n_204),
.B2(n_200),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_240),
.B1(n_241),
.B2(n_249),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_228),
.A2(n_204),
.B1(n_200),
.B2(n_193),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_228),
.A2(n_193),
.B1(n_203),
.B2(n_201),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_224),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_242),
.B(n_232),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_216),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_245),
.A2(n_222),
.B1(n_194),
.B2(n_230),
.Y(n_263)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_210),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_218),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g249 ( 
.A1(n_215),
.A2(n_214),
.B1(n_202),
.B2(n_182),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_260),
.C(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_226),
.B(n_216),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_261),
.B(n_264),
.Y(n_271)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_259),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_205),
.C(n_227),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_196),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_219),
.B(n_222),
.C(n_226),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_232),
.C(n_231),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_240),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_253),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_267),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_272),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_235),
.C(n_237),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_237),
.C(n_250),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_273),
.Y(n_277)
);

BUFx4f_ASAP7_75t_SL g274 ( 
.A(n_261),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_234),
.B(n_257),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_275),
.B(n_144),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_262),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_279),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_268),
.A2(n_238),
.B1(n_252),
.B2(n_261),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_231),
.B(n_230),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_280),
.A2(n_229),
.B(n_167),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g282 ( 
.A1(n_277),
.A2(n_269),
.A3(n_229),
.B1(n_271),
.B2(n_261),
.C1(n_274),
.C2(n_270),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_285),
.B(n_287),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_194),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_284),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_278),
.A2(n_241),
.B1(n_236),
.B2(n_222),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_287),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_293),
.C(n_187),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_276),
.C(n_187),
.Y(n_293)
);

O2A1O1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_291),
.B(n_288),
.C(n_143),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_182),
.B1(n_144),
.B2(n_211),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_11),
.B(n_12),
.Y(n_297)
);


endmodule