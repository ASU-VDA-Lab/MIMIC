module fake_aes_297_n_692 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_692);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_692;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_599;
wire n_305;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_529;
wire n_312;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_613;
wire n_247;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_415;
wire n_482;
wire n_235;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_285;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_62), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_58), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_41), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_67), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_9), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_69), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_36), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_30), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_25), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_74), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_1), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_20), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_1), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_22), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_23), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_33), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_21), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_64), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_15), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_52), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_61), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_71), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_55), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_59), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_12), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_31), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_35), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_60), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_46), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_57), .Y(n_106) );
INVxp33_ASAP7_75t_L g107 ( .A(n_51), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_6), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_9), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_72), .Y(n_110) );
INVx3_ASAP7_75t_L g111 ( .A(n_45), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_2), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_32), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_18), .Y(n_114) );
INVx2_ASAP7_75t_SL g115 ( .A(n_28), .Y(n_115) );
CKINVDCx14_ASAP7_75t_R g116 ( .A(n_26), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_63), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_24), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_19), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_29), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_66), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_44), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_75), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_12), .Y(n_124) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_85), .A2(n_0), .B(n_2), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_95), .A2(n_0), .B1(n_3), .B2(n_4), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_111), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_111), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_111), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_105), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_122), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_114), .B(n_3), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_105), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_115), .B(n_4), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_88), .Y(n_138) );
INVx1_ASAP7_75t_SL g139 ( .A(n_112), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_88), .Y(n_140) );
INVx1_ASAP7_75t_SL g141 ( .A(n_112), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_90), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_122), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_115), .B(n_5), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_90), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_87), .B(n_5), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_91), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_87), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_91), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_120), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_101), .B(n_6), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_120), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_107), .B(n_7), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_121), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_121), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_77), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_79), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_116), .B(n_7), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_80), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_101), .B(n_8), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_82), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_83), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_93), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_96), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_99), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_102), .Y(n_166) );
NOR3xp33_ASAP7_75t_L g167 ( .A(n_126), .B(n_89), .C(n_124), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_135), .A2(n_108), .B1(n_109), .B2(n_81), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_131), .Y(n_169) );
NOR3xp33_ASAP7_75t_L g170 ( .A(n_126), .B(n_84), .C(n_98), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_161), .B(n_123), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_153), .A2(n_95), .B1(n_78), .B2(n_104), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_128), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_139), .B(n_106), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_139), .B(n_106), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_151), .Y(n_176) );
BUFx10_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_127), .B(n_94), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_128), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_135), .A2(n_119), .B1(n_118), .B2(n_117), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_140), .A2(n_110), .B1(n_103), .B2(n_92), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_141), .B(n_113), .Y(n_182) );
INVxp67_ASAP7_75t_L g183 ( .A(n_141), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_127), .B(n_113), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_148), .A2(n_100), .B(n_97), .C(n_94), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_161), .B(n_100), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_144), .B(n_97), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_144), .B(n_42), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_127), .B(n_8), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_163), .B(n_43), .Y(n_191) );
NOR3xp33_ASAP7_75t_L g192 ( .A(n_134), .B(n_10), .C(n_11), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_153), .A2(n_10), .B1(n_11), .B2(n_13), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_127), .B(n_13), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_129), .B(n_14), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_144), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_158), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_151), .Y(n_198) );
INVx2_ASAP7_75t_SL g199 ( .A(n_158), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_151), .Y(n_200) );
INVxp33_ASAP7_75t_L g201 ( .A(n_148), .Y(n_201) );
AND2x6_ASAP7_75t_L g202 ( .A(n_144), .B(n_48), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_153), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_128), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_129), .B(n_16), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_129), .B(n_17), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_129), .B(n_27), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_137), .B(n_34), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_129), .B(n_37), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_128), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_163), .B(n_147), .Y(n_211) );
INVxp67_ASAP7_75t_L g212 ( .A(n_158), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_151), .A2(n_160), .B1(n_147), .B2(n_140), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_142), .B(n_38), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_160), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_142), .B(n_39), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_149), .B(n_40), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_137), .B(n_47), .Y(n_218) );
NOR2xp67_ASAP7_75t_L g219 ( .A(n_137), .B(n_49), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_149), .A2(n_50), .B(n_53), .C(n_54), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_138), .A2(n_56), .B(n_65), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_157), .B(n_68), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_137), .B(n_70), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_137), .B(n_73), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_157), .B(n_76), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_160), .A2(n_136), .B1(n_152), .B2(n_138), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_160), .B(n_145), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_160), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_201), .B(n_132), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_186), .B(n_145), .Y(n_230) );
OR2x6_ASAP7_75t_L g231 ( .A(n_199), .B(n_146), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_183), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_173), .Y(n_233) );
NOR2x1_ASAP7_75t_L g234 ( .A(n_175), .B(n_134), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_186), .B(n_145), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_187), .B(n_145), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_197), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_187), .B(n_145), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_227), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_174), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_179), .Y(n_241) );
INVx4_ASAP7_75t_L g242 ( .A(n_202), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_204), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_171), .B(n_211), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_171), .B(n_154), .Y(n_245) );
NOR2xp33_ASAP7_75t_R g246 ( .A(n_196), .B(n_157), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_210), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_227), .Y(n_248) );
BUFx4f_ASAP7_75t_SL g249 ( .A(n_182), .Y(n_249) );
AO221x1_ASAP7_75t_L g250 ( .A1(n_212), .A2(n_154), .B1(n_155), .B2(n_157), .C(n_162), .Y(n_250) );
CKINVDCx11_ASAP7_75t_R g251 ( .A(n_177), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_178), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_211), .B(n_154), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_226), .B(n_132), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_196), .A2(n_125), .B1(n_162), .B2(n_157), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_226), .B(n_146), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_184), .B(n_155), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_213), .B(n_180), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_167), .A2(n_152), .B(n_150), .C(n_138), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_176), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_180), .B(n_154), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_189), .B(n_162), .Y(n_262) );
BUFx4f_ASAP7_75t_SL g263 ( .A(n_202), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_170), .A2(n_162), .B1(n_154), .B2(n_155), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_198), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_202), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_200), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_177), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_215), .B(n_155), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_228), .B(n_155), .Y(n_270) );
AO22x1_ASAP7_75t_L g271 ( .A1(n_202), .A2(n_136), .B1(n_152), .B2(n_150), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_181), .B(n_162), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_181), .B(n_185), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_168), .B(n_166), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_195), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_168), .B(n_166), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_172), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_202), .A2(n_166), .B1(n_164), .B2(n_159), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_169), .Y(n_279) );
AO22x1_ASAP7_75t_L g280 ( .A1(n_192), .A2(n_136), .B1(n_150), .B2(n_164), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_188), .A2(n_164), .B1(n_159), .B2(n_125), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_169), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_224), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_188), .A2(n_136), .B(n_159), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_169), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_205), .Y(n_286) );
INVx2_ASAP7_75t_SL g287 ( .A(n_190), .Y(n_287) );
INVx4_ASAP7_75t_L g288 ( .A(n_169), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_194), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_191), .B(n_130), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_193), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_191), .B(n_130), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_222), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_219), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_248), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_239), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_256), .B(n_203), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_233), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_232), .B(n_125), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_256), .B(n_125), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_283), .A2(n_207), .B(n_206), .Y(n_301) );
BUFx4f_ASAP7_75t_L g302 ( .A(n_231), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_252), .B(n_125), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_232), .B(n_125), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_258), .A2(n_214), .B1(n_217), .B2(n_216), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_248), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_273), .B(n_209), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_239), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_293), .A2(n_208), .B(n_223), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_286), .B(n_130), .Y(n_310) );
CKINVDCx6p67_ASAP7_75t_R g311 ( .A(n_251), .Y(n_311) );
A2O1A1Ixp33_ASAP7_75t_L g312 ( .A1(n_259), .A2(n_133), .B(n_220), .C(n_221), .Y(n_312) );
NAND2xp33_ASAP7_75t_L g313 ( .A(n_246), .B(n_223), .Y(n_313) );
CKINVDCx12_ASAP7_75t_R g314 ( .A(n_231), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_254), .A2(n_165), .B1(n_156), .B2(n_133), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_244), .B(n_133), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_233), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_293), .A2(n_208), .B(n_218), .Y(n_318) );
INVx5_ASAP7_75t_L g319 ( .A(n_242), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_239), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_254), .B(n_156), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_263), .A2(n_156), .B1(n_165), .B2(n_218), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_241), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_275), .B(n_231), .Y(n_324) );
AND2x2_ASAP7_75t_SL g325 ( .A(n_242), .B(n_156), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_236), .Y(n_326) );
OAI21x1_ASAP7_75t_SL g327 ( .A1(n_242), .A2(n_225), .B(n_156), .Y(n_327) );
OAI21xp33_ASAP7_75t_L g328 ( .A1(n_277), .A2(n_156), .B(n_165), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_266), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_266), .B(n_156), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_231), .B(n_156), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_238), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_250), .A2(n_165), .B1(n_131), .B2(n_143), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_268), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_240), .B(n_165), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_240), .B(n_165), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_251), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_229), .B(n_165), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_269), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_268), .B(n_234), .Y(n_340) );
INVx4_ASAP7_75t_L g341 ( .A(n_237), .Y(n_341) );
A2O1A1Ixp33_ASAP7_75t_L g342 ( .A1(n_260), .A2(n_165), .B(n_131), .C(n_143), .Y(n_342) );
OR2x6_ASAP7_75t_L g343 ( .A(n_291), .B(n_131), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_257), .A2(n_131), .B(n_143), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_270), .A2(n_131), .B(n_143), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_297), .B(n_264), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_314), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_298), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_319), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_295), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_306), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_319), .Y(n_352) );
NAND2x1p5_ASAP7_75t_L g353 ( .A(n_319), .B(n_267), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_298), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_317), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_317), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_339), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_323), .Y(n_358) );
INVx8_ASAP7_75t_L g359 ( .A(n_319), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_323), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_308), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_326), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_302), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_309), .A2(n_284), .B(n_281), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_332), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_316), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_321), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_320), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_335), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_324), .B(n_265), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_296), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_296), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_336), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_329), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_329), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_329), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_310), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_346), .B(n_300), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_358), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_366), .B(n_302), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_358), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_348), .Y(n_382) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_377), .Y(n_383) );
BUFx4f_ASAP7_75t_L g384 ( .A(n_359), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_366), .B(n_260), .Y(n_385) );
INVx1_ASAP7_75t_SL g386 ( .A(n_348), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_360), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_363), .B(n_237), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_357), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_359), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_360), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_357), .Y(n_392) );
NOR2x1_ASAP7_75t_L g393 ( .A(n_352), .B(n_343), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_350), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_350), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_354), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_355), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_377), .B(n_299), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_367), .B(n_265), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_351), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_355), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_362), .B(n_334), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_362), .B(n_334), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_359), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_379), .B(n_356), .Y(n_406) );
OAI21x1_ASAP7_75t_L g407 ( .A1(n_393), .A2(n_364), .B(n_344), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_383), .Y(n_408) );
BUFx3_ASAP7_75t_L g409 ( .A(n_384), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_382), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_384), .Y(n_411) );
INVx4_ASAP7_75t_L g412 ( .A(n_384), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_382), .Y(n_413) );
AOI222xp33_ASAP7_75t_L g414 ( .A1(n_384), .A2(n_365), .B1(n_363), .B2(n_337), .C1(n_351), .C2(n_341), .Y(n_414) );
AOI22xp33_ASAP7_75t_SL g415 ( .A1(n_380), .A2(n_341), .B1(n_337), .B2(n_250), .Y(n_415) );
OR2x6_ASAP7_75t_L g416 ( .A(n_390), .B(n_359), .Y(n_416) );
AOI211xp5_ASAP7_75t_L g417 ( .A1(n_380), .A2(n_388), .B(n_405), .C(n_390), .Y(n_417) );
NAND4xp25_ASAP7_75t_L g418 ( .A(n_395), .B(n_338), .C(n_365), .D(n_304), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_379), .B(n_369), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_405), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_382), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_394), .Y(n_422) );
OA21x2_ASAP7_75t_L g423 ( .A1(n_395), .A2(n_364), .B(n_342), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_399), .A2(n_367), .B1(n_333), .B2(n_370), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_394), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_390), .A2(n_373), .B1(n_369), .B2(n_347), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_405), .A2(n_373), .B1(n_338), .B2(n_340), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_386), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g429 ( .A1(n_385), .A2(n_359), .B(n_307), .C(n_278), .Y(n_429) );
INVx4_ASAP7_75t_L g430 ( .A(n_394), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_381), .B(n_376), .Y(n_431) );
OAI21x1_ASAP7_75t_L g432 ( .A1(n_393), .A2(n_345), .B(n_327), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_396), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_397), .Y(n_434) );
BUFx5_ASAP7_75t_L g435 ( .A(n_381), .Y(n_435) );
OA222x2_ASAP7_75t_L g436 ( .A1(n_396), .A2(n_343), .B1(n_352), .B2(n_303), .C1(n_356), .C2(n_361), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_397), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_389), .A2(n_280), .B1(n_245), .B2(n_368), .C(n_340), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_385), .A2(n_333), .B1(n_343), .B2(n_353), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_401), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_408), .B(n_392), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_430), .B(n_401), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_440), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_435), .Y(n_444) );
NAND4xp25_ASAP7_75t_L g445 ( .A(n_417), .B(n_315), .C(n_294), .D(n_403), .Y(n_445) );
NOR2x1_ASAP7_75t_SL g446 ( .A(n_416), .B(n_337), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_410), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_433), .B(n_387), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_440), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_408), .B(n_387), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_433), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_410), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_420), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_419), .B(n_391), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_428), .B(n_391), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_413), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_417), .B(n_386), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_413), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_419), .B(n_404), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_406), .B(n_402), .Y(n_460) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_428), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_418), .B(n_398), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_418), .B(n_398), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_406), .B(n_402), .Y(n_464) );
AOI211x1_ASAP7_75t_L g465 ( .A1(n_439), .A2(n_280), .B(n_403), .C(n_404), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_421), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_435), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_435), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_435), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_430), .B(n_402), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_426), .B(n_378), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_435), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_430), .B(n_398), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_420), .B(n_378), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_430), .B(n_397), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_435), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_427), .B(n_400), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_421), .B(n_368), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_435), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_435), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_422), .B(n_400), .Y(n_481) );
NOR2xp67_ASAP7_75t_SL g482 ( .A(n_409), .B(n_337), .Y(n_482) );
OAI22xp33_ASAP7_75t_L g483 ( .A1(n_412), .A2(n_311), .B1(n_353), .B2(n_352), .Y(n_483) );
NOR2xp67_ASAP7_75t_L g484 ( .A(n_412), .B(n_349), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_422), .B(n_361), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_425), .B(n_375), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_425), .B(n_315), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_434), .B(n_375), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_434), .B(n_376), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_435), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_437), .Y(n_491) );
NOR2x1_ASAP7_75t_L g492 ( .A(n_483), .B(n_412), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_441), .B(n_437), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_443), .Y(n_494) );
AND2x2_ASAP7_75t_SL g495 ( .A(n_442), .B(n_412), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_441), .B(n_431), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_459), .B(n_431), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_460), .B(n_431), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_460), .B(n_431), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_449), .Y(n_500) );
INVxp33_ASAP7_75t_L g501 ( .A(n_446), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_464), .B(n_436), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_464), .B(n_436), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_470), .Y(n_504) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_444), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_450), .B(n_416), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_451), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_485), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_481), .B(n_442), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_454), .B(n_423), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_450), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_453), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_465), .B(n_415), .C(n_414), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_455), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_445), .B(n_429), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_455), .Y(n_516) );
NAND2xp33_ASAP7_75t_L g517 ( .A(n_444), .B(n_411), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_477), .A2(n_416), .B1(n_409), .B2(n_411), .Y(n_518) );
NAND3xp33_ASAP7_75t_L g519 ( .A(n_482), .B(n_438), .C(n_143), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_481), .B(n_423), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_448), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_478), .Y(n_522) );
NOR2xp33_ASAP7_75t_SL g523 ( .A(n_482), .B(n_409), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_485), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_447), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_447), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_490), .B(n_411), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_478), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_461), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_442), .B(n_416), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_474), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_471), .B(n_423), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_491), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_470), .B(n_423), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_473), .B(n_416), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_473), .B(n_424), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_462), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_462), .B(n_411), .Y(n_538) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_484), .B(n_349), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_490), .B(n_407), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_475), .Y(n_541) );
INVxp67_ASAP7_75t_L g542 ( .A(n_457), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_463), .A2(n_407), .B1(n_372), .B2(n_371), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_452), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_475), .B(n_432), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_463), .B(n_294), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_452), .B(n_432), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_456), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_456), .B(n_331), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_458), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_531), .B(n_457), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_509), .B(n_476), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_511), .B(n_458), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_504), .B(n_466), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_514), .B(n_466), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_494), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_495), .B(n_479), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_500), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_507), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_516), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_533), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_521), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_512), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_515), .B(n_480), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_522), .B(n_486), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_528), .B(n_486), .Y(n_566) );
O2A1O1Ixp5_ASAP7_75t_L g567 ( .A1(n_501), .A2(n_468), .B(n_469), .C(n_472), .Y(n_567) );
AOI21xp5_ASAP7_75t_SL g568 ( .A1(n_515), .A2(n_467), .B(n_487), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_498), .B(n_489), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_508), .B(n_488), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_541), .B(n_489), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_493), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_537), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_524), .B(n_488), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_529), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_497), .B(n_487), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_546), .B(n_131), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_529), .Y(n_578) );
NAND2xp33_ASAP7_75t_L g579 ( .A(n_492), .B(n_349), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_548), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_548), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_546), .B(n_131), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_495), .B(n_349), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_525), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_499), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_550), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_496), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_502), .B(n_143), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_513), .A2(n_372), .B1(n_371), .B2(n_331), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_506), .Y(n_590) );
OAI22xp33_ASAP7_75t_L g591 ( .A1(n_501), .A2(n_353), .B1(n_349), .B2(n_249), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_526), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_544), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_503), .B(n_143), .Y(n_594) );
INVx4_ASAP7_75t_L g595 ( .A(n_539), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_538), .B(n_143), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_538), .B(n_532), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_510), .B(n_542), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_542), .B(n_342), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_547), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_520), .B(n_328), .Y(n_601) );
INVxp67_ASAP7_75t_SL g602 ( .A(n_505), .Y(n_602) );
AOI21xp33_ASAP7_75t_L g603 ( .A1(n_564), .A2(n_512), .B(n_518), .Y(n_603) );
NOR3xp33_ASAP7_75t_L g604 ( .A(n_588), .B(n_519), .C(n_527), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_556), .Y(n_605) );
NAND4xp25_ASAP7_75t_L g606 ( .A(n_564), .B(n_543), .C(n_530), .D(n_545), .Y(n_606) );
NOR2x1_ASAP7_75t_L g607 ( .A(n_579), .B(n_517), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_563), .B(n_535), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_552), .B(n_505), .Y(n_609) );
OAI21xp33_ASAP7_75t_L g610 ( .A1(n_568), .A2(n_598), .B(n_597), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_571), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_562), .B(n_527), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_591), .B(n_505), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_558), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_559), .Y(n_615) );
NOR2x1_ASAP7_75t_L g616 ( .A(n_579), .B(n_517), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_561), .Y(n_617) );
NAND4xp25_ASAP7_75t_L g618 ( .A(n_589), .B(n_543), .C(n_536), .D(n_523), .Y(n_618) );
AND4x1_ASAP7_75t_L g619 ( .A(n_568), .B(n_534), .C(n_255), .D(n_312), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_583), .A2(n_539), .B(n_540), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_575), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_578), .Y(n_622) );
NAND3xp33_ASAP7_75t_SL g623 ( .A(n_583), .B(n_549), .C(n_312), .Y(n_623) );
INVxp67_ASAP7_75t_SL g624 ( .A(n_581), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_591), .A2(n_505), .B(n_540), .C(n_271), .Y(n_625) );
AOI21xp33_ASAP7_75t_L g626 ( .A1(n_594), .A2(n_292), .B(n_290), .Y(n_626) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_595), .B(n_376), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_573), .B(n_307), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_560), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_554), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_557), .A2(n_271), .B(n_313), .Y(n_631) );
NAND3xp33_ASAP7_75t_L g632 ( .A(n_567), .B(n_374), .C(n_318), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_572), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_585), .B(n_374), .Y(n_634) );
NAND4xp25_ASAP7_75t_SL g635 ( .A(n_589), .B(n_274), .C(n_276), .D(n_261), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_569), .B(n_374), .Y(n_636) );
NAND4xp75_ASAP7_75t_L g637 ( .A(n_557), .B(n_325), .C(n_330), .D(n_289), .Y(n_637) );
OAI21xp5_ASAP7_75t_L g638 ( .A1(n_577), .A2(n_325), .B(n_287), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_607), .A2(n_595), .B1(n_587), .B2(n_590), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_616), .A2(n_595), .B1(n_566), .B2(n_565), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_625), .A2(n_602), .B1(n_576), .B2(n_551), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_611), .B(n_580), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_630), .B(n_574), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_603), .A2(n_582), .B1(n_596), .B2(n_599), .C(n_555), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g645 ( .A1(n_610), .A2(n_553), .B1(n_586), .B2(n_600), .C(n_570), .Y(n_645) );
INVxp67_ASAP7_75t_SL g646 ( .A(n_624), .Y(n_646) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_624), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_606), .A2(n_600), .B1(n_581), .B2(n_592), .C(n_593), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_605), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_614), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_618), .A2(n_593), .B1(n_584), .B2(n_601), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_620), .B(n_584), .Y(n_652) );
NAND4xp75_ASAP7_75t_L g653 ( .A(n_613), .B(n_289), .C(n_330), .D(n_272), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_633), .B(n_287), .Y(n_654) );
INVx2_ASAP7_75t_SL g655 ( .A(n_609), .Y(n_655) );
INVxp67_ASAP7_75t_L g656 ( .A(n_612), .Y(n_656) );
AOI221xp5_ASAP7_75t_SL g657 ( .A1(n_608), .A2(n_322), .B1(n_305), .B2(n_230), .C(n_235), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_615), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_617), .Y(n_659) );
O2A1O1Ixp5_ASAP7_75t_L g660 ( .A1(n_612), .A2(n_301), .B(n_253), .C(n_288), .Y(n_660) );
AND4x2_ASAP7_75t_L g661 ( .A(n_644), .B(n_627), .C(n_631), .D(n_619), .Y(n_661) );
NOR3x1_ASAP7_75t_L g662 ( .A(n_639), .B(n_637), .C(n_621), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_651), .B(n_628), .C(n_604), .D(n_626), .Y(n_663) );
OA21x2_ASAP7_75t_L g664 ( .A1(n_646), .A2(n_622), .B(n_629), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_649), .Y(n_665) );
AOI221xp5_ASAP7_75t_SL g666 ( .A1(n_656), .A2(n_634), .B1(n_636), .B2(n_638), .C(n_635), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_650), .Y(n_667) );
OAI211xp5_ASAP7_75t_L g668 ( .A1(n_656), .A2(n_604), .B(n_634), .C(n_623), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_647), .Y(n_669) );
XNOR2x1_ASAP7_75t_L g670 ( .A(n_640), .B(n_632), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_641), .B(n_288), .C(n_262), .Y(n_671) );
NOR3xp33_ASAP7_75t_L g672 ( .A(n_645), .B(n_288), .C(n_267), .Y(n_672) );
A2O1A1Ixp33_ASAP7_75t_L g673 ( .A1(n_646), .A2(n_329), .B(n_243), .C(n_247), .Y(n_673) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_664), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_666), .A2(n_648), .B1(n_652), .B2(n_642), .Y(n_675) );
AO22x2_ASAP7_75t_L g676 ( .A1(n_670), .A2(n_669), .B1(n_665), .B2(n_667), .Y(n_676) );
OAI22xp5_ASAP7_75t_SL g677 ( .A1(n_664), .A2(n_654), .B1(n_655), .B2(n_643), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_663), .A2(n_659), .B1(n_658), .B2(n_657), .C(n_660), .Y(n_678) );
AOI222xp33_ASAP7_75t_L g679 ( .A1(n_668), .A2(n_653), .B1(n_660), .B2(n_247), .C1(n_241), .C2(n_243), .Y(n_679) );
INVx3_ASAP7_75t_L g680 ( .A(n_662), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_663), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_681), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_680), .A2(n_666), .B1(n_671), .B2(n_672), .C(n_673), .Y(n_683) );
OR4x2_ASAP7_75t_L g684 ( .A(n_677), .B(n_661), .C(n_282), .D(n_285), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_678), .B(n_285), .Y(n_685) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_682), .A2(n_675), .B(n_674), .C(n_679), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_685), .B(n_676), .C(n_279), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_683), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_686), .A2(n_676), .B(n_684), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_688), .A2(n_279), .B(n_282), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_690), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_691), .A2(n_689), .B(n_687), .Y(n_692) );
endmodule