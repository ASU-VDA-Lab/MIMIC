module real_aes_2588_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_0), .B(n_131), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_1), .A2(n_140), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_2), .B(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_3), .B(n_131), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_4), .B(n_147), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_5), .B(n_147), .Y(n_523) );
INVx1_ASAP7_75t_L g138 ( .A(n_6), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_7), .B(n_147), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_8), .Y(n_116) );
NAND2xp33_ASAP7_75t_L g544 ( .A(n_9), .B(n_149), .Y(n_544) );
AND2x2_ASAP7_75t_L g167 ( .A(n_10), .B(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g244 ( .A(n_11), .B(n_156), .Y(n_244) );
INVx2_ASAP7_75t_L g153 ( .A(n_12), .Y(n_153) );
AOI221x1_ASAP7_75t_L g568 ( .A1(n_13), .A2(n_26), .B1(n_131), .B2(n_140), .C(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_14), .B(n_147), .Y(n_225) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_15), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_16), .B(n_131), .Y(n_540) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_17), .A2(n_156), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_18), .B(n_151), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_19), .B(n_147), .Y(n_500) );
AO21x1_ASAP7_75t_L g518 ( .A1(n_20), .A2(n_131), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_21), .B(n_131), .Y(n_198) );
INVx1_ASAP7_75t_L g113 ( .A(n_22), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_23), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_24), .A2(n_86), .B1(n_131), .B2(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g474 ( .A(n_25), .Y(n_474) );
NAND2xp33_ASAP7_75t_R g778 ( .A(n_25), .B(n_779), .Y(n_778) );
NAND2x1_ASAP7_75t_L g561 ( .A(n_27), .B(n_147), .Y(n_561) );
NAND2x1_ASAP7_75t_L g510 ( .A(n_28), .B(n_149), .Y(n_510) );
OR2x2_ASAP7_75t_L g154 ( .A(n_29), .B(n_83), .Y(n_154) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_29), .A2(n_83), .B(n_153), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_30), .B(n_149), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_31), .B(n_147), .Y(n_543) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_32), .A2(n_168), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_33), .B(n_149), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_34), .A2(n_140), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_35), .B(n_147), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_36), .A2(n_140), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g137 ( .A(n_37), .B(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g141 ( .A(n_37), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g181 ( .A(n_37), .Y(n_181) );
OR2x6_ASAP7_75t_L g111 ( .A(n_38), .B(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_39), .B(n_131), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_40), .B(n_131), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_41), .B(n_147), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_42), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_43), .B(n_149), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_44), .B(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_45), .A2(n_140), .B(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_46), .A2(n_140), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_47), .B(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_48), .B(n_149), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_49), .B(n_131), .Y(n_222) );
INVx1_ASAP7_75t_L g134 ( .A(n_50), .Y(n_134) );
INVx1_ASAP7_75t_L g144 ( .A(n_50), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_51), .B(n_147), .Y(n_165) );
AOI221xp5_ASAP7_75t_L g98 ( .A1(n_52), .A2(n_99), .B1(n_117), .B2(n_467), .C(n_472), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_52), .A2(n_120), .B1(n_462), .B2(n_463), .Y(n_119) );
INVx1_ASAP7_75t_L g462 ( .A(n_52), .Y(n_462) );
AND2x2_ASAP7_75t_L g188 ( .A(n_53), .B(n_151), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_54), .B(n_149), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_55), .B(n_147), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_56), .B(n_149), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_57), .A2(n_140), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_58), .B(n_131), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_59), .B(n_131), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_60), .A2(n_140), .B(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g204 ( .A(n_61), .B(n_152), .Y(n_204) );
AO21x1_ASAP7_75t_L g520 ( .A1(n_62), .A2(n_140), .B(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_63), .B(n_131), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_64), .B(n_149), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_65), .B(n_131), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_66), .B(n_149), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_67), .A2(n_90), .B1(n_140), .B2(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_68), .B(n_147), .Y(n_201) );
AND2x2_ASAP7_75t_L g534 ( .A(n_69), .B(n_152), .Y(n_534) );
INVx1_ASAP7_75t_L g136 ( .A(n_70), .Y(n_136) );
INVx1_ASAP7_75t_L g142 ( .A(n_70), .Y(n_142) );
AND2x2_ASAP7_75t_L g513 ( .A(n_71), .B(n_168), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_72), .B(n_149), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_73), .A2(n_140), .B(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_74), .A2(n_140), .B(n_145), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_75), .A2(n_140), .B(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g216 ( .A(n_76), .B(n_152), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_77), .B(n_151), .Y(n_170) );
INVx1_ASAP7_75t_L g114 ( .A(n_78), .Y(n_114) );
AND2x2_ASAP7_75t_L g486 ( .A(n_79), .B(n_168), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_80), .B(n_131), .Y(n_502) );
AND2x2_ASAP7_75t_L g155 ( .A(n_81), .B(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g519 ( .A(n_82), .B(n_195), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_84), .B(n_149), .Y(n_501) );
AND2x2_ASAP7_75t_L g564 ( .A(n_85), .B(n_168), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_87), .B(n_147), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_88), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_89), .A2(n_140), .B(n_499), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_91), .A2(n_140), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_92), .B(n_149), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_93), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_94), .B(n_147), .Y(n_491) );
BUFx2_ASAP7_75t_L g203 ( .A(n_95), .Y(n_203) );
BUFx2_ASAP7_75t_SL g105 ( .A(n_96), .Y(n_105) );
BUFx2_ASAP7_75t_L g471 ( .A(n_96), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_97), .A2(n_140), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_SL g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_106), .B(n_115), .Y(n_102) );
CKINVDCx11_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx8_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_R g464 ( .A(n_108), .Y(n_464) );
BUFx2_ASAP7_75t_L g792 ( .A(n_108), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x6_ASAP7_75t_SL g477 ( .A(n_109), .B(n_111), .Y(n_477) );
OR2x6_ASAP7_75t_SL g777 ( .A(n_109), .B(n_110), .Y(n_777) );
OR2x2_ASAP7_75t_L g786 ( .A(n_109), .B(n_111), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OR2x2_ASAP7_75t_SL g470 ( .A(n_115), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g791 ( .A(n_115), .Y(n_791) );
INVxp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_464), .B(n_465), .Y(n_118) );
INVx1_ASAP7_75t_L g463 ( .A(n_120), .Y(n_463) );
AOI22x1_ASAP7_75t_L g476 ( .A1(n_120), .A2(n_477), .B1(n_478), .B2(n_776), .Y(n_476) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_121), .A2(n_477), .B1(n_479), .B2(n_776), .Y(n_780) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_387), .Y(n_121) );
NOR2xp67_ASAP7_75t_L g122 ( .A(n_123), .B(n_306), .Y(n_122) );
NAND5xp2_ASAP7_75t_L g123 ( .A(n_124), .B(n_250), .C(n_260), .D(n_277), .E(n_293), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_184), .B1(n_227), .B2(n_231), .Y(n_125) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_158), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g233 ( .A(n_128), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g252 ( .A(n_128), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g273 ( .A(n_128), .B(n_274), .Y(n_273) );
INVx4_ASAP7_75t_L g287 ( .A(n_128), .Y(n_287) );
AND2x2_ASAP7_75t_L g296 ( .A(n_128), .B(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_SL g318 ( .A(n_128), .B(n_235), .Y(n_318) );
BUFx2_ASAP7_75t_L g361 ( .A(n_128), .Y(n_361) );
AND2x2_ASAP7_75t_L g376 ( .A(n_128), .B(n_159), .Y(n_376) );
OR2x2_ASAP7_75t_L g408 ( .A(n_128), .B(n_409), .Y(n_408) );
NOR4xp25_ASAP7_75t_L g457 ( .A(n_128), .B(n_458), .C(n_459), .D(n_460), .Y(n_457) );
OR2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_155), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_139), .B(n_151), .Y(n_129) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_137), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
AND2x6_ASAP7_75t_L g149 ( .A(n_133), .B(n_142), .Y(n_149) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g147 ( .A(n_135), .B(n_144), .Y(n_147) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx5_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
AND2x2_ASAP7_75t_L g143 ( .A(n_138), .B(n_144), .Y(n_143) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_138), .Y(n_176) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
BUFx3_ASAP7_75t_L g177 ( .A(n_141), .Y(n_177) );
INVx2_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
AND2x4_ASAP7_75t_L g179 ( .A(n_143), .B(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_148), .B(n_150), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_149), .B(n_203), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_150), .A2(n_164), .B(n_165), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_150), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_150), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_150), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_150), .A2(n_225), .B(n_226), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_150), .A2(n_241), .B(n_242), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_150), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_150), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_150), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_150), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_150), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_150), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_150), .A2(n_561), .B(n_562), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_150), .A2(n_570), .B(n_571), .Y(n_569) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_151), .A2(n_172), .B(n_178), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_151), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_151), .A2(n_488), .B(n_489), .Y(n_487) );
OA21x2_ASAP7_75t_L g567 ( .A1(n_151), .A2(n_568), .B(n_572), .Y(n_567) );
OA21x2_ASAP7_75t_L g612 ( .A1(n_151), .A2(n_568), .B(n_572), .Y(n_612) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x4_ASAP7_75t_L g195 ( .A(n_153), .B(n_154), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_156), .A2(n_198), .B(n_199), .Y(n_197) );
BUFx4f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g160 ( .A(n_157), .Y(n_160) );
AOI31xp33_ASAP7_75t_L g325 ( .A1(n_158), .A2(n_326), .A3(n_328), .B(n_330), .Y(n_325) );
INVx2_ASAP7_75t_SL g442 ( .A(n_158), .Y(n_442) );
OR2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_169), .Y(n_158) );
INVx2_ASAP7_75t_L g249 ( .A(n_159), .Y(n_249) );
AND2x2_ASAP7_75t_L g253 ( .A(n_159), .B(n_236), .Y(n_253) );
INVx2_ASAP7_75t_L g276 ( .A(n_159), .Y(n_276) );
AND2x2_ASAP7_75t_L g295 ( .A(n_159), .B(n_235), .Y(n_295) );
AO21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_167), .Y(n_159) );
INVx4_ASAP7_75t_L g168 ( .A(n_160), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_166), .Y(n_161) );
INVx3_ASAP7_75t_L g209 ( .A(n_168), .Y(n_209) );
AND2x2_ASAP7_75t_L g247 ( .A(n_169), .B(n_248), .Y(n_247) );
BUFx3_ASAP7_75t_L g254 ( .A(n_169), .Y(n_254) );
INVx2_ASAP7_75t_L g272 ( .A(n_169), .Y(n_272) );
AND2x2_ASAP7_75t_L g327 ( .A(n_169), .B(n_287), .Y(n_327) );
AND2x4_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
AND2x4_ASAP7_75t_L g298 ( .A(n_170), .B(n_171), .Y(n_298) );
AND2x4_ASAP7_75t_L g173 ( .A(n_174), .B(n_177), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
NOR2x1p5_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_217), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_205), .Y(n_185) );
OR2x2_ASAP7_75t_L g227 ( .A(n_186), .B(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g379 ( .A(n_186), .Y(n_379) );
OR2x2_ASAP7_75t_L g427 ( .A(n_186), .B(n_428), .Y(n_427) );
NAND2x1_ASAP7_75t_L g186 ( .A(n_187), .B(n_196), .Y(n_186) );
OR2x2_ASAP7_75t_SL g218 ( .A(n_187), .B(n_219), .Y(n_218) );
INVx4_ASAP7_75t_L g257 ( .A(n_187), .Y(n_257) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_187), .Y(n_301) );
INVx2_ASAP7_75t_L g309 ( .A(n_187), .Y(n_309) );
OR2x2_ASAP7_75t_L g344 ( .A(n_187), .B(n_207), .Y(n_344) );
AND2x2_ASAP7_75t_L g456 ( .A(n_187), .B(n_311), .Y(n_456) );
AND2x2_ASAP7_75t_L g461 ( .A(n_187), .B(n_220), .Y(n_461) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_195), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_195), .A2(n_222), .B(n_223), .Y(n_221) );
INVx1_ASAP7_75t_SL g496 ( .A(n_195), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_195), .B(n_525), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_195), .A2(n_540), .B(n_541), .Y(n_539) );
OR2x2_ASAP7_75t_L g219 ( .A(n_196), .B(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g285 ( .A(n_196), .B(n_206), .Y(n_285) );
OR2x2_ASAP7_75t_L g292 ( .A(n_196), .B(n_257), .Y(n_292) );
NOR2x1_ASAP7_75t_SL g311 ( .A(n_196), .B(n_230), .Y(n_311) );
BUFx2_ASAP7_75t_L g343 ( .A(n_196), .Y(n_343) );
AND2x2_ASAP7_75t_L g352 ( .A(n_196), .B(n_257), .Y(n_352) );
AND2x2_ASAP7_75t_L g385 ( .A(n_196), .B(n_305), .Y(n_385) );
INVx2_ASAP7_75t_SL g394 ( .A(n_196), .Y(n_394) );
AND2x2_ASAP7_75t_L g397 ( .A(n_196), .B(n_207), .Y(n_397) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_204), .Y(n_196) );
NAND3xp33_ASAP7_75t_L g392 ( .A(n_205), .B(n_262), .C(n_347), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_205), .B(n_309), .Y(n_412) );
INVxp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_206), .B(n_394), .Y(n_415) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_207), .Y(n_259) );
AND2x2_ASAP7_75t_L g303 ( .A(n_207), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g368 ( .A(n_207), .B(n_369), .Y(n_368) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_216), .Y(n_208) );
AO21x1_ASAP7_75t_SL g230 ( .A1(n_209), .A2(n_210), .B(n_216), .Y(n_230) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_209), .A2(n_528), .B(n_534), .Y(n_527) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_209), .A2(n_528), .B(n_534), .Y(n_549) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_209), .A2(n_558), .B(n_564), .Y(n_557) );
AO21x2_ASAP7_75t_L g582 ( .A1(n_209), .A2(n_558), .B(n_564), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_215), .Y(n_210) );
AND2x4_ASAP7_75t_L g263 ( .A(n_217), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g399 ( .A(n_219), .B(n_344), .Y(n_399) );
AND2x2_ASAP7_75t_L g229 ( .A(n_220), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g267 ( .A(n_220), .Y(n_267) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_220), .Y(n_284) );
INVx2_ASAP7_75t_L g305 ( .A(n_220), .Y(n_305) );
INVx1_ASAP7_75t_L g369 ( .A(n_220), .Y(n_369) );
INVx2_ASAP7_75t_L g451 ( .A(n_227), .Y(n_451) );
OR2x2_ASAP7_75t_L g315 ( .A(n_228), .B(n_292), .Y(n_315) );
INVx2_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g455 ( .A(n_229), .B(n_352), .Y(n_455) );
AND2x2_ASAP7_75t_L g348 ( .A(n_230), .B(n_305), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_245), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_233), .A2(n_362), .B1(n_379), .B2(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g275 ( .A(n_235), .Y(n_275) );
AND2x2_ASAP7_75t_L g329 ( .A(n_235), .B(n_249), .Y(n_329) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_235), .Y(n_356) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_236), .Y(n_324) );
AOI21x1_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_244), .Y(n_236) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_237), .A2(n_507), .B(n_513), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_243), .Y(n_238) );
INVxp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_247), .B(n_361), .Y(n_360) );
OAI32xp33_ASAP7_75t_L g377 ( .A1(n_247), .A2(n_378), .A3(n_380), .B1(n_381), .B2(n_383), .Y(n_377) );
BUFx2_ASAP7_75t_L g262 ( .A(n_248), .Y(n_262) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g404 ( .A(n_249), .B(n_298), .Y(n_404) );
OR4x1_ASAP7_75t_L g250 ( .A(n_251), .B(n_254), .C(n_255), .D(n_258), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_251), .A2(n_342), .B1(n_436), .B2(n_437), .Y(n_435) );
INVx2_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_252), .Y(n_444) );
AND2x2_ASAP7_75t_L g286 ( .A(n_253), .B(n_287), .Y(n_286) );
BUFx2_ASAP7_75t_L g366 ( .A(n_253), .Y(n_366) );
INVx1_ASAP7_75t_L g382 ( .A(n_253), .Y(n_382) );
INVx1_ASAP7_75t_L g417 ( .A(n_253), .Y(n_417) );
OR2x2_ASAP7_75t_L g374 ( .A(n_254), .B(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g418 ( .A(n_254), .B(n_419), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_255), .A2(n_292), .B1(n_336), .B2(n_355), .Y(n_357) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g401 ( .A(n_256), .B(n_310), .Y(n_401) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
BUFx2_ASAP7_75t_L g268 ( .A(n_257), .Y(n_268) );
NOR2xp67_ASAP7_75t_L g283 ( .A(n_257), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g264 ( .A(n_258), .Y(n_264) );
NAND4xp25_ASAP7_75t_L g391 ( .A(n_258), .B(n_262), .C(n_343), .D(n_355), .Y(n_391) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g428 ( .A(n_259), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_263), .B1(n_265), .B2(n_269), .Y(n_260) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_261), .A2(n_262), .B1(n_412), .B2(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVxp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx3_ASAP7_75t_L g290 ( .A(n_267), .Y(n_290) );
AOI32xp33_ASAP7_75t_L g406 ( .A1(n_267), .A2(n_407), .A3(n_411), .B1(n_416), .B2(n_420), .Y(n_406) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_273), .Y(n_269) );
NOR2xp67_ASAP7_75t_L g312 ( .A(n_270), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g365 ( .A(n_270), .B(n_366), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_270), .A2(n_278), .B1(n_390), .B2(n_395), .C(n_398), .Y(n_389) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g322 ( .A(n_271), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g437 ( .A(n_271), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_272), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g279 ( .A(n_274), .Y(n_279) );
AND2x2_ASAP7_75t_L g297 ( .A(n_274), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_SL g337 ( .A(n_275), .Y(n_337) );
INVx1_ASAP7_75t_L g321 ( .A(n_276), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_280), .B1(n_286), .B2(n_288), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g423 ( .A(n_279), .B(n_353), .Y(n_423) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g363 ( .A(n_282), .Y(n_363) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
AND2x2_ASAP7_75t_L g294 ( .A(n_287), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_287), .B(n_324), .Y(n_323) );
NAND2x1p5_ASAP7_75t_L g336 ( .A(n_287), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_287), .B(n_329), .Y(n_450) );
AOI22xp33_ASAP7_75t_SL g447 ( .A1(n_288), .A2(n_448), .B1(n_449), .B2(n_451), .Y(n_447) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
OR2x2_ASAP7_75t_L g330 ( .A(n_290), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g340 ( .A(n_290), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_290), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_290), .B(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_SL g395 ( .A(n_290), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g371 ( .A(n_292), .B(n_372), .Y(n_371) );
OAI21xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_296), .B(n_299), .Y(n_293) );
INVx1_ASAP7_75t_L g313 ( .A(n_295), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_296), .A2(n_333), .B1(n_340), .B2(n_345), .Y(n_332) );
INVx3_ASAP7_75t_L g335 ( .A(n_298), .Y(n_335) );
INVx2_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
OAI32xp33_ASAP7_75t_SL g390 ( .A1(n_301), .A2(n_361), .A3(n_391), .B1(n_392), .B2(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g310 ( .A(n_304), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND4xp25_ASAP7_75t_SL g306 ( .A(n_307), .B(n_332), .C(n_349), .D(n_364), .Y(n_306) );
AOI221xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_312), .B1(n_314), .B2(n_316), .C(n_325), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx2_ASAP7_75t_L g347 ( .A(n_309), .Y(n_347) );
AND2x2_ASAP7_75t_L g396 ( .A(n_309), .B(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_309), .B(n_348), .Y(n_434) );
AND2x2_ASAP7_75t_L g445 ( .A(n_309), .B(n_368), .Y(n_445) );
INVx2_ASAP7_75t_L g331 ( .A(n_311), .Y(n_331) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI21xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_319), .B(n_322), .Y(n_316) );
AND2x2_ASAP7_75t_L g448 ( .A(n_317), .B(n_319), .Y(n_448) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_318), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g425 ( .A(n_323), .Y(n_425) );
INVx1_ASAP7_75t_L g410 ( .A(n_324), .Y(n_410) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_327), .B(n_382), .Y(n_381) );
NOR2x1_ASAP7_75t_L g339 ( .A(n_328), .B(n_335), .Y(n_339) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g438 ( .A(n_329), .Y(n_438) );
INVx1_ASAP7_75t_L g420 ( .A(n_331), .Y(n_420) );
OR2x2_ASAP7_75t_L g436 ( .A(n_331), .B(n_347), .Y(n_436) );
NAND2xp33_ASAP7_75t_SL g333 ( .A(n_334), .B(n_338), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx2_ASAP7_75t_L g353 ( .A(n_335), .Y(n_353) );
AND2x2_ASAP7_75t_L g358 ( .A(n_335), .B(n_348), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_335), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g432 ( .A(n_336), .Y(n_432) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_341), .A2(n_422), .B1(n_424), .B2(n_426), .Y(n_421) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g386 ( .A(n_344), .Y(n_386) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g372 ( .A(n_348), .Y(n_372) );
AOI322xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_353), .A3(n_354), .B1(n_357), .B2(n_358), .C1(n_359), .C2(n_362), .Y(n_349) );
OAI21xp5_ASAP7_75t_SL g400 ( .A1(n_350), .A2(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g367 ( .A(n_352), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g424 ( .A(n_353), .B(n_425), .Y(n_424) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_360), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g380 ( .A(n_361), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_361), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B1(n_370), .B2(n_373), .C(n_377), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_366), .A2(n_453), .B1(n_455), .B2(n_456), .C(n_457), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_368), .B(n_379), .Y(n_378) );
BUFx2_ASAP7_75t_L g419 ( .A(n_369), .Y(n_419) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OAI21xp5_ASAP7_75t_L g443 ( .A1(n_373), .A2(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp33_ASAP7_75t_SL g453 ( .A(n_382), .B(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
NOR4xp75_ASAP7_75t_L g387 ( .A(n_388), .B(n_405), .C(n_429), .D(n_446), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_400), .Y(n_388) );
INVx1_ASAP7_75t_L g459 ( .A(n_397), .Y(n_459) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g431 ( .A(n_404), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g458 ( .A(n_404), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_406), .B(n_421), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_SL g454 ( .A(n_425), .Y(n_454) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND3x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_439), .C(n_443), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B(n_435), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_452), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_464), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g790 ( .A(n_471), .B(n_791), .Y(n_790) );
AOI31xp33_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_778), .A3(n_781), .B(n_787), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_661), .Y(n_479) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_616), .C(n_645), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_482), .B(n_589), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_514), .B1(n_535), .B2(n_546), .C(n_550), .Y(n_482) );
INVx3_ASAP7_75t_SL g706 ( .A(n_483), .Y(n_706) );
AND2x2_ASAP7_75t_SL g483 ( .A(n_484), .B(n_493), .Y(n_483) );
NAND2x1p5_ASAP7_75t_L g552 ( .A(n_484), .B(n_505), .Y(n_552) );
INVx4_ASAP7_75t_L g587 ( .A(n_484), .Y(n_587) );
AND2x2_ASAP7_75t_L g609 ( .A(n_484), .B(n_506), .Y(n_609) );
AND2x2_ASAP7_75t_L g615 ( .A(n_484), .B(n_554), .Y(n_615) );
INVx5_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx2_ASAP7_75t_L g584 ( .A(n_485), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_485), .B(n_505), .Y(n_660) );
AND2x2_ASAP7_75t_L g665 ( .A(n_485), .B(n_506), .Y(n_665) );
AND2x2_ASAP7_75t_L g677 ( .A(n_485), .B(n_538), .Y(n_677) );
NOR2x1_ASAP7_75t_SL g716 ( .A(n_485), .B(n_554), .Y(n_716) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
INVx2_ASAP7_75t_L g545 ( .A(n_493), .Y(n_545) );
AND2x2_ASAP7_75t_L g649 ( .A(n_493), .B(n_598), .Y(n_649) );
AND2x2_ASAP7_75t_L g746 ( .A(n_493), .B(n_677), .Y(n_746) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_505), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g578 ( .A(n_495), .Y(n_578) );
INVx2_ASAP7_75t_L g600 ( .A(n_495), .Y(n_600) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B(n_503), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_496), .B(n_504), .Y(n_503) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_496), .A2(n_497), .B(n_503), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_502), .Y(n_497) );
AND2x2_ASAP7_75t_L g575 ( .A(n_505), .B(n_537), .Y(n_575) );
INVx2_ASAP7_75t_L g579 ( .A(n_505), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_505), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g678 ( .A(n_505), .B(n_643), .Y(n_678) );
OR2x2_ASAP7_75t_L g725 ( .A(n_505), .B(n_538), .Y(n_725) );
INVx4_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_506), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .Y(n_507) );
AND2x2_ASAP7_75t_L g722 ( .A(n_514), .B(n_603), .Y(n_722) );
AND2x2_ASAP7_75t_L g772 ( .A(n_514), .B(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g648 ( .A(n_515), .B(n_592), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_526), .Y(n_515) );
AND2x2_ASAP7_75t_L g581 ( .A(n_516), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g611 ( .A(n_516), .B(n_612), .Y(n_611) );
AND2x4_ASAP7_75t_L g632 ( .A(n_516), .B(n_612), .Y(n_632) );
AND2x4_ASAP7_75t_L g667 ( .A(n_516), .B(n_655), .Y(n_667) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g548 ( .A(n_517), .Y(n_548) );
OAI21x1_ASAP7_75t_SL g517 ( .A1(n_518), .A2(n_520), .B(n_524), .Y(n_517) );
INVx1_ASAP7_75t_L g525 ( .A(n_519), .Y(n_525) );
AND2x2_ASAP7_75t_L g594 ( .A(n_526), .B(n_547), .Y(n_594) );
AND2x2_ASAP7_75t_L g680 ( .A(n_526), .B(n_612), .Y(n_680) );
AND2x2_ASAP7_75t_L g691 ( .A(n_526), .B(n_556), .Y(n_691) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g555 ( .A(n_527), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g622 ( .A(n_527), .B(n_557), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_529), .B(n_533), .Y(n_528) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_545), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_537), .B(n_587), .Y(n_644) );
AND2x2_ASAP7_75t_L g688 ( .A(n_537), .B(n_554), .Y(n_688) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_538), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g598 ( .A(n_538), .Y(n_598) );
BUFx3_ASAP7_75t_L g607 ( .A(n_538), .Y(n_607) );
AND2x2_ASAP7_75t_L g630 ( .A(n_538), .B(n_600), .Y(n_630) );
OAI322xp33_ASAP7_75t_L g550 ( .A1(n_545), .A2(n_551), .A3(n_555), .B1(n_565), .B2(n_573), .C1(n_580), .C2(n_585), .Y(n_550) );
INVx1_ASAP7_75t_L g711 ( .A(n_545), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_546), .B(n_586), .Y(n_585) );
AND2x4_ASAP7_75t_L g624 ( .A(n_546), .B(n_566), .Y(n_624) );
INVx2_ASAP7_75t_L g669 ( .A(n_546), .Y(n_669) );
AND2x2_ASAP7_75t_L g685 ( .A(n_546), .B(n_627), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_546), .B(n_703), .Y(n_733) );
AND2x4_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
AND2x2_ASAP7_75t_SL g636 ( .A(n_547), .B(n_612), .Y(n_636) );
OR2x2_ASAP7_75t_L g657 ( .A(n_547), .B(n_574), .Y(n_657) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx2_ASAP7_75t_L g629 ( .A(n_548), .Y(n_629) );
INVx2_ASAP7_75t_L g574 ( .A(n_549), .Y(n_574) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_549), .Y(n_576) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx2_ASAP7_75t_L g619 ( .A(n_552), .Y(n_619) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_553), .Y(n_639) );
INVx1_ASAP7_75t_L g737 ( .A(n_553), .Y(n_737) );
INVxp67_ASAP7_75t_SL g752 ( .A(n_553), .Y(n_752) );
NAND2x1_ASAP7_75t_L g762 ( .A(n_555), .B(n_566), .Y(n_762) );
INVx1_ASAP7_75t_L g769 ( .A(n_555), .Y(n_769) );
BUFx2_ASAP7_75t_L g603 ( .A(n_556), .Y(n_603) );
AND2x2_ASAP7_75t_L g679 ( .A(n_556), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx3_ASAP7_75t_L g588 ( .A(n_557), .Y(n_588) );
INVxp67_ASAP7_75t_L g592 ( .A(n_557), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_563), .Y(n_558) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_565), .B(n_581), .C(n_583), .Y(n_580) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_SL g601 ( .A(n_566), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_566), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g753 ( .A(n_566), .B(n_702), .Y(n_753) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g655 ( .A(n_567), .Y(n_655) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_567), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_573) );
AND2x4_ASAP7_75t_SL g702 ( .A(n_574), .B(n_582), .Y(n_702) );
AND2x2_ASAP7_75t_L g715 ( .A(n_575), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_576), .Y(n_717) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx2_ASAP7_75t_L g674 ( .A(n_578), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_578), .B(n_587), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_579), .B(n_597), .Y(n_596) );
AND3x2_ASAP7_75t_L g614 ( .A(n_579), .B(n_607), .C(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g638 ( .A(n_579), .Y(n_638) );
AND2x2_ASAP7_75t_L g751 ( .A(n_579), .B(n_752), .Y(n_751) );
BUFx2_ASAP7_75t_L g627 ( .A(n_582), .Y(n_627) );
INVx1_ASAP7_75t_L g705 ( .A(n_582), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_583), .B(n_606), .Y(n_744) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_584), .B(n_688), .Y(n_693) );
AND2x4_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
AND2x2_ASAP7_75t_L g684 ( .A(n_587), .B(n_630), .Y(n_684) );
INVx1_ASAP7_75t_SL g635 ( .A(n_588), .Y(n_635) );
AND2x2_ASAP7_75t_L g743 ( .A(n_588), .B(n_655), .Y(n_743) );
AND2x2_ASAP7_75t_L g764 ( .A(n_588), .B(n_636), .Y(n_764) );
AOI221xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_595), .B1(n_601), .B2(n_604), .C(n_610), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g756 ( .A(n_592), .Y(n_756) );
AOI21xp33_ASAP7_75t_SL g610 ( .A1(n_593), .A2(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g602 ( .A(n_594), .B(n_603), .Y(n_602) );
AOI222xp33_ASAP7_75t_L g625 ( .A1(n_594), .A2(n_626), .B1(n_628), .B2(n_633), .C1(n_637), .C2(n_640), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_594), .B(n_743), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_595), .A2(n_624), .B1(n_647), .B2(n_649), .Y(n_646) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g631 ( .A(n_598), .Y(n_631) );
AND2x2_ASAP7_75t_L g750 ( .A(n_598), .B(n_716), .Y(n_750) );
OAI32xp33_ASAP7_75t_L g754 ( .A1(n_598), .A2(n_623), .A3(n_675), .B1(n_683), .B2(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g759 ( .A(n_598), .B(n_609), .Y(n_759) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g643 ( .A(n_600), .Y(n_643) );
OAI21xp5_ASAP7_75t_SL g650 ( .A1(n_601), .A2(n_651), .B(n_658), .Y(n_650) );
INVx1_ASAP7_75t_L g714 ( .A(n_603), .Y(n_714) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
AND2x2_ASAP7_75t_L g618 ( .A(n_606), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g626 ( .A(n_609), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g699 ( .A(n_609), .B(n_630), .Y(n_699) );
INVx1_ASAP7_75t_SL g770 ( .A(n_611), .Y(n_770) );
AND2x2_ASAP7_75t_L g704 ( .A(n_612), .B(n_705), .Y(n_704) );
OAI222xp33_ASAP7_75t_L g757 ( .A1(n_613), .A2(n_666), .B1(n_745), .B2(n_758), .C1(n_760), .C2(n_762), .Y(n_757) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x4_ASAP7_75t_L g730 ( .A(n_615), .B(n_731), .Y(n_730) );
OAI21xp33_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_620), .B(n_625), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_619), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g698 ( .A(n_621), .Y(n_698) );
INVx1_ASAP7_75t_L g666 ( .A(n_622), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_622), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g720 ( .A(n_627), .Y(n_720) );
AO22x1_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_628) );
OAI322xp33_ASAP7_75t_L g740 ( .A1(n_629), .A2(n_690), .A3(n_693), .B1(n_741), .B2(n_742), .C1(n_744), .C2(n_745), .Y(n_740) );
AND2x2_ASAP7_75t_SL g664 ( .A(n_630), .B(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g659 ( .A(n_631), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_632), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g761 ( .A(n_632), .B(n_691), .Y(n_761) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g741 ( .A(n_635), .Y(n_741) );
INVx1_ASAP7_75t_SL g670 ( .A(n_636), .Y(n_670) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
OR2x2_ASAP7_75t_L g672 ( .A(n_644), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g710 ( .A(n_644), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_650), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_656), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g683 ( .A(n_654), .B(n_669), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_654), .B(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g713 ( .A(n_657), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_662), .B(n_726), .Y(n_661) );
NAND4xp25_ASAP7_75t_L g662 ( .A(n_663), .B(n_681), .C(n_694), .D(n_707), .Y(n_662) );
AOI322xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .A3(n_667), .B1(n_668), .B2(n_671), .C1(n_676), .C2(n_679), .Y(n_663) );
AOI211xp5_ASAP7_75t_L g763 ( .A1(n_664), .A2(n_764), .B(n_765), .C(n_768), .Y(n_763) );
AND2x2_ASAP7_75t_L g775 ( .A(n_665), .B(n_752), .Y(n_775) );
INVx1_ASAP7_75t_L g697 ( .A(n_667), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_667), .B(n_702), .Y(n_739) );
NAND2xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_675), .B(n_688), .Y(n_755) );
AND2x4_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B1(n_685), .B2(n_686), .C1(n_689), .C2(n_692), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_684), .A2(n_695), .B1(n_698), .B2(n_699), .C(n_700), .Y(n_694) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI21xp33_ASAP7_75t_SL g700 ( .A1(n_701), .A2(n_703), .B(n_706), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_712), .B1(n_715), .B2(n_717), .C(n_718), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g767 ( .A(n_716), .Y(n_767) );
AOI21xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_721), .B(n_723), .Y(n_718) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx2_ASAP7_75t_L g731 ( .A(n_725), .Y(n_731) );
OR2x2_ASAP7_75t_L g766 ( .A(n_725), .B(n_767), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_747), .C(n_763), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_740), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_732), .B(n_734), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_738), .Y(n_734) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI221xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_753), .B1(n_754), .B2(n_756), .C(n_757), .Y(n_747) );
INVxp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NOR2x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_762), .B(n_766), .Y(n_765) );
O2A1O1Ixp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .B(n_771), .C(n_774), .Y(n_768) );
INVxp67_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
CKINVDCx11_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVxp67_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx3_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_792), .Y(n_788) );
INVxp67_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
endmodule