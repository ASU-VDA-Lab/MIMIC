module fake_jpeg_7483_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_17),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_24),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_26),
.B1(n_22),
.B2(n_27),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_46),
.B1(n_17),
.B2(n_19),
.Y(n_55)
);

INVx5_ASAP7_75t_SL g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_24),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_26),
.B1(n_27),
.B2(n_25),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_4),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_3),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_52),
.B(n_58),
.C(n_69),
.Y(n_84)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_59),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

AND2x6_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_3),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_54),
.Y(n_72)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_31),
.B1(n_29),
.B2(n_19),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_29),
.B1(n_15),
.B2(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_61),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_64),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_28),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_8),
.B(n_11),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_15),
.B1(n_18),
.B2(n_14),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_20),
.B(n_14),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_5),
.B(n_6),
.Y(n_77)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_38),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_50),
.C(n_47),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_89),
.C(n_92),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_93),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_94),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_52),
.B1(n_68),
.B2(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_49),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_100),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_61),
.B1(n_11),
.B2(n_12),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_77),
.Y(n_108)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_79),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_84),
.B(n_81),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_95),
.B(n_84),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_87),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_111),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_117),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_106),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_119),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_101),
.C(n_108),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_101),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_80),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_80),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_76),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_128),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_103),
.B(n_120),
.C(n_124),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_105),
.C(n_110),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_130),
.B1(n_75),
.B2(n_88),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);

OAI21x1_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_70),
.B(n_75),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_136),
.B(n_132),
.Y(n_138)
);

AOI221xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_126),
.B1(n_70),
.B2(n_12),
.C(n_79),
.Y(n_139)
);


endmodule