module fake_jpeg_1995_n_188 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_16),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_32),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_31),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_5),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_69),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_73),
.Y(n_83)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_67),
.B1(n_55),
.B2(n_63),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_86),
.B1(n_74),
.B2(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_49),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_79),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_67),
.B1(n_55),
.B2(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

BUFx2_ASAP7_75t_SL g89 ( 
.A(n_88),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_72),
.B(n_75),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_57),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_98),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

XOR2x2_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_57),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_101),
.C(n_104),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_52),
.C(n_58),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_47),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_48),
.B1(n_2),
.B2(n_3),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_61),
.C(n_60),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_18),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_80),
.B1(n_56),
.B2(n_54),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_103),
.B1(n_5),
.B2(n_6),
.Y(n_132)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_0),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_119),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_48),
.B1(n_59),
.B2(n_3),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_122),
.B1(n_10),
.B2(n_11),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_1),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_22),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_1),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_2),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_92),
.B(n_89),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_136),
.B(n_46),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_133),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_25),
.B1(n_44),
.B2(n_42),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_8),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_143),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_8),
.B(n_9),
.Y(n_136)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_142),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_26),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_134),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_11),
.B(n_12),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_141),
.A2(n_15),
.B(n_27),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_144),
.B(n_145),
.Y(n_148)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_109),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_30),
.C(n_41),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_161),
.C(n_162),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_14),
.A3(n_15),
.B1(n_23),
.B2(n_24),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_132),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_157),
.B(n_159),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_131),
.B(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_125),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_158),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_126),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_162),
.B(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_166),
.Y(n_175)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

BUFx12f_ASAP7_75t_SL g171 ( 
.A(n_165),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_171),
.A2(n_168),
.B(n_148),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_147),
.B(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_174),
.Y(n_180)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_169),
.B(n_151),
.CI(n_153),
.CON(n_174),
.SN(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_175),
.B1(n_171),
.B2(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_181),
.B(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_182),
.Y(n_184)
);

NOR2x1_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_180),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_173),
.C(n_155),
.Y(n_186)
);

AO21x1_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_152),
.B(n_174),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_150),
.Y(n_188)
);


endmodule