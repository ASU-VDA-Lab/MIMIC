module fake_aes_11015_n_631 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_631);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_631;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_599;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g73 ( .A(n_63), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_69), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_36), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_41), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_47), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_34), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_65), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_22), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_3), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_19), .Y(n_82) );
BUFx10_ASAP7_75t_L g83 ( .A(n_46), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_6), .Y(n_84) );
NOR2xp33_ASAP7_75t_L g85 ( .A(n_17), .B(n_62), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_4), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_0), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_35), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_26), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_72), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_57), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_44), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_59), .Y(n_93) );
BUFx2_ASAP7_75t_SL g94 ( .A(n_42), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_30), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_7), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_40), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_14), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_8), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_58), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_50), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_28), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_43), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_51), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_67), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_27), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_23), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_66), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_21), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_7), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_8), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_70), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_12), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_53), .Y(n_114) );
BUFx5_ASAP7_75t_L g115 ( .A(n_32), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_52), .Y(n_116) );
NOR2x1_ASAP7_75t_L g117 ( .A(n_86), .B(n_25), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_115), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_110), .Y(n_119) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_102), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_120) );
CKINVDCx8_ASAP7_75t_R g121 ( .A(n_94), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_87), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_83), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_107), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
INVx1_ASAP7_75t_SL g126 ( .A(n_84), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_96), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_98), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_111), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_107), .B(n_1), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_102), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_108), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_99), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_106), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_110), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_108), .B(n_2), .Y(n_137) );
INVx4_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
NOR2x1_ASAP7_75t_L g139 ( .A(n_73), .B(n_31), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_115), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_74), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_106), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_112), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_75), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_88), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_112), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_115), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_82), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_115), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_89), .B(n_3), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_90), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_115), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_91), .B(n_4), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_92), .B(n_116), .Y(n_154) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_93), .B(n_33), .Y(n_155) );
AND2x6_ASAP7_75t_L g156 ( .A(n_95), .B(n_37), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_124), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_124), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_130), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_130), .Y(n_160) );
NAND3xp33_ASAP7_75t_L g161 ( .A(n_127), .B(n_101), .C(n_114), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_130), .B(n_115), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_138), .B(n_97), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_135), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_124), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_138), .B(n_113), .Y(n_167) );
OR2x6_ASAP7_75t_L g168 ( .A(n_138), .B(n_100), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_123), .B(n_76), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_125), .Y(n_170) );
INVx5_ASAP7_75t_L g171 ( .A(n_156), .Y(n_171) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_156), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_123), .B(n_115), .Y(n_173) );
AO22x1_ASAP7_75t_L g174 ( .A1(n_156), .A2(n_80), .B1(n_105), .B2(n_104), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_150), .B(n_109), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_150), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_133), .B(n_103), .Y(n_177) );
INVx1_ASAP7_75t_SL g178 ( .A(n_126), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_150), .B(n_85), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_141), .B(n_79), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_134), .A2(n_78), .B1(n_77), .B2(n_85), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_132), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
NAND2xp33_ASAP7_75t_L g186 ( .A(n_156), .B(n_29), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_118), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_155), .B(n_38), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_144), .B(n_5), .Y(n_190) );
AND2x6_ASAP7_75t_L g191 ( .A(n_139), .B(n_71), .Y(n_191) );
INVxp67_ASAP7_75t_SL g192 ( .A(n_154), .Y(n_192) );
INVx1_ASAP7_75t_SL g193 ( .A(n_143), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_122), .B(n_5), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_118), .Y(n_195) );
OR2x6_ASAP7_75t_L g196 ( .A(n_153), .B(n_6), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_128), .B(n_9), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_129), .Y(n_198) );
AND2x6_ASAP7_75t_L g199 ( .A(n_117), .B(n_39), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_132), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_155), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_145), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_148), .B(n_13), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_156), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_132), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_132), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_137), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_140), .B(n_48), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_172), .B(n_121), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_172), .B(n_152), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_172), .B(n_152), .Y(n_211) );
NOR2xp33_ASAP7_75t_R g212 ( .A(n_165), .B(n_131), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_192), .B(n_147), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_207), .B(n_147), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_160), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_178), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_171), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_188), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_198), .B(n_146), .Y(n_219) );
INVxp67_ASAP7_75t_L g220 ( .A(n_170), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_162), .A2(n_149), .B(n_140), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_171), .B(n_149), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_188), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_171), .B(n_146), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_160), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_188), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_164), .B(n_181), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_167), .B(n_142), .Y(n_228) );
INVx1_ASAP7_75t_SL g229 ( .A(n_193), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_160), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_173), .Y(n_231) );
INVx1_ASAP7_75t_SL g232 ( .A(n_165), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_194), .B(n_142), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_195), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_176), .B(n_131), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_195), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_173), .Y(n_237) );
INVx5_ASAP7_75t_L g238 ( .A(n_163), .Y(n_238) );
INVx5_ASAP7_75t_L g239 ( .A(n_163), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_195), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_159), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_204), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_175), .B(n_120), .Y(n_243) );
AND2x6_ASAP7_75t_SL g244 ( .A(n_196), .B(n_136), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_163), .Y(n_245) );
NOR2xp33_ASAP7_75t_R g246 ( .A(n_186), .B(n_136), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_175), .B(n_13), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_168), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_171), .B(n_119), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_163), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_196), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_168), .B(n_180), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_204), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_200), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_162), .Y(n_255) );
NOR2x2_ASAP7_75t_L g256 ( .A(n_196), .B(n_119), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_194), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_197), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_171), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_189), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_168), .B(n_18), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_168), .B(n_20), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_180), .B(n_24), .Y(n_263) );
NAND3xp33_ASAP7_75t_SL g264 ( .A(n_201), .B(n_45), .C(n_49), .Y(n_264) );
INVx5_ASAP7_75t_SL g265 ( .A(n_216), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_225), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_225), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_231), .B(n_189), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_229), .Y(n_269) );
AOI22xp33_ASAP7_75t_SL g270 ( .A1(n_251), .A2(n_196), .B1(n_177), .B2(n_180), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_212), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_251), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_220), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_231), .B(n_180), .Y(n_274) );
AOI221xp5_ASAP7_75t_L g275 ( .A1(n_257), .A2(n_202), .B1(n_190), .B2(n_161), .C(n_203), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_225), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_225), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_227), .A2(n_186), .B(n_174), .Y(n_278) );
INVxp67_ASAP7_75t_L g279 ( .A(n_219), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_232), .B(n_177), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_SL g281 ( .A1(n_258), .A2(n_182), .B(n_179), .C(n_183), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_215), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_257), .B(n_177), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_219), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_233), .B(n_169), .Y(n_285) );
OAI21x1_ASAP7_75t_SL g286 ( .A1(n_252), .A2(n_180), .B(n_185), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_237), .B(n_180), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_243), .B(n_208), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_233), .B(n_179), .Y(n_289) );
BUFx12f_ASAP7_75t_L g290 ( .A(n_244), .Y(n_290) );
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_241), .A2(n_208), .B(n_187), .C(n_179), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_214), .A2(n_158), .B(n_205), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_213), .Y(n_293) );
BUFx4f_ASAP7_75t_L g294 ( .A(n_262), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_256), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_242), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_228), .B(n_199), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_236), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_215), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_242), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_262), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_241), .A2(n_158), .B(n_205), .C(n_184), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_248), .A2(n_235), .B1(n_258), .B2(n_249), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_242), .B(n_206), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_230), .Y(n_305) );
AND2x2_ASAP7_75t_SL g306 ( .A(n_244), .B(n_199), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_221), .A2(n_157), .B(n_184), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_237), .B(n_199), .Y(n_308) );
AND2x2_ASAP7_75t_SL g309 ( .A(n_246), .B(n_199), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_SL g310 ( .A1(n_281), .A2(n_291), .B(n_263), .C(n_302), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_288), .A2(n_255), .B(n_230), .C(n_247), .Y(n_311) );
BUFx12f_ASAP7_75t_L g312 ( .A(n_269), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_282), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_293), .B(n_255), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_299), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_273), .Y(n_317) );
AOI22xp33_ASAP7_75t_SL g318 ( .A1(n_295), .A2(n_294), .B1(n_265), .B2(n_290), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_286), .A2(n_261), .B(n_210), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_305), .Y(n_320) );
OAI21x1_ASAP7_75t_L g321 ( .A1(n_307), .A2(n_211), .B(n_254), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_294), .Y(n_322) );
OAI21x1_ASAP7_75t_SL g323 ( .A1(n_268), .A2(n_260), .B(n_218), .Y(n_323) );
OAI21x1_ASAP7_75t_L g324 ( .A1(n_307), .A2(n_254), .B(n_245), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_266), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_277), .Y(n_326) );
AO21x2_ASAP7_75t_L g327 ( .A1(n_278), .A2(n_264), .B(n_166), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_293), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_276), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_268), .Y(n_330) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_297), .A2(n_240), .B(n_236), .C(n_218), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_276), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_272), .B(n_253), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_265), .B(n_236), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_278), .A2(n_222), .B(n_253), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_274), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_274), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_287), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_328), .A2(n_284), .B1(n_270), .B2(n_306), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_317), .A2(n_279), .B1(n_283), .B2(n_285), .C(n_275), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_312), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_328), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_315), .A2(n_301), .B1(n_309), .B2(n_265), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_312), .B(n_301), .Y(n_344) );
AOI22xp33_ASAP7_75t_SL g345 ( .A1(n_312), .A2(n_271), .B1(n_280), .B2(n_283), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_320), .B(n_287), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_320), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_320), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_315), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_314), .Y(n_350) );
AO221x2_ASAP7_75t_L g351 ( .A1(n_316), .A2(n_267), .B1(n_303), .B2(n_218), .C(n_226), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_310), .A2(n_308), .B(n_304), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_316), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_314), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_315), .A2(n_275), .B1(n_209), .B2(n_289), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_314), .Y(n_356) );
OAI211xp5_ASAP7_75t_L g357 ( .A1(n_318), .A2(n_224), .B(n_240), .C(n_236), .Y(n_357) );
OAI21x1_ASAP7_75t_L g358 ( .A1(n_324), .A2(n_292), .B(n_254), .Y(n_358) );
OA21x2_ASAP7_75t_L g359 ( .A1(n_324), .A2(n_166), .B(n_157), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_330), .Y(n_360) );
AOI31xp33_ASAP7_75t_SL g361 ( .A1(n_334), .A2(n_199), .A3(n_191), .B(n_226), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_330), .A2(n_298), .B1(n_240), .B2(n_199), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_315), .A2(n_240), .B1(n_191), .B2(n_300), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_342), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_347), .B(n_325), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_350), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_347), .B(n_325), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_342), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_348), .B(n_325), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_348), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_354), .Y(n_371) );
OA21x2_ASAP7_75t_L g372 ( .A1(n_358), .A2(n_323), .B(n_321), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_354), .B(n_326), .Y(n_373) );
NOR4xp25_ASAP7_75t_SL g374 ( .A(n_344), .B(n_360), .C(n_356), .D(n_353), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_356), .B(n_326), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_350), .Y(n_376) );
NOR4xp25_ASAP7_75t_SL g377 ( .A(n_360), .B(n_331), .C(n_311), .D(n_336), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_345), .B(n_322), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_346), .B(n_326), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_341), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_346), .B(n_338), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_349), .B(n_338), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_351), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_351), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_351), .B(n_337), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_359), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_341), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_351), .B(n_334), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_359), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_359), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_355), .B(n_337), .Y(n_391) );
OA21x2_ASAP7_75t_L g392 ( .A1(n_358), .A2(n_323), .B(n_321), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_339), .B(n_336), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_359), .B(n_327), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_343), .B(n_327), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_379), .B(n_340), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_370), .B(n_313), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_371), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g399 ( .A(n_378), .B(n_357), .C(n_322), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_393), .B(n_333), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_381), .B(n_327), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_370), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_381), .B(n_327), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_370), .Y(n_404) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_393), .A2(n_329), .B1(n_332), .B2(n_313), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_368), .B(n_313), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_379), .B(n_332), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_376), .Y(n_408) );
OAI33xp33_ASAP7_75t_L g409 ( .A1(n_383), .A2(n_329), .A3(n_332), .B1(n_226), .B2(n_223), .B3(n_234), .Y(n_409) );
OAI22xp5_ASAP7_75t_SL g410 ( .A1(n_380), .A2(n_363), .B1(n_362), .B2(n_361), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_387), .A2(n_352), .B1(n_329), .B2(n_335), .C(n_313), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_385), .B(n_319), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_365), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_365), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_366), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_379), .B(n_333), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_365), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_391), .A2(n_333), .B1(n_191), .B2(n_319), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_376), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_391), .B(n_333), .Y(n_420) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_380), .B(n_234), .C(n_223), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_367), .B(n_206), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_367), .B(n_206), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_391), .B(n_191), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_366), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_367), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_366), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_385), .A2(n_191), .B1(n_296), .B2(n_300), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_369), .B(n_191), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_369), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_385), .B(n_54), .Y(n_431) );
INVx4_ASAP7_75t_L g432 ( .A(n_380), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_388), .A2(n_300), .B1(n_296), .B2(n_253), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_369), .B(n_206), .Y(n_434) );
OAI322xp33_ASAP7_75t_L g435 ( .A1(n_368), .A2(n_200), .A3(n_245), .B1(n_250), .B2(n_61), .C1(n_64), .C2(n_68), .Y(n_435) );
OR2x6_ASAP7_75t_SL g436 ( .A(n_388), .B(n_55), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_376), .A2(n_238), .B(n_239), .Y(n_437) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_373), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_373), .B(n_56), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_373), .B(n_200), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_386), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_438), .B(n_395), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_438), .B(n_395), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_438), .B(n_395), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_438), .B(n_394), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_401), .B(n_394), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_441), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_441), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_403), .B(n_412), .Y(n_449) );
BUFx2_ASAP7_75t_L g450 ( .A(n_408), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_412), .B(n_394), .Y(n_451) );
INVx3_ASAP7_75t_L g452 ( .A(n_419), .Y(n_452) );
NAND4xp25_ASAP7_75t_SL g453 ( .A(n_436), .B(n_383), .C(n_384), .D(n_374), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_412), .B(n_384), .Y(n_454) );
AND2x4_ASAP7_75t_SL g455 ( .A(n_431), .B(n_364), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_404), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_415), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_398), .B(n_389), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_432), .B(n_375), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_404), .B(n_389), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_415), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_425), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_408), .B(n_390), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_425), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_427), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_413), .B(n_390), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_436), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_414), .B(n_390), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_417), .B(n_386), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_427), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_402), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_426), .B(n_386), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_430), .B(n_419), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_419), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_416), .B(n_375), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_396), .B(n_432), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_407), .B(n_382), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_420), .B(n_375), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_400), .B(n_382), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_432), .B(n_392), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_400), .B(n_374), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_406), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_431), .B(n_439), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_431), .B(n_392), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_397), .B(n_392), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_397), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
AND2x2_ASAP7_75t_SL g488 ( .A(n_397), .B(n_392), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_405), .B(n_392), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_434), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_399), .B(n_377), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_409), .B(n_377), .C(n_245), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_421), .B(n_200), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_405), .B(n_372), .Y(n_494) );
NOR3xp33_ASAP7_75t_SL g495 ( .A(n_410), .B(n_60), .C(n_372), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_458), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_455), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_475), .B(n_440), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_475), .B(n_422), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_477), .B(n_423), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_458), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_446), .B(n_372), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_446), .B(n_372), .Y(n_503) );
NAND3xp33_ASAP7_75t_L g504 ( .A(n_467), .B(n_418), .C(n_428), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_466), .B(n_372), .Y(n_505) );
NAND4xp25_ASAP7_75t_L g506 ( .A(n_476), .B(n_418), .C(n_424), .D(n_411), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_445), .B(n_433), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_471), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_479), .B(n_429), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_471), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_466), .B(n_437), .Y(n_511) );
AND3x2_ASAP7_75t_L g512 ( .A(n_487), .B(n_435), .C(n_250), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_445), .B(n_238), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_456), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_482), .B(n_238), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_469), .B(n_238), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_455), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_455), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_469), .B(n_238), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_482), .B(n_238), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_449), .B(n_239), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_449), .B(n_239), .Y(n_522) );
NOR2x1_ASAP7_75t_L g523 ( .A(n_453), .B(n_217), .Y(n_523) );
NAND2x1p5_ASAP7_75t_L g524 ( .A(n_459), .B(n_239), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_456), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_451), .B(n_239), .Y(n_526) );
AOI21xp33_ASAP7_75t_SL g527 ( .A1(n_481), .A2(n_239), .B(n_217), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_450), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_473), .Y(n_529) );
NOR2xp67_ASAP7_75t_SL g530 ( .A(n_483), .B(n_259), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_478), .B(n_217), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_473), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_486), .B(n_451), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_478), .B(n_217), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_454), .B(n_259), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_463), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_447), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_447), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_448), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_454), .B(n_259), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_463), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_480), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_491), .B(n_483), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_448), .Y(n_544) );
OAI221xp5_ASAP7_75t_SL g545 ( .A1(n_504), .A2(n_480), .B1(n_484), .B2(n_450), .C(n_489), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_543), .A2(n_484), .B1(n_488), .B2(n_444), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_499), .Y(n_547) );
INVxp67_ASAP7_75t_L g548 ( .A(n_528), .Y(n_548) );
OAI322xp33_ASAP7_75t_L g549 ( .A1(n_496), .A2(n_501), .A3(n_532), .B1(n_529), .B2(n_498), .C1(n_502), .C2(n_503), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_533), .B(n_442), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_514), .B(n_460), .Y(n_551) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_528), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_542), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_517), .B(n_486), .Y(n_554) );
XOR2xp5_ASAP7_75t_L g555 ( .A(n_500), .B(n_472), .Y(n_555) );
OAI21xp33_ASAP7_75t_L g556 ( .A1(n_542), .A2(n_495), .B(n_488), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_508), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_525), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_510), .Y(n_559) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_523), .B(n_493), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_537), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_536), .B(n_468), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_538), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_539), .Y(n_564) );
NAND2xp33_ASAP7_75t_L g565 ( .A(n_518), .B(n_486), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_497), .A2(n_488), .B1(n_485), .B2(n_468), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_544), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_509), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_568) );
XOR2xp5_ASAP7_75t_L g569 ( .A(n_533), .B(n_472), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_511), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_497), .B(n_486), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_502), .B(n_460), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_507), .B(n_443), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_524), .A2(n_452), .B1(n_485), .B2(n_494), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_511), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_515), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_520), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_506), .A2(n_490), .B1(n_452), .B2(n_474), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_570), .Y(n_579) );
INVxp67_ASAP7_75t_SL g580 ( .A(n_560), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_575), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_551), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_547), .B(n_503), .Y(n_583) );
INVxp67_ASAP7_75t_L g584 ( .A(n_552), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_551), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_557), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_549), .B(n_541), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_548), .B(n_505), .Y(n_588) );
OAI322xp33_ASAP7_75t_L g589 ( .A1(n_555), .A2(n_505), .A3(n_489), .B1(n_494), .B2(n_531), .C1(n_534), .C2(n_516), .Y(n_589) );
OAI211xp5_ASAP7_75t_L g590 ( .A1(n_578), .A2(n_527), .B(n_534), .C(n_531), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_550), .B(n_526), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_559), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g593 ( .A1(n_545), .A2(n_530), .B(n_522), .C(n_521), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_572), .B(n_490), .Y(n_594) );
NOR2xp33_ASAP7_75t_SL g595 ( .A(n_556), .B(n_512), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_558), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_561), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_553), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_572), .B(n_462), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_593), .A2(n_569), .B1(n_545), .B2(n_546), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_587), .B(n_568), .Y(n_601) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_587), .B(n_565), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_579), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_595), .A2(n_566), .B1(n_554), .B2(n_574), .Y(n_604) );
OAI211xp5_ASAP7_75t_L g605 ( .A1(n_580), .A2(n_571), .B(n_566), .C(n_576), .Y(n_605) );
OAI21x1_ASAP7_75t_SL g606 ( .A1(n_583), .A2(n_562), .B(n_563), .Y(n_606) );
XNOR2x1_ASAP7_75t_L g607 ( .A(n_591), .B(n_512), .Y(n_607) );
NOR2x1_ASAP7_75t_L g608 ( .A(n_589), .B(n_567), .Y(n_608) );
AO22x2_ASAP7_75t_L g609 ( .A1(n_580), .A2(n_584), .B1(n_586), .B2(n_597), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_582), .A2(n_577), .B1(n_573), .B2(n_564), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_581), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_602), .A2(n_588), .B(n_584), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_605), .B(n_598), .Y(n_613) );
NOR5xp2_ASAP7_75t_SL g614 ( .A(n_600), .B(n_590), .C(n_598), .D(n_585), .E(n_594), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_603), .Y(n_615) );
AOI321xp33_ASAP7_75t_L g616 ( .A1(n_608), .A2(n_592), .A3(n_596), .B1(n_599), .B2(n_540), .C(n_535), .Y(n_616) );
AOI222xp33_ASAP7_75t_L g617 ( .A1(n_601), .A2(n_516), .B1(n_519), .B2(n_513), .C1(n_452), .C2(n_474), .Y(n_617) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_609), .A2(n_519), .B(n_524), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_612), .A2(n_607), .B1(n_609), .B2(n_604), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g620 ( .A(n_613), .B(n_611), .C(n_492), .Y(n_620) );
NAND5xp2_ASAP7_75t_L g621 ( .A(n_616), .B(n_610), .C(n_606), .D(n_464), .E(n_462), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_617), .B(n_452), .C(n_464), .Y(n_622) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_619), .B(n_618), .C(n_614), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_620), .B(n_615), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_623), .A2(n_621), .B(n_622), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_624), .Y(n_626) );
OAI21xp5_ASAP7_75t_L g627 ( .A1(n_625), .A2(n_465), .B(n_461), .Y(n_627) );
AOI221x1_ASAP7_75t_L g628 ( .A1(n_627), .A2(n_626), .B1(n_465), .B2(n_461), .C(n_457), .Y(n_628) );
AOI21xp33_ASAP7_75t_L g629 ( .A1(n_628), .A2(n_457), .B(n_461), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_629), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_630), .A2(n_457), .B(n_470), .Y(n_631) );
endmodule