module fake_jpeg_23668_n_100 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx10_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

AND2x6_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_26),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_16),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_25),
.A2(n_18),
.B1(n_9),
.B2(n_10),
.Y(n_48)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_1),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_32),
.C(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_29),
.Y(n_35)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_2),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_17),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_27),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_17),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_15),
.C(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_5),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_8),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_18),
.B1(n_27),
.B2(n_31),
.Y(n_60)
);

BUFx24_ASAP7_75t_SL g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_63),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_58),
.C(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_60),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_24),
.B(n_11),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_9),
.B(n_11),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_51),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_74),
.B(n_12),
.C(n_40),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_61),
.B1(n_30),
.B2(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_29),
.A3(n_12),
.B1(n_30),
.B2(n_31),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_68),
.C(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_86),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_64),
.B(n_59),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_82),
.B(n_79),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_87),
.B(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_75),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_83),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_90),
.C(n_86),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_95),
.B(n_89),
.Y(n_96)
);

AOI31xp33_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_97),
.A3(n_93),
.B(n_12),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_80),
.B(n_65),
.Y(n_99)
);

AOI221xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_50),
.B1(n_62),
.B2(n_12),
.C(n_40),
.Y(n_100)
);


endmodule