module real_jpeg_30761_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g157 ( 
.A(n_0),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_0),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_0),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_1),
.B(n_488),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_1),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_19),
.B1(n_20),
.B2(n_24),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_2),
.B(n_178),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_2),
.A2(n_19),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_2),
.A2(n_19),
.B1(n_427),
.B2(n_430),
.Y(n_426)
);

INVx3_ASAP7_75t_R g100 ( 
.A(n_3),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_3),
.A2(n_100),
.B1(n_147),
.B2(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_3),
.A2(n_100),
.B1(n_216),
.B2(n_219),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_3),
.B(n_29),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_3),
.B(n_358),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_3),
.B(n_368),
.C(n_371),
.Y(n_367)
);

NAND2xp67_ASAP7_75t_L g383 ( 
.A(n_3),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_3),
.B(n_201),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_5),
.Y(n_94)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_6),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_6),
.Y(n_130)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_6),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_6),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_7),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_7),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_8),
.Y(n_279)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_9),
.Y(n_128)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_9),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_9),
.Y(n_139)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_10),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_10),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_10),
.Y(n_440)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_11),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_12),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_12),
.A2(n_46),
.B1(n_162),
.B2(n_166),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_12),
.A2(n_46),
.B1(n_194),
.B2(n_198),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g435 ( 
.A1(n_12),
.A2(n_46),
.B1(n_436),
.B2(n_438),
.Y(n_435)
);

OAI311xp33_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_65),
.A3(n_487),
.B1(n_489),
.C1(n_494),
.Y(n_13)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_14),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_63),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_62),
.Y(n_15)
);

OR2x6_ASAP7_75t_SL g64 ( 
.A(n_16),
.B(n_62),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_16),
.B(n_486),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_17),
.B(n_458),
.Y(n_457)
);

OA22x2_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_28),
.B1(n_42),
.B2(n_49),
.Y(n_17)
);

AO21x1_ASAP7_75t_L g62 ( 
.A1(n_18),
.A2(n_28),
.B(n_49),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g171 ( 
.A1(n_19),
.A2(n_172),
.B(n_177),
.Y(n_171)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_28),
.A2(n_42),
.B1(n_49),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_50),
.Y(n_49)
);

OAI21x1_ASAP7_75t_L g107 ( 
.A1(n_29),
.A2(n_51),
.B(n_108),
.Y(n_107)
);

OAI22x1_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_32),
.Y(n_267)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_36),
.Y(n_284)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_39),
.Y(n_437)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2x1_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_61),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_L g494 ( 
.A(n_65),
.B(n_495),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_414),
.B(n_480),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_401),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_313),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_286),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_250),
.Y(n_69)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_70),
.Y(n_403)
);

NAND2x1p5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_227),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_71),
.B(n_227),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_181),
.C(n_207),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_73),
.B(n_181),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_118),
.B1(n_179),
.B2(n_180),
.Y(n_73)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_74),
.B(n_213),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_74),
.A2(n_179),
.B1(n_258),
.B2(n_290),
.Y(n_289)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_107),
.B1(n_116),
.B2(n_117),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_75),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_75),
.B(n_117),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_75),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_75),
.B(n_119),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_86),
.B(n_99),
.Y(n_75)
);

NOR2x1p5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_87),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_76),
.Y(n_358)
);

OAI22x1_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_79),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_79),
.Y(n_336)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_81),
.Y(n_197)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_85),
.Y(n_238)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_85),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g433 ( 
.A(n_86),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_86),
.A2(n_99),
.B1(n_358),
.B2(n_435),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B1(n_95),
.B2(n_96),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_90),
.Y(n_432)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_98),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_105),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_109),
.B(n_112),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_104),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_105),
.Y(n_342)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_107),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_108),
.Y(n_454)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_112),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_117),
.Y(n_249)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_118),
.A2(n_208),
.B(n_224),
.Y(n_242)
);

NAND2x1p5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_153),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_119),
.B(n_214),
.Y(n_213)
);

XOR2x2_ASAP7_75t_SL g256 ( 
.A(n_119),
.B(n_153),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_119),
.A2(n_214),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_119),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_119),
.B(n_209),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_119),
.B(n_211),
.Y(n_307)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_119),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_119),
.A2(n_259),
.B1(n_260),
.B2(n_292),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_119),
.A2(n_292),
.B1(n_362),
.B2(n_363),
.Y(n_391)
);

OA21x2_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_135),
.B(n_150),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_121),
.B(n_135),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_125),
.B1(n_129),
.B2(n_131),
.Y(n_121)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_128),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22x1_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_140),
.B1(n_144),
.B2(n_147),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_143),
.Y(n_327)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_148),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_150),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_161),
.B1(n_168),
.B2(n_170),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_154),
.A2(n_161),
.B1(n_215),
.B2(n_220),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx4f_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2x1_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_191),
.B1(n_192),
.B2(n_206),
.Y(n_181)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_182),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_182),
.A2(n_306),
.B1(n_442),
.B2(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OR2x6_ASAP7_75t_L g260 ( 
.A(n_184),
.B(n_215),
.Y(n_260)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_190),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_189),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_201),
.B(n_203),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_193),
.A2(n_201),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_193),
.B(n_201),
.Y(n_246)
);

INVx3_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g423 ( 
.A1(n_201),
.A2(n_233),
.B(n_234),
.Y(n_423)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

NOR2xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

AOI22x1_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_209),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_212),
.B(n_224),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_208),
.A2(n_226),
.B(n_258),
.Y(n_257)
);

NOR2x1p5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_209),
.Y(n_306)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_209),
.Y(n_443)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_232),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_214),
.Y(n_293)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AND3x1_ASAP7_75t_L g295 ( 
.A(n_226),
.B(n_296),
.C(n_297),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_241),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_229),
.B(n_243),
.C(n_479),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B(n_239),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_230),
.B(n_259),
.C(n_311),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_230),
.A2(n_317),
.B(n_319),
.C(n_343),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_230),
.B(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_239),
.B(n_465),
.C(n_470),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_239),
.A2(n_240),
.B1(n_466),
.B2(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_242),
.Y(n_479)
);

XOR2x1_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_244),
.Y(n_471)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_250),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_251),
.B(n_253),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.C(n_257),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_255),
.B(n_256),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_262),
.Y(n_308)
);

NAND2x1p5_ASAP7_75t_L g347 ( 
.A(n_259),
.B(n_320),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_259),
.A2(n_260),
.B1(n_311),
.B2(n_312),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_259),
.B(n_348),
.C(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_259),
.B(n_391),
.Y(n_390)
);

CKINVDCx11_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_260),
.B(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_260),
.B(n_382),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_260),
.B(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OA21x2_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_271),
.B(n_276),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx4f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_270),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_280),
.B(n_285),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx2_ASAP7_75t_SL g281 ( 
.A(n_282),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_300),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_287),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_298),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_288),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.C(n_294),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_294),
.B1(n_295),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_292),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_295),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_296),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g407 ( 
.A(n_298),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_304),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_301),
.B(n_304),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_308),
.C(n_309),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_305),
.B(n_399),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_306),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_306),
.B(n_446),
.C(n_447),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_319),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_308),
.B(n_310),
.Y(n_399)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

OAI21x1_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_396),
.B(n_400),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_353),
.B(n_395),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_344),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_316),
.B(n_344),
.Y(n_395)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_318),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_318),
.B(n_347),
.C(n_349),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_324),
.B(n_332),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_337),
.B(n_341),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_340),
.Y(n_366)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_349),
.B1(n_350),
.B2(n_352),
.Y(n_344)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_345),
.Y(n_352)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

OAI21x1_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_359),
.B(n_394),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_355),
.B(n_356),
.Y(n_394)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_357),
.Y(n_378)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_379),
.B(n_392),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_375),
.Y(n_360)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_390),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_388),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_385),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NOR2x1_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_397),
.B(n_398),
.Y(n_400)
);

AOI21x1_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_405),
.B(n_411),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g411 ( 
.A1(n_403),
.A2(n_412),
.B(n_413),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_461),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_415),
.A2(n_481),
.B(n_485),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_457),
.Y(n_415)
);

NOR2x1_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_449),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_417),
.B(n_449),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_443),
.C(n_444),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_420),
.B(n_442),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_422),
.B1(n_441),
.B2(n_442),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_423),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_423),
.A2(n_446),
.B1(n_448),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_424),
.Y(n_456)
);

OA22x2_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_433),
.B2(n_434),
.Y(n_424)
);

AO21x1_ASAP7_75t_L g451 ( 
.A1(n_425),
.A2(n_426),
.B(n_433),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx8_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_447),
.C(n_456),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_442),
.A2(n_443),
.B1(n_467),
.B2(n_468),
.Y(n_466)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_445),
.B(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_446),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_450),
.B(n_455),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_451),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_452),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_455),
.B(n_459),
.C(n_460),
.Y(n_458)
);

INVxp33_ASAP7_75t_SL g486 ( 
.A(n_458),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_474),
.Y(n_461)
);

OAI211xp5_ASAP7_75t_SL g481 ( 
.A1(n_462),
.A2(n_482),
.B(n_483),
.C(n_484),
.Y(n_481)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_472),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_472),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_466),
.Y(n_477)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_470),
.B(n_476),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_478),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_475),
.B(n_478),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_487),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_487),
.B(n_496),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_492),
.Y(n_491)
);

INVx6_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);


endmodule