module real_jpeg_19068_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_167;
wire n_128;
wire n_179;
wire n_244;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_0),
.A2(n_64),
.B1(n_70),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_0),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_0),
.A2(n_52),
.B1(n_54),
.B2(n_75),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_75),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_0),
.A2(n_27),
.B1(n_29),
.B2(n_75),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_1),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_64),
.B1(n_70),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_2),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_2),
.A2(n_52),
.B1(n_54),
.B2(n_94),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_94),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_94),
.Y(n_226)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_3),
.A2(n_52),
.B1(n_54),
.B2(n_66),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_5),
.A2(n_38),
.B1(n_52),
.B2(n_54),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_38),
.Y(n_146)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_6),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_6),
.B(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_6),
.A2(n_237),
.B(n_261),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_7),
.A2(n_64),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_7),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_7),
.A2(n_52),
.B1(n_54),
.B2(n_71),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_71),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_71),
.Y(n_251)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_9),
.A2(n_27),
.B1(n_29),
.B2(n_46),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_9),
.A2(n_46),
.B1(n_52),
.B2(n_54),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_53),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_10),
.A2(n_53),
.B1(n_64),
.B2(n_70),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_53),
.Y(n_194)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_11),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_11),
.A2(n_52),
.B(n_144),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_11),
.A2(n_64),
.B1(n_70),
.B2(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_11),
.B(n_73),
.Y(n_191)
);

A2O1A1O1Ixp25_ASAP7_75t_L g203 ( 
.A1(n_11),
.A2(n_35),
.B(n_40),
.C(n_204),
.D(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_11),
.B(n_35),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_11),
.B(n_58),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_11),
.A2(n_25),
.B(n_219),
.Y(n_239)
);

A2O1A1O1Ixp25_ASAP7_75t_L g252 ( 
.A1(n_11),
.A2(n_54),
.B(n_55),
.C(n_152),
.D(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_11),
.B(n_54),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_14),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_110)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_16),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_20),
.B(n_102),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.C(n_82),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_21),
.A2(n_22),
.B1(n_76),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_23),
.B(n_50),
.C(n_61),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_24),
.B(n_33),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_25),
.A2(n_26),
.B(n_31),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_25),
.A2(n_28),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_25),
.A2(n_85),
.B1(n_88),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_25),
.A2(n_26),
.B1(n_146),
.B2(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_25),
.A2(n_218),
.B(n_219),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_25),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_25),
.B(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_26),
.Y(n_229)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_29),
.B1(n_41),
.B2(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_27),
.A2(n_42),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_29),
.B(n_41),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_29),
.B(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_45),
.B2(n_47),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_34),
.A2(n_39),
.B1(n_47),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_36),
.B1(n_56),
.B2(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_35),
.A2(n_253),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_41),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_36),
.B(n_59),
.Y(n_258)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_39),
.A2(n_45),
.B1(n_47),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_39),
.A2(n_47),
.B1(n_216),
.B2(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_39),
.A2(n_251),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_40),
.A2(n_43),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_40),
.B(n_168),
.Y(n_167)
);

CKINVDCx9p33_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_47),
.A2(n_90),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_47),
.B(n_169),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_47),
.A2(n_167),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_47),
.B(n_142),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_61),
.B2(n_62),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B1(n_58),
.B2(n_60),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_51),
.Y(n_97)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_56),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_55),
.A2(n_58),
.B1(n_60),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_55),
.Y(n_150)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_57),
.Y(n_259)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_69),
.B(n_72),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_68),
.B1(n_69),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_66),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_64),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_64),
.A2(n_66),
.B(n_142),
.C(n_143),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_68),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_68),
.A2(n_93),
.B(n_122),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_72),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_78),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_79),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_80),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_82),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_91),
.C(n_95),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_84),
.B(n_89),
.Y(n_163)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_88),
.A2(n_226),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_88),
.B(n_142),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B(n_99),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_101),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_98),
.A2(n_149),
.B1(n_150),
.B2(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_98),
.A2(n_99),
.B(n_175),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_125),
.B2(n_126),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_114),
.B2(n_115),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_111),
.B(n_113),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_111),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_124),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_125),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_156),
.B(n_284),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_153),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_131),
.B(n_153),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_135),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_134),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_136),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.C(n_147),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_138),
.B1(n_147),
.B2(n_148),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_145),
.Y(n_139)
);

AOI22x1_ASAP7_75t_SL g185 ( 
.A1(n_140),
.A2(n_141),
.B1(n_145),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_145),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B(n_151),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_196),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_179),
.B(n_195),
.Y(n_158)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_159),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_176),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_176),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.C(n_164),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_164),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.C(n_173),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_166),
.B1(n_173),
.B2(n_174),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_180),
.B(n_182),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.C(n_187),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_183),
.B(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_185),
.A2(n_187),
.B1(n_188),
.B2(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_185),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.C(n_192),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_189),
.A2(n_190),
.B1(n_268),
.B2(n_270),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_191),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_194),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_282),
.C(n_283),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_276),
.B(n_281),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_264),
.B(n_275),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_245),
.B(n_263),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_222),
.B(n_244),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_210),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_202),
.B(n_210),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_203),
.A2(n_206),
.B1(n_207),
.B2(n_231),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_217),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_215),
.C(n_217),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_218),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_232),
.B(n_243),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_230),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_230),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_238),
.B(n_242),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_234),
.B(n_235),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_246),
.B(n_247),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_256),
.B2(n_262),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_252),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_255),
.C(n_262),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_256),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_260),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_272),
.C(n_273),
.Y(n_277)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);


endmodule