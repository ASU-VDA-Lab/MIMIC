module fake_jpeg_28398_n_293 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_20),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_32),
.Y(n_47)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_28),
.B1(n_16),
.B2(n_4),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_1),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_29),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_23),
.B1(n_17),
.B2(n_25),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_43),
.A2(n_39),
.B1(n_49),
.B2(n_44),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_25),
.B1(n_21),
.B2(n_17),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_45),
.A2(n_31),
.B1(n_5),
.B2(n_6),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_61),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_26),
.C(n_32),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_18),
.C(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_35),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_13),
.B(n_15),
.Y(n_78)
);

FAx1_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_40),
.CI(n_39),
.CON(n_62),
.SN(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_95),
.B(n_4),
.C(n_57),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_92),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_65),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_67),
.B(n_9),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_70),
.B(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_36),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_77),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_41),
.B1(n_37),
.B2(n_38),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_78),
.B1(n_80),
.B2(n_87),
.Y(n_97)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_37),
.Y(n_77)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

OA22x2_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_39),
.B1(n_35),
.B2(n_16),
.Y(n_85)
);

AO22x2_ASAP7_75t_L g114 ( 
.A1(n_85),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_114)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_33),
.B1(n_24),
.B2(n_29),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_14),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_60),
.A2(n_33),
.B1(n_24),
.B2(n_16),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_94),
.B1(n_4),
.B2(n_7),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_2),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_2),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_7),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_19),
.B1(n_31),
.B2(n_3),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_3),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_88),
.B1(n_62),
.B2(n_89),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_99),
.B(n_120),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_31),
.B(n_5),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_100),
.A2(n_105),
.B(n_95),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_114),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_112),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_8),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_68),
.A2(n_15),
.B(n_10),
.C(n_11),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_78),
.B(n_70),
.Y(n_131)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_117),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_9),
.Y(n_120)
);

BUFx24_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_11),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_74),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_125),
.B(n_132),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_62),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_126),
.B(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_129),
.B(n_133),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_68),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_131),
.B(n_152),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_74),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_64),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_68),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_64),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_106),
.C(n_112),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_149),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_63),
.B1(n_76),
.B2(n_85),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_97),
.B1(n_113),
.B2(n_107),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_90),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_114),
.Y(n_146)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_147),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_71),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_93),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_119),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_92),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_105),
.B(n_113),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_156),
.A2(n_146),
.B(n_148),
.Y(n_185)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_170),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_127),
.B1(n_126),
.B2(n_142),
.Y(n_193)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_174),
.B(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_95),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_182),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_115),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_141),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_109),
.Y(n_184)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_185),
.A2(n_186),
.B(n_189),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_156),
.A2(n_131),
.B(n_127),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_138),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_196),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_167),
.A2(n_184),
.B(n_160),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_207),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_145),
.B1(n_139),
.B2(n_152),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_193),
.A2(n_164),
.B1(n_165),
.B2(n_169),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_127),
.B(n_142),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_198),
.B(n_200),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_141),
.C(n_150),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_206),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_85),
.B(n_91),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_166),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_155),
.A2(n_89),
.B1(n_86),
.B2(n_73),
.Y(n_205)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_104),
.C(n_123),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_169),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_183),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_158),
.Y(n_211)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_221),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_157),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_162),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_161),
.B1(n_159),
.B2(n_171),
.Y(n_220)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_224),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_204),
.A2(n_171),
.B1(n_157),
.B2(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_227),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_194),
.A2(n_163),
.B1(n_180),
.B2(n_175),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_188),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_222),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_224),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_197),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_234),
.Y(n_250)
);

AOI21xp33_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_186),
.B(n_189),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_233),
.A2(n_185),
.B(n_236),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_162),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_213),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_196),
.C(n_190),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_242),
.C(n_229),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_226),
.A2(n_190),
.B1(n_195),
.B2(n_198),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_214),
.B1(n_220),
.B2(n_200),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_195),
.C(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_178),
.Y(n_268)
);

OAI22x1_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_213),
.B1(n_227),
.B2(n_200),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_248),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_240),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_253),
.C(n_238),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_226),
.B1(n_212),
.B2(n_180),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_191),
.B1(n_202),
.B2(n_174),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_228),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_258),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_257),
.A2(n_245),
.B(n_181),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_170),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_263),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_237),
.C(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_264),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_236),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_237),
.C(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_179),
.C(n_178),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_66),
.Y(n_277)
);

O2A1O1Ixp33_ASAP7_75t_SL g274 ( 
.A1(n_268),
.A2(n_104),
.B(n_123),
.C(n_12),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_268),
.A2(n_247),
.B1(n_248),
.B2(n_250),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_273),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_11),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_271),
.A2(n_277),
.B(n_12),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_265),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_274),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_264),
.Y(n_278)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_272),
.B(n_269),
.Y(n_280)
);

AOI21x1_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_271),
.B(n_273),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_283),
.C(n_279),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_262),
.C(n_261),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_261),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_285),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_290),
.A2(n_289),
.B1(n_286),
.B2(n_66),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_13),
.C(n_104),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_13),
.Y(n_293)
);


endmodule