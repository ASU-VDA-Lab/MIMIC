module fake_netlist_1_12194_n_37 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_0), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
BUFx10_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_3), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_0), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_13), .B(n_1), .C(n_2), .Y(n_20) );
INVx3_ASAP7_75t_L g21 ( .A(n_12), .Y(n_21) );
NOR3xp33_ASAP7_75t_SL g22 ( .A(n_15), .B(n_2), .C(n_3), .Y(n_22) );
OR2x6_ASAP7_75t_L g23 ( .A(n_22), .B(n_16), .Y(n_23) );
NAND3xp33_ASAP7_75t_L g24 ( .A(n_20), .B(n_12), .C(n_14), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_21), .A2(n_18), .B1(n_17), .B2(n_12), .Y(n_25) );
OAI31xp33_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_21), .A3(n_15), .B(n_18), .Y(n_26) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
INVxp67_ASAP7_75t_SL g28 ( .A(n_27), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
NAND2xp5_ASAP7_75t_SL g30 ( .A(n_28), .B(n_26), .Y(n_30) );
NOR3xp33_ASAP7_75t_SL g31 ( .A(n_29), .B(n_23), .C(n_6), .Y(n_31) );
AOI21xp33_ASAP7_75t_SL g32 ( .A1(n_30), .A2(n_29), .B(n_6), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g33 ( .A(n_31), .B(n_4), .Y(n_33) );
NOR3xp33_ASAP7_75t_SL g34 ( .A(n_33), .B(n_7), .C(n_8), .Y(n_34) );
NAND5xp2_ASAP7_75t_L g35 ( .A(n_32), .B(n_7), .C(n_9), .D(n_10), .E(n_11), .Y(n_35) );
BUFx2_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
NAND3xp33_ASAP7_75t_L g37 ( .A(n_36), .B(n_19), .C(n_35), .Y(n_37) );
endmodule