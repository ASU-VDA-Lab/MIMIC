module fake_netlist_1_7487_n_15 (n_1, n_2, n_0, n_15);
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_10;
wire n_8;
NAND2xp5_ASAP7_75t_SL g3 ( .A(n_1), .B(n_2), .Y(n_3) );
BUFx3_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
AND2x2_ASAP7_75t_L g5 ( .A(n_0), .B(n_2), .Y(n_5) );
INVx1_ASAP7_75t_SL g6 ( .A(n_5), .Y(n_6) );
AOI21x1_ASAP7_75t_L g7 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_4), .Y(n_8) );
OR2x2_ASAP7_75t_L g9 ( .A(n_7), .B(n_4), .Y(n_9) );
NAND2xp5_ASAP7_75t_SL g10 ( .A(n_8), .B(n_7), .Y(n_10) );
OR3x2_ASAP7_75t_L g11 ( .A(n_9), .B(n_0), .C(n_5), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
AOI22xp5_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_13), .B1(n_11), .B2(n_8), .Y(n_15) );
endmodule