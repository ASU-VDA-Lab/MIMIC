module fake_jpeg_11559_n_96 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_96);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_10),
.Y(n_11)
);

INVx2_ASAP7_75t_SL g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_29),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_1),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_12),
.B1(n_19),
.B2(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_30),
.B1(n_13),
.B2(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_15),
.B1(n_16),
.B2(n_12),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_27),
.B1(n_12),
.B2(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_26),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_52),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_45),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_27),
.C(n_29),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_38),
.C(n_36),
.Y(n_55)
);

XNOR2x1_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_49),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_21),
.B1(n_17),
.B2(n_19),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_21),
.B1(n_17),
.B2(n_18),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_16),
.C(n_37),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_37),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_14),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_38),
.B(n_13),
.C(n_34),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_62),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_63),
.C(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_20),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_20),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_63),
.B(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_65),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_69),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_52),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_59),
.B1(n_62),
.B2(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_54),
.B(n_53),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_68),
.B(n_67),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_59),
.B1(n_54),
.B2(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_78),
.Y(n_81)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_82),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_67),
.B(n_47),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_67),
.B(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_77),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_88),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_75),
.B1(n_74),
.B2(n_20),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_10),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_5),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_88),
.C(n_7),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_89),
.B1(n_93),
.B2(n_9),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_9),
.Y(n_96)
);


endmodule