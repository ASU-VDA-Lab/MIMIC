module fake_jpeg_21258_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

OR2x2_ASAP7_75t_SL g13 ( 
.A(n_0),
.B(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_15),
.A2(n_21),
.B1(n_22),
.B2(n_10),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_16),
.A2(n_14),
.B1(n_7),
.B2(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_10),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_9),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_12),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_31),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_10),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_18),
.Y(n_38)
);

A2O1A1O1Ixp25_ASAP7_75t_L g30 ( 
.A1(n_16),
.A2(n_11),
.B(n_21),
.C(n_22),
.D(n_17),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_11),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_20),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_29),
.C(n_36),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_29),
.B1(n_24),
.B2(n_20),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_SL g39 ( 
.A(n_37),
.B(n_25),
.C(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_42),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_35),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_47),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_42),
.C(n_44),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_49),
.Y(n_51)
);


endmodule