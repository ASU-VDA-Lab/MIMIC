module fake_netlist_1_8108_n_728 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_728);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_728;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_721;
wire n_438;
wire n_134;
wire n_656;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_50), .Y(n_82) );
INVxp67_ASAP7_75t_L g83 ( .A(n_27), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_16), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_59), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_78), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_38), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_75), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_32), .Y(n_89) );
BUFx2_ASAP7_75t_L g90 ( .A(n_79), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_68), .Y(n_91) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_25), .Y(n_92) );
INVx2_ASAP7_75t_SL g93 ( .A(n_2), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_10), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_23), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_42), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_70), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_39), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_29), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_54), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_43), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_3), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_80), .Y(n_103) );
CKINVDCx14_ASAP7_75t_R g104 ( .A(n_72), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_44), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_4), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_52), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_74), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_62), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_3), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_67), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_53), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_19), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_1), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_66), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_4), .Y(n_116) );
INVxp33_ASAP7_75t_L g117 ( .A(n_28), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_25), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_56), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_46), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_10), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_12), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_37), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_14), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_36), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_13), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_33), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_71), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_8), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_22), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_24), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_121), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_121), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_90), .B(n_0), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_90), .B(n_0), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_121), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_86), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_124), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_124), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_105), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_124), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_105), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_85), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_84), .B(n_1), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_93), .B(n_102), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_105), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_84), .B(n_2), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_85), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_89), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_89), .Y(n_152) );
CKINVDCx6p67_ASAP7_75t_R g153 ( .A(n_108), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_106), .B(n_5), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_91), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_91), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_96), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_93), .B(n_5), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_93), .B(n_6), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_96), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_106), .B(n_6), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_107), .B(n_7), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_107), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_107), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_97), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_102), .B(n_7), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_94), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_92), .Y(n_168) );
NAND2x1_ASAP7_75t_L g169 ( .A(n_97), .B(n_8), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_98), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_98), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_99), .Y(n_172) );
INVx1_ASAP7_75t_SL g173 ( .A(n_108), .Y(n_173) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_110), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_92), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_115), .B(n_9), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_162), .Y(n_177) );
BUFx10_ASAP7_75t_L g178 ( .A(n_167), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_153), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_147), .B(n_111), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_162), .Y(n_181) );
OR2x6_ASAP7_75t_L g182 ( .A(n_146), .B(n_114), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_153), .Y(n_183) );
INVx1_ASAP7_75t_SL g184 ( .A(n_173), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_132), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_162), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_162), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_162), .Y(n_188) );
INVx4_ASAP7_75t_SL g189 ( .A(n_136), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_173), .B(n_115), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_132), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_153), .B(n_119), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_132), .Y(n_193) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_167), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_174), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_158), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_147), .B(n_117), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_136), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_170), .B(n_99), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_136), .B(n_114), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_158), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_137), .B(n_119), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_170), .B(n_101), .Y(n_203) );
INVx4_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
NAND2x1p5_ASAP7_75t_L g206 ( .A(n_137), .B(n_116), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_145), .B(n_104), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_174), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_132), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_146), .B(n_116), .Y(n_210) );
BUFx4f_ASAP7_75t_L g211 ( .A(n_145), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_150), .B(n_83), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_176), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_132), .Y(n_214) );
NOR2x1p5_ASAP7_75t_L g215 ( .A(n_169), .B(n_146), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_150), .B(n_83), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_151), .B(n_131), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_149), .A2(n_95), .B1(n_130), .B2(n_131), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_151), .B(n_120), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_152), .B(n_130), .Y(n_220) );
AND2x6_ASAP7_75t_L g221 ( .A(n_176), .B(n_103), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_149), .A2(n_122), .B1(n_126), .B2(n_118), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_132), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_132), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_163), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_132), .Y(n_226) );
INVxp67_ASAP7_75t_L g227 ( .A(n_176), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_149), .B(n_122), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_154), .Y(n_229) );
NAND3xp33_ASAP7_75t_L g230 ( .A(n_159), .B(n_126), .C(n_113), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_152), .B(n_87), .Y(n_231) );
AOI21x1_ASAP7_75t_L g232 ( .A1(n_170), .A2(n_120), .B(n_128), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_170), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_155), .B(n_112), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_165), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_154), .B(n_161), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_154), .B(n_92), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_155), .B(n_112), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_156), .B(n_123), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_156), .B(n_123), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_165), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_165), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_161), .B(n_92), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_194), .B(n_161), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_221), .A2(n_82), .B1(n_169), .B2(n_171), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_196), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_201), .A2(n_157), .B1(n_171), .B2(n_160), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_180), .B(n_157), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_205), .A2(n_160), .B1(n_172), .B2(n_163), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_225), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_237), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_180), .B(n_172), .Y(n_252) );
CKINVDCx16_ASAP7_75t_R g253 ( .A(n_178), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_197), .B(n_172), .Y(n_254) );
OR2x6_ASAP7_75t_L g255 ( .A(n_182), .B(n_169), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_225), .Y(n_256) );
OR2x2_ASAP7_75t_SL g257 ( .A(n_194), .B(n_129), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_197), .B(n_166), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_195), .B(n_166), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_184), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_198), .B(n_163), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_211), .B(n_142), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_198), .B(n_163), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_204), .B(n_163), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_204), .B(n_109), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_221), .A2(n_109), .B1(n_100), .B2(n_88), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_178), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_207), .B(n_138), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_206), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_183), .B(n_134), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_206), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_177), .A2(n_135), .B1(n_139), .B2(n_164), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_202), .B(n_138), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_243), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_237), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_200), .B(n_140), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_189), .B(n_134), .Y(n_277) );
INVx4_ASAP7_75t_L g278 ( .A(n_189), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_181), .A2(n_139), .B(n_135), .C(n_164), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_237), .Y(n_280) );
OR2x6_ASAP7_75t_L g281 ( .A(n_182), .B(n_92), .Y(n_281) );
CKINVDCx14_ASAP7_75t_R g282 ( .A(n_179), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_185), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_233), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_195), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_208), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_185), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_211), .A2(n_139), .B(n_135), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_185), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_185), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_208), .Y(n_291) );
CKINVDCx6p67_ASAP7_75t_R g292 ( .A(n_182), .Y(n_292) );
INVx5_ASAP7_75t_L g293 ( .A(n_221), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_200), .B(n_101), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_213), .A2(n_164), .B(n_144), .C(n_140), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_221), .Y(n_296) );
BUFx8_ASAP7_75t_L g297 ( .A(n_229), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_186), .B(n_148), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_217), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_221), .A2(n_128), .B1(n_103), .B2(n_125), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_217), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_213), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_236), .B(n_141), .Y(n_303) );
INVx5_ASAP7_75t_L g304 ( .A(n_214), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_231), .B(n_212), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_227), .A2(n_125), .B1(n_127), .B2(n_144), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_228), .B(n_133), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_218), .A2(n_144), .B1(n_143), .B2(n_133), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_217), .Y(n_309) );
INVxp67_ASAP7_75t_SL g310 ( .A(n_187), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_216), .B(n_143), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_188), .B(n_148), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_220), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_220), .B(n_148), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_235), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_246), .A2(n_220), .B1(n_215), .B2(n_228), .Y(n_316) );
OR2x6_ASAP7_75t_L g317 ( .A(n_281), .B(n_192), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_285), .A2(n_190), .B1(n_222), .B2(n_210), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_278), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_281), .B(n_260), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_299), .Y(n_322) );
AND2x4_ASAP7_75t_SL g323 ( .A(n_292), .B(n_189), .Y(n_323) );
NOR2xp67_ASAP7_75t_SL g324 ( .A(n_293), .B(n_240), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_305), .A2(n_238), .B(n_199), .Y(n_325) );
AND2x6_ASAP7_75t_L g326 ( .A(n_296), .B(n_241), .Y(n_326) );
OAI22xp33_ASAP7_75t_L g327 ( .A1(n_281), .A2(n_141), .B1(n_230), .B2(n_242), .Y(n_327) );
INVx3_ASAP7_75t_SL g328 ( .A(n_253), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_259), .B(n_239), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_296), .A2(n_239), .B1(n_234), .B2(n_219), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_297), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_258), .B(n_234), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_251), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_269), .B(n_238), .Y(n_334) );
A2O1A1Ixp33_ASAP7_75t_L g335 ( .A1(n_279), .A2(n_219), .B(n_199), .C(n_203), .Y(n_335) );
CKINVDCx11_ASAP7_75t_R g336 ( .A(n_267), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_293), .B(n_232), .Y(n_337) );
BUFx12f_ASAP7_75t_L g338 ( .A(n_297), .Y(n_338) );
BUFx4_ASAP7_75t_SL g339 ( .A(n_286), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_271), .B(n_203), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_310), .A2(n_92), .B1(n_113), .B2(n_127), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_278), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_293), .B(n_113), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_293), .B(n_113), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_251), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_315), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_248), .B(n_113), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_301), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_310), .A2(n_113), .B1(n_142), .B2(n_148), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_298), .A2(n_193), .B(n_224), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_265), .B(n_9), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_247), .B(n_142), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_309), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_244), .B(n_11), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_291), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_270), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_265), .B(n_11), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_277), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_313), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_302), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_277), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_283), .Y(n_362) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_283), .Y(n_363) );
INVx5_ASAP7_75t_L g364 ( .A(n_255), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_266), .B(n_12), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_283), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_303), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_274), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_270), .B(n_13), .Y(n_369) );
NOR2xp67_ASAP7_75t_L g370 ( .A(n_245), .B(n_14), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_275), .A2(n_142), .B1(n_148), .B2(n_193), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g372 ( .A1(n_360), .A2(n_255), .B1(n_300), .B2(n_254), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_346), .Y(n_373) );
INVx6_ASAP7_75t_L g374 ( .A(n_342), .Y(n_374) );
INVx4_ASAP7_75t_L g375 ( .A(n_326), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_346), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_362), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_348), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_328), .B(n_257), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_351), .A2(n_255), .B1(n_274), .B2(n_280), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g381 ( .A1(n_355), .A2(n_252), .B1(n_307), .B2(n_273), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_367), .A2(n_294), .B1(n_308), .B2(n_276), .C(n_295), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_351), .A2(n_294), .B1(n_247), .B2(n_282), .Y(n_384) );
OA21x2_ASAP7_75t_L g385 ( .A1(n_335), .A2(n_279), .B(n_288), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_329), .A2(n_249), .B1(n_306), .B2(n_282), .C(n_264), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_319), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_356), .A2(n_249), .B1(n_261), .B2(n_263), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_322), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_342), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_352), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_332), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_357), .A2(n_314), .B1(n_256), .B2(n_250), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_362), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_362), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_316), .A2(n_317), .B1(n_357), .B2(n_369), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_316), .A2(n_272), .B1(n_311), .B2(n_268), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_328), .B(n_272), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_317), .A2(n_314), .B1(n_312), .B2(n_298), .Y(n_400) );
AND2x6_ASAP7_75t_L g401 ( .A(n_321), .B(n_287), .Y(n_401) );
OAI222xp33_ASAP7_75t_L g402 ( .A1(n_364), .A2(n_262), .B1(n_312), .B2(n_168), .C1(n_18), .C2(n_19), .Y(n_402) );
A2O1A1Ixp33_ASAP7_75t_L g403 ( .A1(n_325), .A2(n_262), .B(n_148), .C(n_142), .Y(n_403) );
INVx5_ASAP7_75t_L g404 ( .A(n_326), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_364), .B(n_304), .Y(n_405) );
NOR2x1_ASAP7_75t_SL g406 ( .A(n_317), .B(n_304), .Y(n_406) );
AOI21xp33_ASAP7_75t_L g407 ( .A1(n_397), .A2(n_369), .B(n_347), .Y(n_407) );
OAI21x1_ASAP7_75t_L g408 ( .A1(n_392), .A2(n_337), .B(n_349), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_373), .Y(n_409) );
OAI21xp5_ASAP7_75t_SL g410 ( .A1(n_381), .A2(n_321), .B(n_365), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_372), .B(n_364), .Y(n_411) );
AOI21xp33_ASAP7_75t_L g412 ( .A1(n_392), .A2(n_365), .B(n_368), .Y(n_412) );
OAI21x1_ASAP7_75t_L g413 ( .A1(n_377), .A2(n_337), .B(n_350), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_393), .A2(n_370), .B1(n_354), .B2(n_368), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_375), .B(n_364), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_373), .Y(n_416) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_404), .Y(n_417) );
AO31x2_ASAP7_75t_L g418 ( .A1(n_403), .A2(n_335), .A3(n_330), .B(n_341), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_379), .Y(n_419) );
A2O1A1Ixp33_ASAP7_75t_L g420 ( .A1(n_393), .A2(n_318), .B(n_334), .C(n_340), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_376), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_384), .A2(n_379), .B1(n_399), .B2(n_386), .Y(n_422) );
AOI21xp33_ASAP7_75t_L g423 ( .A1(n_385), .A2(n_327), .B(n_344), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_399), .A2(n_336), .B1(n_331), .B2(n_345), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_401), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_375), .A2(n_338), .B1(n_333), .B2(n_345), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_376), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_378), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_383), .A2(n_336), .B1(n_333), .B2(n_334), .Y(n_429) );
NAND2xp33_ASAP7_75t_SL g430 ( .A(n_375), .B(n_324), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g431 ( .A1(n_398), .A2(n_340), .B(n_323), .C(n_344), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_388), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_380), .A2(n_361), .B1(n_358), .B2(n_323), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_401), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_378), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_382), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_419), .B(n_382), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_409), .Y(n_438) );
NAND4xp25_ASAP7_75t_L g439 ( .A(n_422), .B(n_387), .C(n_394), .D(n_390), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_428), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_409), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_425), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_412), .A2(n_387), .B1(n_390), .B2(n_388), .Y(n_443) );
NOR2x1p5_ASAP7_75t_L g444 ( .A(n_434), .B(n_391), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_432), .B(n_385), .Y(n_445) );
BUFx4f_ASAP7_75t_L g446 ( .A(n_415), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_409), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_412), .A2(n_385), .B1(n_389), .B2(n_401), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_428), .Y(n_449) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_410), .A2(n_385), .B1(n_391), .B2(n_374), .C(n_400), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_435), .B(n_401), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_416), .Y(n_452) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_423), .A2(n_402), .B(n_377), .Y(n_453) );
AOI33xp33_ASAP7_75t_L g454 ( .A1(n_424), .A2(n_339), .A3(n_327), .B1(n_343), .B2(n_209), .B3(n_191), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_416), .B(n_406), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_435), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_425), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_436), .Y(n_458) );
OAI21xp33_ASAP7_75t_SL g459 ( .A1(n_421), .A2(n_396), .B(n_395), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_436), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_434), .B(n_406), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_410), .B(n_358), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_421), .B(n_395), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_427), .Y(n_464) );
OAI321xp33_ASAP7_75t_L g465 ( .A1(n_429), .A2(n_142), .A3(n_148), .B1(n_371), .B2(n_175), .C(n_339), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_427), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_434), .Y(n_467) );
AOI31xp33_ASAP7_75t_L g468 ( .A1(n_411), .A2(n_405), .A3(n_396), .B(n_404), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_413), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_420), .B(n_391), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_414), .B(n_407), .C(n_431), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_418), .B(n_405), .Y(n_472) );
OAI211xp5_ASAP7_75t_L g473 ( .A1(n_433), .A2(n_404), .B(n_361), .C(n_320), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_440), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_438), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_452), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_437), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_452), .B(n_418), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_440), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_446), .A2(n_443), .B1(n_450), .B2(n_462), .Y(n_480) );
BUFx3_ASAP7_75t_L g481 ( .A(n_446), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_449), .B(n_426), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_471), .B(n_142), .C(n_148), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_449), .B(n_407), .Y(n_484) );
NAND4xp25_ASAP7_75t_SL g485 ( .A(n_454), .B(n_423), .C(n_16), .D(n_17), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_456), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_472), .B(n_418), .Y(n_487) );
NOR3xp33_ASAP7_75t_L g488 ( .A(n_439), .B(n_168), .C(n_430), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_438), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_472), .B(n_417), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_445), .B(n_472), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_439), .B(n_168), .C(n_320), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_471), .A2(n_415), .B1(n_401), .B2(n_374), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_446), .A2(n_415), .B1(n_404), .B2(n_374), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_456), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_445), .B(n_418), .Y(n_496) );
OAI31xp33_ASAP7_75t_L g497 ( .A1(n_450), .A2(n_415), .A3(n_405), .B(n_343), .Y(n_497) );
OAI211xp5_ASAP7_75t_L g498 ( .A1(n_443), .A2(n_142), .B(n_168), .C(n_404), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_464), .B(n_418), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_464), .B(n_418), .Y(n_500) );
NAND4xp25_ASAP7_75t_L g501 ( .A(n_448), .B(n_460), .C(n_458), .D(n_470), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_458), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_464), .B(n_408), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_460), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_455), .Y(n_505) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_446), .A2(n_468), .B1(n_465), .B2(n_442), .Y(n_506) );
BUFx3_ASAP7_75t_L g507 ( .A(n_455), .Y(n_507) );
BUFx3_ASAP7_75t_L g508 ( .A(n_455), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_466), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_448), .A2(n_404), .B1(n_374), .B2(n_417), .Y(n_510) );
OAI31xp33_ASAP7_75t_L g511 ( .A1(n_444), .A2(n_405), .A3(n_168), .B(n_209), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_438), .B(n_408), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_444), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_441), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_441), .B(n_408), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_441), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_451), .A2(n_401), .B1(n_326), .B2(n_417), .Y(n_517) );
OAI211xp5_ASAP7_75t_L g518 ( .A1(n_459), .A2(n_175), .B(n_417), .C(n_191), .Y(n_518) );
OAI221xp5_ASAP7_75t_L g519 ( .A1(n_470), .A2(n_417), .B1(n_175), .B2(n_224), .C(n_226), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_463), .B(n_15), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_447), .B(n_417), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_447), .B(n_413), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_461), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_447), .B(n_15), .Y(n_524) );
AOI211xp5_ASAP7_75t_L g525 ( .A1(n_480), .A2(n_465), .B(n_473), .C(n_461), .Y(n_525) );
INVx1_ASAP7_75t_SL g526 ( .A(n_507), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_474), .B(n_463), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_491), .B(n_442), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_505), .B(n_457), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_487), .B(n_469), .Y(n_530) );
NAND3xp33_ASAP7_75t_SL g531 ( .A(n_511), .B(n_473), .C(n_467), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_491), .B(n_457), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_475), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_509), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_507), .B(n_463), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_474), .B(n_451), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_487), .B(n_469), .Y(n_537) );
OAI21xp33_ASAP7_75t_L g538 ( .A1(n_501), .A2(n_459), .B(n_175), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_476), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_508), .B(n_467), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_499), .B(n_500), .Y(n_541) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_477), .B(n_175), .C(n_468), .Y(n_542) );
NOR3xp33_ASAP7_75t_L g543 ( .A(n_485), .B(n_461), .C(n_469), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_508), .B(n_461), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_509), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_479), .B(n_453), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_514), .B(n_453), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_490), .B(n_453), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_524), .B(n_453), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_482), .B(n_17), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_479), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_518), .A2(n_366), .B(n_363), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_514), .B(n_18), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_524), .B(n_20), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_486), .B(n_20), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_486), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_495), .Y(n_557) );
NOR2x1p5_ASAP7_75t_SL g558 ( .A(n_515), .B(n_175), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_506), .A2(n_326), .B1(n_175), .B2(n_223), .Y(n_559) );
AND2x4_ASAP7_75t_SL g560 ( .A(n_513), .B(n_366), .Y(n_560) );
AOI21xp33_ASAP7_75t_SL g561 ( .A1(n_513), .A2(n_21), .B(n_22), .Y(n_561) );
INVx3_ASAP7_75t_L g562 ( .A(n_490), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_499), .B(n_175), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_481), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_490), .B(n_21), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_523), .B(n_63), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_516), .B(n_23), .Y(n_567) );
AND2x4_ASAP7_75t_SL g568 ( .A(n_521), .B(n_366), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_516), .B(n_24), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_495), .B(n_326), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_502), .Y(n_571) );
INVx3_ASAP7_75t_L g572 ( .A(n_475), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_502), .B(n_226), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_489), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_500), .B(n_26), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_489), .B(n_30), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_504), .B(n_31), .Y(n_577) );
NAND3xp33_ASAP7_75t_SL g578 ( .A(n_497), .B(n_34), .C(n_35), .Y(n_578) );
XNOR2x2_ASAP7_75t_L g579 ( .A(n_484), .B(n_40), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_496), .B(n_41), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_520), .Y(n_581) );
INVx3_ASAP7_75t_SL g582 ( .A(n_481), .Y(n_582) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_515), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_541), .B(n_496), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_539), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_541), .B(n_478), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_542), .A2(n_517), .B1(n_494), .B2(n_478), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_539), .B(n_503), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_528), .B(n_503), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_561), .A2(n_488), .B(n_498), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_530), .B(n_512), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_526), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_532), .B(n_521), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_530), .B(n_512), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_534), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_581), .B(n_545), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_537), .B(n_522), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_537), .B(n_522), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_551), .B(n_493), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_556), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_550), .B(n_510), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_557), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_535), .B(n_519), .Y(n_603) );
NAND4xp75_ASAP7_75t_SL g604 ( .A(n_550), .B(n_492), .C(n_483), .D(n_48), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_549), .B(n_226), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_571), .B(n_223), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_582), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_527), .B(n_223), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_555), .B(n_45), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_562), .B(n_214), .Y(n_610) );
INVx2_ASAP7_75t_SL g611 ( .A(n_544), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_563), .B(n_214), .Y(n_612) );
NAND2x1_ASAP7_75t_L g613 ( .A(n_544), .B(n_366), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_562), .B(n_47), .Y(n_614) );
OR2x6_ASAP7_75t_L g615 ( .A(n_544), .B(n_540), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_525), .A2(n_363), .B1(n_362), .B2(n_214), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_562), .B(n_49), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_563), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_583), .B(n_51), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_538), .B(n_363), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_548), .B(n_55), .Y(n_621) );
NAND4xp25_ASAP7_75t_SL g622 ( .A(n_564), .B(n_57), .C(n_58), .D(n_60), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_536), .Y(n_623) );
NAND2x1_ASAP7_75t_SL g624 ( .A(n_582), .B(n_61), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_548), .B(n_64), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_572), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_583), .B(n_65), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_572), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_572), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_529), .B(n_69), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_533), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_574), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_574), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_553), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_567), .Y(n_635) );
AND2x4_ASAP7_75t_SL g636 ( .A(n_565), .B(n_363), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_592), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_584), .B(n_546), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_585), .Y(n_639) );
INVxp67_ASAP7_75t_SL g640 ( .A(n_620), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_584), .B(n_580), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_596), .Y(n_642) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_601), .A2(n_579), .B1(n_580), .B2(n_554), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_601), .B(n_543), .C(n_547), .Y(n_644) );
AOI32xp33_ASAP7_75t_L g645 ( .A1(n_607), .A2(n_543), .A3(n_575), .B1(n_577), .B2(n_548), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_586), .B(n_575), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_586), .B(n_569), .Y(n_647) );
AOI211x1_ASAP7_75t_L g648 ( .A1(n_587), .A2(n_578), .B(n_531), .C(n_570), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_589), .B(n_588), .Y(n_649) );
XNOR2xp5_ASAP7_75t_L g650 ( .A(n_592), .B(n_593), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_623), .B(n_577), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_595), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_634), .B(n_577), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_615), .A2(n_559), .B1(n_566), .B2(n_576), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_600), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_611), .B(n_568), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_635), .B(n_579), .Y(n_657) );
NOR2x1_ASAP7_75t_L g658 ( .A(n_620), .B(n_566), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_615), .B(n_558), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_602), .A2(n_566), .B1(n_573), .B2(n_560), .C(n_552), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_591), .B(n_560), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_615), .Y(n_662) );
O2A1O1Ixp33_ASAP7_75t_L g663 ( .A1(n_590), .A2(n_73), .B(n_76), .C(n_77), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_594), .B(n_81), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_603), .A2(n_304), .B1(n_289), .B2(n_290), .Y(n_665) );
OAI21xp5_ASAP7_75t_L g666 ( .A1(n_622), .A2(n_624), .B(n_616), .Y(n_666) );
NAND4xp75_ASAP7_75t_L g667 ( .A(n_621), .B(n_287), .C(n_289), .D(n_290), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_625), .B(n_287), .Y(n_668) );
NAND3xp33_ASAP7_75t_SL g669 ( .A(n_619), .B(n_287), .C(n_289), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_618), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_615), .B(n_289), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_613), .A2(n_290), .B(n_627), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_612), .A2(n_290), .B(n_614), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_614), .A2(n_625), .B(n_617), .Y(n_674) );
XOR2x2_ASAP7_75t_L g675 ( .A(n_604), .B(n_597), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_597), .Y(n_676) );
XNOR2xp5_ASAP7_75t_L g677 ( .A(n_598), .B(n_594), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_598), .B(n_633), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_614), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_609), .A2(n_636), .B(n_625), .C(n_621), .Y(n_680) );
INVxp67_ASAP7_75t_L g681 ( .A(n_599), .Y(n_681) );
OA22x2_ASAP7_75t_L g682 ( .A1(n_636), .A2(n_617), .B1(n_629), .B2(n_628), .Y(n_682) );
OAI21xp33_ASAP7_75t_L g683 ( .A1(n_626), .A2(n_609), .B(n_605), .Y(n_683) );
OAI22xp5_ASAP7_75t_SL g684 ( .A1(n_630), .A2(n_633), .B1(n_632), .B2(n_631), .Y(n_684) );
NOR2x1_ASAP7_75t_L g685 ( .A(n_632), .B(n_610), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_606), .Y(n_686) );
INVx2_ASAP7_75t_SL g687 ( .A(n_610), .Y(n_687) );
XNOR2xp5_ASAP7_75t_L g688 ( .A(n_605), .B(n_608), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_601), .A2(n_480), .B1(n_550), .B2(n_477), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_586), .B(n_585), .Y(n_690) );
XNOR2x2_ASAP7_75t_L g691 ( .A(n_607), .B(n_579), .Y(n_691) );
AOI211xp5_ASAP7_75t_L g692 ( .A1(n_657), .A2(n_644), .B(n_666), .C(n_680), .Y(n_692) );
INVxp33_ASAP7_75t_SL g693 ( .A(n_650), .Y(n_693) );
OAI21xp5_ASAP7_75t_L g694 ( .A1(n_643), .A2(n_657), .B(n_637), .Y(n_694) );
XNOR2xp5_ASAP7_75t_L g695 ( .A(n_675), .B(n_689), .Y(n_695) );
OAI21xp5_ASAP7_75t_L g696 ( .A1(n_637), .A2(n_658), .B(n_640), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_648), .B(n_645), .C(n_681), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_674), .A2(n_659), .B(n_662), .C(n_679), .Y(n_698) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_685), .Y(n_699) );
NOR2x1_ASAP7_75t_L g700 ( .A(n_669), .B(n_667), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_690), .Y(n_701) );
OA22x2_ASAP7_75t_L g702 ( .A1(n_677), .A2(n_659), .B1(n_684), .B2(n_642), .Y(n_702) );
OAI22xp5_ASAP7_75t_SL g703 ( .A1(n_659), .A2(n_640), .B1(n_691), .B2(n_651), .Y(n_703) );
OAI211xp5_ASAP7_75t_L g704 ( .A1(n_683), .A2(n_660), .B(n_668), .C(n_664), .Y(n_704) );
AOI21xp33_ASAP7_75t_L g705 ( .A1(n_682), .A2(n_663), .B(n_653), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_676), .B(n_670), .Y(n_706) );
AO22x2_ASAP7_75t_L g707 ( .A1(n_697), .A2(n_639), .B1(n_654), .B2(n_655), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_692), .B(n_652), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_703), .A2(n_690), .B1(n_651), .B2(n_647), .C(n_678), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_701), .B(n_638), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_706), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_694), .A2(n_682), .B1(n_661), .B2(n_665), .C(n_687), .Y(n_712) );
AOI211x1_ASAP7_75t_SL g713 ( .A1(n_696), .A2(n_678), .B(n_668), .C(n_673), .Y(n_713) );
OAI211xp5_ASAP7_75t_L g714 ( .A1(n_705), .A2(n_665), .B(n_671), .C(n_686), .Y(n_714) );
AOI211x1_ASAP7_75t_L g715 ( .A1(n_712), .A2(n_708), .B(n_714), .C(n_702), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_709), .A2(n_702), .B1(n_695), .B2(n_693), .Y(n_716) );
NAND2x1p5_ASAP7_75t_L g717 ( .A(n_711), .B(n_700), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_707), .A2(n_698), .B(n_699), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_710), .Y(n_719) );
NAND5xp2_ASAP7_75t_L g720 ( .A(n_717), .B(n_704), .C(n_707), .D(n_713), .E(n_672), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_719), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_716), .A2(n_649), .B1(n_646), .B2(n_641), .Y(n_722) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_720), .B(n_718), .Y(n_723) );
XNOR2xp5_ASAP7_75t_L g724 ( .A(n_722), .B(n_715), .Y(n_724) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_723), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_725), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_726), .A2(n_724), .B(n_721), .Y(n_727) );
AOI21xp33_ASAP7_75t_SL g728 ( .A1(n_727), .A2(n_688), .B(n_656), .Y(n_728) );
endmodule