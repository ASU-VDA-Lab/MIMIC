module fake_netlist_1_9392_n_681 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_681);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_681;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_74), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_10), .Y(n_87) );
INVx1_ASAP7_75t_SL g88 ( .A(n_13), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_49), .Y(n_89) );
INVx2_ASAP7_75t_SL g90 ( .A(n_60), .Y(n_90) );
BUFx2_ASAP7_75t_L g91 ( .A(n_59), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_76), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_40), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_56), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_38), .Y(n_95) );
OR2x2_ASAP7_75t_L g96 ( .A(n_21), .B(n_5), .Y(n_96) );
HB1xp67_ASAP7_75t_L g97 ( .A(n_9), .Y(n_97) );
BUFx2_ASAP7_75t_L g98 ( .A(n_67), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_22), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_41), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_83), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_48), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_64), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_58), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_4), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_19), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_10), .Y(n_107) );
INVx4_ASAP7_75t_R g108 ( .A(n_0), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_13), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_61), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_14), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_72), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_44), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_68), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_46), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_11), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_57), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_17), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_7), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_7), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_81), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_34), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_93), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_92), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_92), .Y(n_127) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_97), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_87), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_94), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_91), .B(n_1), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_93), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_91), .B(n_3), .Y(n_133) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_94), .A2(n_37), .B(n_84), .Y(n_134) );
BUFx12f_ASAP7_75t_L g135 ( .A(n_98), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_98), .B(n_4), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_95), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_90), .B(n_5), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_90), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_124), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_95), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_105), .B(n_6), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_99), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_99), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_105), .B(n_6), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_86), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_106), .B(n_120), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_100), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_100), .Y(n_149) );
NOR2x1_ASAP7_75t_L g150 ( .A(n_102), .B(n_8), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_102), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_107), .A2(n_8), .B1(n_9), .B2(n_11), .Y(n_152) );
INVx4_ASAP7_75t_L g153 ( .A(n_89), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_110), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_112), .B(n_12), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_153), .B(n_103), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_140), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_153), .B(n_110), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_153), .B(n_113), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_146), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_153), .B(n_104), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_126), .B(n_122), .Y(n_163) );
OAI22xp33_ASAP7_75t_SL g164 ( .A1(n_152), .A2(n_96), .B1(n_121), .B2(n_112), .Y(n_164) );
OAI22xp33_ASAP7_75t_L g165 ( .A1(n_152), .A2(n_114), .B1(n_121), .B2(n_118), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_140), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_129), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_142), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_125), .Y(n_169) );
AOI21x1_ASAP7_75t_L g170 ( .A1(n_126), .A2(n_124), .B(n_123), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_131), .B(n_114), .Y(n_171) );
NOR2x1_ASAP7_75t_L g172 ( .A(n_133), .B(n_136), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_127), .B(n_115), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_140), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_139), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_135), .B(n_119), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_125), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_127), .B(n_123), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_131), .B(n_117), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_131), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_125), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_125), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_135), .B(n_117), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_131), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_142), .B(n_118), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_142), .A2(n_116), .B1(n_109), .B2(n_111), .Y(n_188) );
INVxp67_ASAP7_75t_SL g189 ( .A(n_130), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_135), .B(n_113), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_140), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_147), .B(n_101), .Y(n_192) );
NOR3xp33_ASAP7_75t_L g193 ( .A(n_128), .B(n_155), .C(n_88), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_142), .A2(n_96), .B1(n_108), .B2(n_15), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_189), .B(n_130), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_192), .B(n_137), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_172), .B(n_137), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_172), .B(n_149), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_163), .B(n_149), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_181), .B(n_139), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_181), .B(n_139), .Y(n_201) );
NOR2xp67_ASAP7_75t_L g202 ( .A(n_167), .B(n_144), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_180), .A2(n_145), .B1(n_138), .B2(n_144), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_168), .A2(n_134), .B(n_154), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_181), .B(n_139), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_181), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_185), .B(n_139), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_185), .Y(n_208) );
OR2x2_ASAP7_75t_L g209 ( .A(n_160), .B(n_155), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_173), .B(n_145), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_185), .B(n_154), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_185), .B(n_154), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_168), .A2(n_134), .B(n_148), .Y(n_213) );
NAND2xp33_ASAP7_75t_L g214 ( .A(n_180), .B(n_139), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_171), .B(n_141), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_176), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_171), .B(n_186), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_186), .B(n_141), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_180), .A2(n_150), .B1(n_141), .B2(n_148), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_180), .A2(n_150), .B1(n_143), .B2(n_148), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_186), .B(n_143), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_180), .A2(n_128), .B1(n_143), .B2(n_132), .Y(n_222) );
OAI22xp5_ASAP7_75t_SL g223 ( .A1(n_188), .A2(n_134), .B1(n_132), .B2(n_151), .Y(n_223) );
OR2x2_ASAP7_75t_L g224 ( .A(n_188), .B(n_132), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_186), .B(n_151), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_158), .B(n_151), .Y(n_226) );
INVxp67_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
AND2x6_ASAP7_75t_SL g228 ( .A(n_164), .B(n_12), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_159), .B(n_151), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_168), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_168), .B(n_151), .Y(n_231) );
AND2x4_ASAP7_75t_SL g232 ( .A(n_194), .B(n_151), .Y(n_232) );
AND2x6_ASAP7_75t_SL g233 ( .A(n_164), .B(n_14), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_165), .B(n_15), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_179), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_180), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_180), .B(n_140), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_180), .A2(n_134), .B1(n_17), .B2(n_18), .Y(n_238) );
NOR3xp33_ASAP7_75t_SL g239 ( .A(n_177), .B(n_16), .C(n_18), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_156), .B(n_16), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_193), .A2(n_19), .B1(n_20), .B2(n_23), .Y(n_241) );
AND2x6_ASAP7_75t_SL g242 ( .A(n_184), .B(n_20), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_170), .B(n_24), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_161), .B(n_25), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_176), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_211), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_209), .B(n_176), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_235), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_224), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_234), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_200), .A2(n_201), .B(n_205), .Y(n_251) );
NAND2xp33_ASAP7_75t_L g252 ( .A(n_245), .B(n_191), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_202), .B(n_170), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_200), .A2(n_201), .B(n_205), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_227), .B(n_191), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_207), .A2(n_157), .B(n_162), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_217), .B(n_175), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_224), .A2(n_157), .B(n_162), .C(n_166), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_232), .A2(n_175), .B1(n_166), .B2(n_182), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_210), .B(n_26), .Y(n_260) );
BUFx10_ASAP7_75t_L g261 ( .A(n_242), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_207), .A2(n_187), .B(n_183), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_199), .A2(n_187), .B(n_183), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_196), .B(n_187), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_204), .A2(n_183), .B(n_182), .Y(n_265) );
AO32x2_ASAP7_75t_L g266 ( .A1(n_223), .A2(n_182), .A3(n_178), .B1(n_174), .B2(n_169), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_195), .B(n_178), .Y(n_267) );
INVxp67_ASAP7_75t_L g268 ( .A(n_234), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_213), .A2(n_178), .B(n_174), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g270 ( .A1(n_197), .A2(n_174), .B(n_169), .C(n_29), .Y(n_270) );
CKINVDCx8_ASAP7_75t_R g271 ( .A(n_228), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
NOR2x1_ASAP7_75t_L g273 ( .A(n_240), .B(n_169), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_198), .A2(n_27), .B(n_28), .Y(n_274) );
O2A1O1Ixp5_ASAP7_75t_SL g275 ( .A1(n_231), .A2(n_30), .B(n_31), .C(n_32), .Y(n_275) );
NOR2xp67_ASAP7_75t_L g276 ( .A(n_222), .B(n_33), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_211), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_212), .B(n_35), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_231), .A2(n_36), .B(n_39), .Y(n_279) );
AOI21x1_ASAP7_75t_L g280 ( .A1(n_237), .A2(n_42), .B(n_43), .Y(n_280) );
NOR2xp33_ASAP7_75t_R g281 ( .A(n_214), .B(n_45), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_230), .A2(n_47), .B(n_50), .Y(n_282) );
AO21x1_ASAP7_75t_L g283 ( .A1(n_238), .A2(n_51), .B(n_52), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_203), .B(n_215), .Y(n_284) );
AO21x1_ASAP7_75t_L g285 ( .A1(n_243), .A2(n_53), .B(n_54), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_208), .B(n_55), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_208), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_218), .A2(n_62), .B(n_63), .C(n_65), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_212), .B(n_66), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_221), .A2(n_69), .B(n_70), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_225), .A2(n_71), .B(n_73), .Y(n_291) );
A2O1A1Ixp33_ASAP7_75t_SL g292 ( .A1(n_219), .A2(n_75), .B(n_77), .C(n_78), .Y(n_292) );
XOR2xp5_ASAP7_75t_L g293 ( .A(n_220), .B(n_79), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_208), .B(n_80), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_239), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_267), .Y(n_296) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_253), .A2(n_236), .B(n_214), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_275), .A2(n_244), .B(n_226), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_248), .B(n_206), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g300 ( .A1(n_260), .A2(n_232), .B(n_229), .C(n_241), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_272), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_249), .B(n_233), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_247), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g304 ( .A1(n_268), .A2(n_243), .B(n_216), .C(n_245), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_278), .A2(n_243), .B(n_216), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_264), .Y(n_306) );
OA21x2_ASAP7_75t_L g307 ( .A1(n_285), .A2(n_82), .B(n_85), .Y(n_307) );
AO31x2_ASAP7_75t_L g308 ( .A1(n_283), .A2(n_288), .A3(n_284), .B(n_290), .Y(n_308) );
OAI21x1_ASAP7_75t_L g309 ( .A1(n_280), .A2(n_270), .B(n_265), .Y(n_309) );
AOI221x1_ASAP7_75t_L g310 ( .A1(n_274), .A2(n_282), .B1(n_269), .B2(n_291), .C(n_278), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_272), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_251), .A2(n_254), .B(n_263), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_264), .A2(n_267), .B(n_294), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_294), .A2(n_256), .B(n_262), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_246), .B(n_277), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_272), .B(n_250), .Y(n_316) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_273), .A2(n_279), .B(n_276), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_258), .A2(n_289), .B(n_255), .Y(n_318) );
NAND3x1_ASAP7_75t_L g319 ( .A(n_271), .B(n_261), .C(n_295), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_259), .A2(n_286), .B(n_266), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_257), .A2(n_252), .B(n_287), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_287), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_292), .A2(n_293), .B(n_266), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_261), .A2(n_250), .B1(n_268), .B2(n_249), .Y(n_324) );
INVx5_ASAP7_75t_L g325 ( .A(n_281), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_266), .B(n_248), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_248), .B(n_235), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_264), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_267), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_272), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_268), .A2(n_164), .B(n_165), .C(n_227), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_267), .Y(n_332) );
AO222x2_ASAP7_75t_L g333 ( .A1(n_319), .A2(n_327), .B1(n_331), .B2(n_324), .C1(n_302), .C2(n_299), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_296), .B(n_332), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_313), .A2(n_305), .B(n_312), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_296), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_303), .B(n_332), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_329), .Y(n_338) );
CKINVDCx8_ASAP7_75t_R g339 ( .A(n_325), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_329), .B(n_306), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_306), .B(n_328), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_327), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_314), .A2(n_318), .B(n_300), .Y(n_343) );
AOI21xp33_ASAP7_75t_SL g344 ( .A1(n_316), .A2(n_328), .B(n_307), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_315), .Y(n_345) );
AO21x2_ASAP7_75t_L g346 ( .A1(n_326), .A2(n_323), .B(n_320), .Y(n_346) );
INVx6_ASAP7_75t_L g347 ( .A(n_311), .Y(n_347) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_309), .A2(n_320), .B(n_310), .Y(n_348) );
OAI21xp5_ASAP7_75t_L g349 ( .A1(n_297), .A2(n_321), .B(n_304), .Y(n_349) );
INVx4_ASAP7_75t_SL g350 ( .A(n_311), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_303), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_299), .B(n_322), .Y(n_352) );
OAI21x1_ASAP7_75t_L g353 ( .A1(n_309), .A2(n_298), .B(n_317), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_298), .A2(n_317), .B(n_310), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_299), .B(n_322), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_325), .A2(n_307), .B(n_299), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_330), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_308), .B(n_301), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_330), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_301), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_307), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_338), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_338), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_343), .A2(n_358), .B(n_335), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_348), .Y(n_365) );
AO21x2_ASAP7_75t_L g366 ( .A1(n_344), .A2(n_307), .B(n_308), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_341), .A2(n_325), .B1(n_319), .B2(n_308), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_336), .Y(n_368) );
AO21x2_ASAP7_75t_L g369 ( .A1(n_344), .A2(n_308), .B(n_325), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_336), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_336), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_338), .B(n_308), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_348), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_336), .B(n_325), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_336), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_336), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_348), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_339), .Y(n_378) );
AO31x2_ASAP7_75t_L g379 ( .A1(n_343), .A2(n_325), .A3(n_335), .B(n_358), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_337), .B(n_341), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_348), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_351), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_361), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_334), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_334), .B(n_340), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_361), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_340), .B(n_337), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_361), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_345), .B(n_355), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_342), .B(n_345), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_371), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_362), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_362), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_386), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_372), .B(n_346), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_363), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_386), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_386), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_384), .B(n_342), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_372), .B(n_346), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_386), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_372), .B(n_346), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_384), .B(n_355), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_363), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_383), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_382), .B(n_351), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_382), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_385), .B(n_346), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_383), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_383), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_382), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_371), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_388), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_388), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_385), .B(n_352), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_388), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_365), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_365), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_365), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_385), .B(n_354), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_370), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_371), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_375), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_387), .B(n_390), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_365), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_390), .B(n_352), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_373), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_387), .B(n_354), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_368), .B(n_353), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_418), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_392), .Y(n_431) );
INVxp67_ASAP7_75t_L g432 ( .A(n_407), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_420), .B(n_364), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_420), .B(n_364), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_408), .B(n_380), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_428), .B(n_381), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_424), .B(n_390), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_428), .B(n_381), .Y(n_438) );
NOR2xp67_ASAP7_75t_L g439 ( .A(n_417), .B(n_356), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_395), .B(n_379), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_392), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_393), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_393), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_408), .B(n_381), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_396), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_400), .B(n_381), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_400), .B(n_373), .Y(n_448) );
NOR2x1_ASAP7_75t_L g449 ( .A(n_396), .B(n_378), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_424), .B(n_387), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_404), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_400), .B(n_380), .Y(n_452) );
NOR2x1_ASAP7_75t_L g453 ( .A(n_404), .B(n_378), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_399), .B(n_380), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_417), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_421), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_419), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_419), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_395), .B(n_373), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_399), .B(n_389), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_395), .B(n_373), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_395), .B(n_377), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_415), .B(n_389), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_421), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_418), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_391), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_418), .Y(n_467) );
INVx4_ASAP7_75t_L g468 ( .A(n_412), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_415), .B(n_367), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_402), .B(n_377), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_402), .B(n_377), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_402), .B(n_379), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_425), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_427), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_402), .B(n_379), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_411), .B(n_379), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_394), .B(n_379), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_403), .B(n_367), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_394), .B(n_379), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_411), .B(n_379), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_406), .B(n_379), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_394), .B(n_375), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_397), .B(n_375), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_429), .B(n_369), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_433), .B(n_423), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_452), .B(n_416), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_440), .B(n_429), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_452), .B(n_416), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_456), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_433), .B(n_423), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_434), .B(n_446), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_430), .Y(n_492) );
INVxp67_ASAP7_75t_SL g493 ( .A(n_447), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_434), .B(n_429), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_430), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_435), .B(n_405), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_430), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_450), .B(n_426), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_437), .B(n_426), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_435), .B(n_406), .Y(n_500) );
OAI21xp33_ASAP7_75t_L g501 ( .A1(n_472), .A2(n_475), .B(n_440), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_481), .B(n_409), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_463), .B(n_403), .Y(n_503) );
NAND2x1p5_ASAP7_75t_L g504 ( .A(n_449), .B(n_378), .Y(n_504) );
AND2x2_ASAP7_75t_SL g505 ( .A(n_440), .B(n_397), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_454), .B(n_414), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_481), .B(n_405), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_434), .B(n_429), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_434), .B(n_427), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_444), .B(n_414), .Y(n_510) );
NOR2x1_ASAP7_75t_L g511 ( .A(n_449), .B(n_378), .Y(n_511) );
INVxp67_ASAP7_75t_L g512 ( .A(n_456), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_460), .B(n_413), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_431), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_465), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_465), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_453), .B(n_374), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_431), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_440), .B(n_409), .Y(n_519) );
INVxp67_ASAP7_75t_SL g520 ( .A(n_465), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_446), .B(n_425), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_441), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_467), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_448), .B(n_425), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_467), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_444), .B(n_413), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_441), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_442), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_448), .B(n_401), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_459), .B(n_401), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_436), .B(n_401), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_436), .B(n_438), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_438), .B(n_398), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_442), .B(n_398), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_443), .B(n_398), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_459), .B(n_397), .Y(n_536) );
AOI21xp33_ASAP7_75t_SL g537 ( .A1(n_476), .A2(n_333), .B(n_410), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_467), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_469), .B(n_410), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_461), .B(n_410), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_473), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_484), .B(n_422), .Y(n_542) );
AND2x4_ASAP7_75t_L g543 ( .A(n_484), .B(n_422), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_443), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_473), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_432), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_491), .B(n_472), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_537), .B(n_478), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_514), .Y(n_549) );
OAI221xp5_ASAP7_75t_L g550 ( .A1(n_501), .A2(n_453), .B1(n_480), .B2(n_476), .C(n_464), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_514), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_485), .B(n_477), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_510), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_491), .B(n_475), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_485), .B(n_477), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_518), .Y(n_556) );
AOI21xp33_ASAP7_75t_L g557 ( .A1(n_546), .A2(n_480), .B(n_445), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_518), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_510), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_490), .B(n_479), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_520), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_493), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_505), .A2(n_464), .B1(n_468), .B2(n_474), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_519), .A2(n_461), .B1(n_462), .B2(n_470), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_492), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_489), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_522), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_490), .B(n_462), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_532), .B(n_470), .Y(n_569) );
NAND2x1_ASAP7_75t_L g570 ( .A(n_511), .B(n_468), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_503), .B(n_479), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g572 ( .A(n_500), .B(n_484), .C(n_439), .D(n_445), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_519), .A2(n_484), .B1(n_471), .B2(n_451), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_489), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_519), .A2(n_471), .B1(n_451), .B2(n_455), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_522), .Y(n_576) );
NOR3xp33_ASAP7_75t_L g577 ( .A(n_512), .B(n_357), .C(n_360), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_527), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_509), .B(n_457), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_527), .Y(n_580) );
NOR2xp67_ASAP7_75t_L g581 ( .A(n_487), .B(n_468), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_528), .Y(n_582) );
NOR2xp67_ASAP7_75t_L g583 ( .A(n_487), .B(n_468), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_509), .B(n_455), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_494), .B(n_474), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_539), .B(n_457), .Y(n_586) );
NAND3x1_ASAP7_75t_L g587 ( .A(n_494), .B(n_458), .C(n_466), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_508), .B(n_458), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_539), .B(n_483), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_496), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_498), .B(n_473), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_499), .B(n_483), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_496), .B(n_482), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_528), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_544), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_502), .B(n_482), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_492), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_586), .Y(n_598) );
INVxp67_ASAP7_75t_L g599 ( .A(n_548), .Y(n_599) );
NAND2x1_ASAP7_75t_L g600 ( .A(n_581), .B(n_487), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_583), .A2(n_505), .B(n_502), .C(n_507), .Y(n_601) );
A2O1A1Ixp33_ASAP7_75t_SL g602 ( .A1(n_577), .A2(n_544), .B(n_466), .C(n_349), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_579), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_584), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_561), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_547), .B(n_508), .Y(n_606) );
OAI31xp33_ASAP7_75t_L g607 ( .A1(n_550), .A2(n_504), .A3(n_517), .B(n_543), .Y(n_607) );
INVxp33_ASAP7_75t_L g608 ( .A(n_591), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_561), .B(n_504), .Y(n_609) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_562), .A2(n_513), .B(n_506), .Y(n_610) );
OAI211xp5_ASAP7_75t_SL g611 ( .A1(n_562), .A2(n_486), .B(n_488), .C(n_507), .Y(n_611) );
AOI222xp33_ASAP7_75t_L g612 ( .A1(n_553), .A2(n_526), .B1(n_540), .B2(n_530), .C1(n_536), .C2(n_543), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_565), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_591), .B(n_488), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_554), .B(n_521), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g616 ( .A(n_577), .B(n_439), .C(n_486), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_590), .B(n_521), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_559), .B(n_533), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_568), .B(n_524), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_596), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_587), .A2(n_504), .B1(n_517), .B2(n_531), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_549), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_557), .A2(n_524), .B1(n_529), .B2(n_536), .C(n_530), .Y(n_623) );
OAI21xp33_ASAP7_75t_L g624 ( .A1(n_573), .A2(n_543), .B(n_542), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_573), .A2(n_529), .B1(n_540), .B2(n_542), .C(n_534), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_564), .A2(n_542), .B1(n_535), .B2(n_545), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_563), .B(n_517), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_587), .A2(n_356), .B(n_541), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_572), .A2(n_516), .B1(n_515), .B2(n_497), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_571), .A2(n_516), .B1(n_515), .B2(n_497), .Y(n_630) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_599), .A2(n_566), .B(n_574), .C(n_570), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_607), .B(n_574), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_611), .A2(n_566), .B1(n_592), .B2(n_589), .C(n_575), .Y(n_633) );
XOR2x2_ASAP7_75t_L g634 ( .A(n_600), .B(n_569), .Y(n_634) );
AND3x4_ASAP7_75t_L g635 ( .A(n_627), .B(n_597), .C(n_565), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_602), .A2(n_576), .B(n_595), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_608), .B(n_598), .Y(n_637) );
OAI31xp33_ASAP7_75t_L g638 ( .A1(n_601), .A2(n_588), .A3(n_585), .B(n_552), .Y(n_638) );
OAI22xp33_ASAP7_75t_SL g639 ( .A1(n_627), .A2(n_555), .B1(n_560), .B2(n_593), .Y(n_639) );
AOI322xp5_ASAP7_75t_L g640 ( .A1(n_620), .A2(n_551), .A3(n_594), .B1(n_582), .B2(n_580), .C1(n_578), .C2(n_567), .Y(n_640) );
OA21x2_ASAP7_75t_L g641 ( .A1(n_609), .A2(n_597), .B(n_558), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_625), .A2(n_556), .B1(n_545), .B2(n_495), .C(n_541), .Y(n_642) );
O2A1O1Ixp5_ASAP7_75t_L g643 ( .A1(n_609), .A2(n_538), .B(n_525), .C(n_495), .Y(n_643) );
AOI21xp33_ASAP7_75t_SL g644 ( .A1(n_621), .A2(n_525), .B(n_523), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_610), .A2(n_538), .B1(n_523), .B2(n_349), .C(n_360), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_622), .Y(n_646) );
OAI32xp33_ASAP7_75t_L g647 ( .A1(n_624), .A2(n_466), .A3(n_422), .B1(n_412), .B2(n_376), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_601), .A2(n_466), .B1(n_339), .B2(n_359), .C(n_357), .Y(n_648) );
AOI32xp33_ASAP7_75t_L g649 ( .A1(n_623), .A2(n_374), .A3(n_412), .B1(n_422), .B2(n_368), .Y(n_649) );
AOI222xp33_ASAP7_75t_L g650 ( .A1(n_616), .A2(n_350), .B1(n_374), .B2(n_359), .C1(n_412), .C2(n_354), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_602), .A2(n_374), .B(n_391), .C(n_353), .Y(n_651) );
AOI21xp33_ASAP7_75t_L g652 ( .A1(n_605), .A2(n_369), .B(n_366), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_612), .B(n_369), .Y(n_653) );
NOR3xp33_ASAP7_75t_L g654 ( .A(n_628), .B(n_353), .C(n_368), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_603), .A2(n_369), .B1(n_366), .B2(n_368), .C(n_374), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g656 ( .A1(n_626), .A2(n_391), .B(n_376), .C(n_370), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_629), .A2(n_368), .B1(n_376), .B2(n_370), .Y(n_657) );
OAI21xp5_ASAP7_75t_SL g658 ( .A1(n_629), .A2(n_391), .B(n_371), .Y(n_658) );
XOR2xp5_ASAP7_75t_L g659 ( .A(n_614), .B(n_370), .Y(n_659) );
NAND3xp33_ASAP7_75t_SL g660 ( .A(n_630), .B(n_350), .C(n_347), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_630), .A2(n_347), .B1(n_376), .B2(n_391), .C(n_371), .Y(n_661) );
AOI211x1_ASAP7_75t_SL g662 ( .A1(n_632), .A2(n_636), .B(n_660), .C(n_652), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_637), .B(n_640), .Y(n_663) );
NOR3xp33_ASAP7_75t_L g664 ( .A(n_639), .B(n_631), .C(n_644), .Y(n_664) );
NAND3xp33_ASAP7_75t_SL g665 ( .A(n_635), .B(n_638), .C(n_651), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_634), .A2(n_641), .B(n_643), .Y(n_666) );
AOI311xp33_ASAP7_75t_L g667 ( .A1(n_642), .A2(n_633), .A3(n_654), .B(n_656), .C(n_655), .Y(n_667) );
NAND3x2_ASAP7_75t_L g668 ( .A(n_662), .B(n_653), .C(n_646), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_664), .B(n_606), .Y(n_669) );
NOR3xp33_ASAP7_75t_L g670 ( .A(n_665), .B(n_658), .C(n_647), .Y(n_670) );
NOR4xp25_ASAP7_75t_L g671 ( .A(n_663), .B(n_649), .C(n_648), .D(n_645), .Y(n_671) );
INVxp67_ASAP7_75t_L g672 ( .A(n_669), .Y(n_672) );
AND2x4_ASAP7_75t_L g673 ( .A(n_670), .B(n_604), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_672), .B(n_666), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_673), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_674), .A2(n_668), .B1(n_671), .B2(n_667), .Y(n_676) );
OA21x2_ASAP7_75t_L g677 ( .A1(n_676), .A2(n_675), .B(n_674), .Y(n_677) );
OA22x2_ASAP7_75t_L g678 ( .A1(n_677), .A2(n_659), .B1(n_617), .B2(n_615), .Y(n_678) );
OAI21x1_ASAP7_75t_L g679 ( .A1(n_678), .A2(n_641), .B(n_618), .Y(n_679) );
AO21x2_ASAP7_75t_L g680 ( .A1(n_679), .A2(n_661), .B(n_619), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_680), .A2(n_650), .B1(n_657), .B2(n_613), .Y(n_681) );
endmodule