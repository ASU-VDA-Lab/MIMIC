module fake_jpeg_28053_n_135 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_6),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_29),
.B1(n_27),
.B2(n_30),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_41),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_11),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_24),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_54),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_11),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_50),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_14),
.B(n_12),
.Y(n_49)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_17),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_23),
.C(n_15),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_21),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_16),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_14),
.C(n_12),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_59),
.B(n_68),
.Y(n_83)
);

AND2x4_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_35),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_72),
.B(n_36),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_19),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_16),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_38),
.Y(n_72)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_88),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_36),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_79),
.B(n_81),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_73),
.A2(n_55),
.B1(n_48),
.B2(n_21),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_87),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_16),
.B(n_19),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_61),
.B(n_58),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_36),
.C(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_96),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_64),
.B1(n_62),
.B2(n_58),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_98),
.B1(n_79),
.B2(n_83),
.Y(n_101)
);

AO22x1_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_60),
.B1(n_59),
.B2(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_63),
.C(n_66),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_59),
.C(n_63),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_100),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_105),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_80),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_106),
.C(n_91),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_88),
.B1(n_78),
.B2(n_67),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_60),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_75),
.B1(n_82),
.B2(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_111),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_78),
.B(n_75),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_94),
.C(n_100),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_18),
.C(n_2),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g114 ( 
.A(n_105),
.B(n_87),
.CI(n_60),
.CON(n_114),
.SN(n_114)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_115),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_68),
.B(n_81),
.Y(n_115)
);

OAI321xp33_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_107),
.A3(n_113),
.B1(n_114),
.B2(n_102),
.C(n_112),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_4),
.B(n_5),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_103),
.B1(n_102),
.B2(n_106),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_122),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_113),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_4),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_127),
.A3(n_119),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_120),
.B(n_4),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_5),
.B(n_8),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_129),
.B(n_5),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_130),
.A2(n_131),
.B(n_123),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.C(n_122),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_9),
.Y(n_135)
);


endmodule