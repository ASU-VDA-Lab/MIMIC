module real_aes_873_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_330;
wire n_388;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_484;
wire n_326;
wire n_492;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g218 ( .A(n_0), .B(n_219), .Y(n_218) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_1), .A2(n_55), .B1(n_90), .B2(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g166 ( .A(n_2), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_3), .B(n_224), .Y(n_246) );
NAND2xp33_ASAP7_75t_SL g204 ( .A(n_4), .B(n_205), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_4), .A2(n_81), .B1(n_82), .B2(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_4), .Y(n_493) );
INVx1_ASAP7_75t_L g178 ( .A(n_5), .Y(n_178) );
INVx1_ASAP7_75t_L g147 ( .A(n_6), .Y(n_147) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_7), .A2(n_20), .B1(n_90), .B2(n_91), .Y(n_89) );
AND2x2_ASAP7_75t_L g244 ( .A(n_8), .B(n_227), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_9), .A2(n_44), .B1(n_140), .B2(n_141), .Y(n_139) );
INVx2_ASAP7_75t_L g181 ( .A(n_10), .Y(n_181) );
AOI221x1_ASAP7_75t_L g196 ( .A1(n_11), .A2(n_197), .B1(n_199), .B2(n_200), .C(n_203), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g136 ( .A1(n_12), .A2(n_66), .B1(n_137), .B2(n_138), .Y(n_136) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_13), .A2(n_34), .B1(n_120), .B2(n_123), .Y(n_119) );
INVx1_ASAP7_75t_L g145 ( .A(n_14), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_15), .B(n_224), .Y(n_282) );
INVx1_ASAP7_75t_L g150 ( .A(n_16), .Y(n_150) );
AOI221xp5_ASAP7_75t_SL g291 ( .A1(n_16), .A2(n_32), .B1(n_199), .B2(n_224), .C(n_292), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_17), .A2(n_199), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_18), .B(n_219), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g86 ( .A1(n_19), .A2(n_26), .B1(n_87), .B2(n_103), .Y(n_86) );
OAI221xp5_ASAP7_75t_L g158 ( .A1(n_20), .A2(n_55), .B1(n_57), .B2(n_159), .C(n_161), .Y(n_158) );
OR2x2_ASAP7_75t_L g180 ( .A(n_21), .B(n_68), .Y(n_180) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_21), .A2(n_68), .B(n_181), .Y(n_202) );
INVxp67_ASAP7_75t_L g195 ( .A(n_22), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_23), .B(n_221), .Y(n_286) );
AND2x2_ASAP7_75t_L g238 ( .A(n_24), .B(n_226), .Y(n_238) );
INVx3_ASAP7_75t_L g90 ( .A(n_25), .Y(n_90) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_27), .A2(n_199), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_28), .B(n_221), .Y(n_293) );
INVx1_ASAP7_75t_SL g98 ( .A(n_29), .Y(n_98) );
INVx1_ASAP7_75t_L g168 ( .A(n_30), .Y(n_168) );
AND2x2_ASAP7_75t_L g187 ( .A(n_30), .B(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g205 ( .A(n_30), .B(n_166), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_31), .A2(n_75), .B1(n_132), .B2(n_133), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_33), .A2(n_62), .B1(n_189), .B2(n_199), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_35), .B(n_219), .Y(n_235) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_36), .A2(n_57), .B1(n_90), .B2(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g225 ( .A(n_37), .B(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_38), .B(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_39), .B(n_226), .Y(n_295) );
INVx1_ASAP7_75t_L g185 ( .A(n_40), .Y(n_185) );
INVx1_ASAP7_75t_L g209 ( .A(n_40), .Y(n_209) );
INVx1_ASAP7_75t_L g99 ( .A(n_41), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_42), .B(n_224), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_43), .A2(n_81), .B1(n_82), .B2(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_43), .Y(n_501) );
AND2x2_ASAP7_75t_L g267 ( .A(n_45), .B(n_226), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_46), .B(n_221), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_47), .A2(n_58), .B1(n_128), .B2(n_129), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_48), .B(n_219), .Y(n_265) );
AND2x2_ASAP7_75t_SL g287 ( .A(n_49), .B(n_227), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_50), .A2(n_199), .B(n_233), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g148 ( .A1(n_51), .A2(n_149), .B1(n_150), .B2(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_51), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_52), .B(n_221), .Y(n_250) );
AND2x2_ASAP7_75t_SL g259 ( .A(n_53), .B(n_255), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g112 ( .A1(n_54), .A2(n_59), .B1(n_113), .B2(n_116), .Y(n_112) );
INVxp33_ASAP7_75t_L g163 ( .A(n_55), .Y(n_163) );
INVx1_ASAP7_75t_L g188 ( .A(n_56), .Y(n_188) );
INVx1_ASAP7_75t_L g211 ( .A(n_56), .Y(n_211) );
INVxp67_ASAP7_75t_L g162 ( .A(n_57), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_60), .A2(n_63), .B1(n_182), .B2(n_224), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_61), .B(n_224), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_64), .B(n_219), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_65), .B(n_219), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_67), .A2(n_199), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_69), .B(n_221), .Y(n_264) );
BUFx2_ASAP7_75t_L g80 ( .A(n_70), .Y(n_80) );
INVxp67_ASAP7_75t_L g198 ( .A(n_71), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_72), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_73), .B(n_221), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_74), .A2(n_199), .B(n_284), .Y(n_283) );
BUFx2_ASAP7_75t_SL g160 ( .A(n_76), .Y(n_160) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_155), .B1(n_169), .B2(n_490), .C(n_491), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_143), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_142), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g142 ( .A(n_80), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
NAND2xp5_ASAP7_75t_L g83 ( .A(n_84), .B(n_125), .Y(n_83) );
NOR2xp33_ASAP7_75t_L g84 ( .A(n_85), .B(n_111), .Y(n_84) );
NAND2xp5_ASAP7_75t_SL g85 ( .A(n_86), .B(n_106), .Y(n_85) );
AND2x4_ASAP7_75t_L g87 ( .A(n_88), .B(n_95), .Y(n_87) );
AND2x2_ASAP7_75t_L g120 ( .A(n_88), .B(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g138 ( .A(n_88), .B(n_134), .Y(n_138) );
AND2x4_ASAP7_75t_L g88 ( .A(n_89), .B(n_92), .Y(n_88) );
AND2x2_ASAP7_75t_L g105 ( .A(n_89), .B(n_93), .Y(n_105) );
INVx1_ASAP7_75t_L g110 ( .A(n_89), .Y(n_110) );
INVx1_ASAP7_75t_L g115 ( .A(n_89), .Y(n_115) );
INVx2_ASAP7_75t_L g91 ( .A(n_90), .Y(n_91) );
INVx1_ASAP7_75t_L g94 ( .A(n_90), .Y(n_94) );
OAI22x1_ASAP7_75t_L g96 ( .A1(n_90), .A2(n_97), .B1(n_98), .B2(n_99), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_90), .Y(n_97) );
INVx1_ASAP7_75t_L g102 ( .A(n_90), .Y(n_102) );
AND2x4_ASAP7_75t_L g109 ( .A(n_92), .B(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g124 ( .A(n_92), .Y(n_124) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
AND2x2_ASAP7_75t_L g114 ( .A(n_93), .B(n_115), .Y(n_114) );
AND2x4_ASAP7_75t_L g113 ( .A(n_95), .B(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g132 ( .A(n_95), .B(n_109), .Y(n_132) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_100), .Y(n_95) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_96), .Y(n_104) );
AND2x2_ASAP7_75t_L g108 ( .A(n_96), .B(n_101), .Y(n_108) );
INVx2_ASAP7_75t_L g122 ( .A(n_96), .Y(n_122) );
AND2x4_ASAP7_75t_L g134 ( .A(n_100), .B(n_122), .Y(n_134) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g121 ( .A(n_101), .B(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g130 ( .A(n_101), .Y(n_130) );
AND2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x4_ASAP7_75t_L g129 ( .A(n_105), .B(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g133 ( .A(n_105), .B(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x2_ASAP7_75t_L g116 ( .A(n_108), .B(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g123 ( .A(n_108), .B(n_124), .Y(n_123) );
AND2x6_ASAP7_75t_L g137 ( .A(n_109), .B(n_121), .Y(n_137) );
AND2x2_ASAP7_75t_L g140 ( .A(n_109), .B(n_134), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_119), .Y(n_111) );
AND2x2_ASAP7_75t_L g128 ( .A(n_114), .B(n_121), .Y(n_128) );
AND2x6_ASAP7_75t_L g141 ( .A(n_114), .B(n_134), .Y(n_141) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_115), .Y(n_118) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_135), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_131), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_139), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B1(n_146), .B2(n_154), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_146), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B1(n_152), .B2(n_153), .Y(n_146) );
INVx1_ASAP7_75t_L g152 ( .A(n_147), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_148), .Y(n_153) );
INVx1_ASAP7_75t_L g151 ( .A(n_150), .Y(n_151) );
INVx1_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_157), .Y(n_156) );
AND3x1_ASAP7_75t_SL g157 ( .A(n_158), .B(n_164), .C(n_167), .Y(n_157) );
INVxp67_ASAP7_75t_L g499 ( .A(n_158), .Y(n_499) );
CKINVDCx8_ASAP7_75t_R g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_164), .Y(n_497) );
AO21x1_ASAP7_75t_SL g505 ( .A1(n_164), .A2(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g183 ( .A(n_165), .B(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_SL g504 ( .A(n_165), .B(n_167), .Y(n_504) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g193 ( .A(n_166), .B(n_185), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_167), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2x1p5_ASAP7_75t_L g190 ( .A(n_168), .B(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_171), .B(n_367), .Y(n_170) );
NOR4xp25_ASAP7_75t_L g171 ( .A(n_172), .B(n_310), .C(n_349), .D(n_356), .Y(n_171) );
OAI221xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_228), .B1(n_268), .B2(n_277), .C(n_296), .Y(n_172) );
OR2x2_ASAP7_75t_L g440 ( .A(n_173), .B(n_302), .Y(n_440) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g355 ( .A(n_174), .B(n_280), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_174), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_174), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g174 ( .A(n_175), .B(n_212), .Y(n_174) );
AND2x4_ASAP7_75t_SL g279 ( .A(n_175), .B(n_280), .Y(n_279) );
INVx3_ASAP7_75t_L g301 ( .A(n_175), .Y(n_301) );
AND2x2_ASAP7_75t_L g336 ( .A(n_175), .B(n_309), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_175), .B(n_213), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_175), .B(n_303), .Y(n_388) );
OR2x2_ASAP7_75t_L g466 ( .A(n_175), .B(n_280), .Y(n_466) );
AND2x4_ASAP7_75t_L g175 ( .A(n_176), .B(n_196), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_182), .B1(n_189), .B2(n_194), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_179), .B(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_179), .B(n_198), .Y(n_197) );
NOR3xp33_ASAP7_75t_L g203 ( .A(n_179), .B(n_204), .C(n_206), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_179), .A2(n_246), .B(n_247), .Y(n_245) );
AND2x4_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
AND2x2_ASAP7_75t_SL g227 ( .A(n_180), .B(n_181), .Y(n_227) );
AND2x4_ASAP7_75t_L g182 ( .A(n_183), .B(n_186), .Y(n_182) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_184), .Y(n_507) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x4_ASAP7_75t_L g221 ( .A(n_185), .B(n_210), .Y(n_221) );
BUFx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x6_ASAP7_75t_L g199 ( .A(n_187), .B(n_193), .Y(n_199) );
INVx2_ASAP7_75t_L g192 ( .A(n_188), .Y(n_192) );
AND2x6_ASAP7_75t_L g219 ( .A(n_188), .B(n_208), .Y(n_219) );
AND2x4_ASAP7_75t_L g189 ( .A(n_190), .B(n_193), .Y(n_189) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_190), .Y(n_506) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx4_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AOI21x1_ASAP7_75t_L g214 ( .A1(n_201), .A2(n_215), .B(n_225), .Y(n_214) );
INVx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx4f_ASAP7_75t_L g255 ( .A(n_202), .Y(n_255) );
INVx5_ASAP7_75t_L g222 ( .A(n_205), .Y(n_222) );
AND2x4_ASAP7_75t_L g224 ( .A(n_205), .B(n_207), .Y(n_224) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_210), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g288 ( .A(n_213), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_213), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g314 ( .A(n_213), .Y(n_314) );
OR2x2_ASAP7_75t_L g319 ( .A(n_213), .B(n_303), .Y(n_319) );
AND2x2_ASAP7_75t_L g332 ( .A(n_213), .B(n_290), .Y(n_332) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_213), .Y(n_335) );
INVx1_ASAP7_75t_L g347 ( .A(n_213), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_213), .B(n_301), .Y(n_412) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_223), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_220), .B(n_222), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_222), .A2(n_234), .B(n_235), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_222), .A2(n_249), .B(n_250), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_222), .A2(n_264), .B(n_265), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_222), .A2(n_285), .B(n_286), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_222), .A2(n_293), .B(n_294), .Y(n_292) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_224), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_226), .Y(n_237) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_226), .A2(n_291), .B(n_295), .Y(n_290) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_229), .B(n_239), .Y(n_228) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g276 ( .A(n_230), .B(n_260), .Y(n_276) );
AND2x4_ASAP7_75t_L g306 ( .A(n_230), .B(n_243), .Y(n_306) );
INVx2_ASAP7_75t_L g340 ( .A(n_230), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_230), .B(n_260), .Y(n_398) );
AND2x2_ASAP7_75t_L g445 ( .A(n_230), .B(n_274), .Y(n_445) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_237), .B(n_238), .Y(n_230) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_231), .A2(n_237), .B(n_238), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_236), .Y(n_231) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_237), .A2(n_261), .B(n_267), .Y(n_260) );
AOI222xp33_ASAP7_75t_L g433 ( .A1(n_239), .A2(n_305), .B1(n_348), .B2(n_408), .C1(n_434), .C2(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_251), .Y(n_240) );
AND2x2_ASAP7_75t_L g352 ( .A(n_241), .B(n_272), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_241), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g481 ( .A(n_241), .B(n_321), .Y(n_481) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_242), .A2(n_312), .B(n_316), .Y(n_311) );
AND2x2_ASAP7_75t_L g392 ( .A(n_242), .B(n_275), .Y(n_392) );
OR2x2_ASAP7_75t_L g417 ( .A(n_242), .B(n_276), .Y(n_417) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx5_ASAP7_75t_L g271 ( .A(n_243), .Y(n_271) );
AND2x2_ASAP7_75t_L g358 ( .A(n_243), .B(n_340), .Y(n_358) );
AND2x2_ASAP7_75t_L g384 ( .A(n_243), .B(n_260), .Y(n_384) );
OR2x2_ASAP7_75t_L g387 ( .A(n_243), .B(n_274), .Y(n_387) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_243), .Y(n_405) );
AND2x4_ASAP7_75t_SL g462 ( .A(n_243), .B(n_339), .Y(n_462) );
OR2x2_ASAP7_75t_L g471 ( .A(n_243), .B(n_298), .Y(n_471) );
OR2x6_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g304 ( .A(n_251), .Y(n_304) );
AOI221xp5_ASAP7_75t_SL g422 ( .A1(n_251), .A2(n_306), .B1(n_423), .B2(n_425), .C(n_426), .Y(n_422) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_260), .Y(n_251) );
OR2x2_ASAP7_75t_L g361 ( .A(n_252), .B(n_331), .Y(n_361) );
OR2x2_ASAP7_75t_L g371 ( .A(n_252), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g397 ( .A(n_252), .B(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g403 ( .A(n_252), .B(n_322), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_252), .B(n_386), .Y(n_415) );
INVx2_ASAP7_75t_L g428 ( .A(n_252), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_252), .B(n_306), .Y(n_449) );
AND2x2_ASAP7_75t_L g453 ( .A(n_252), .B(n_275), .Y(n_453) );
AND2x2_ASAP7_75t_L g461 ( .A(n_252), .B(n_462), .Y(n_461) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g274 ( .A(n_253), .Y(n_274) );
AOI21x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_256), .B(n_259), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_255), .A2(n_282), .B(n_283), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_260), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g305 ( .A(n_260), .B(n_274), .Y(n_305) );
INVx2_ASAP7_75t_L g322 ( .A(n_260), .Y(n_322) );
AND2x4_ASAP7_75t_L g339 ( .A(n_260), .B(n_340), .Y(n_339) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_260), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_266), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g451 ( .A(n_270), .B(n_273), .Y(n_451) );
AND2x4_ASAP7_75t_L g297 ( .A(n_271), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g338 ( .A(n_271), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g365 ( .A(n_271), .B(n_305), .Y(n_365) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
AND2x2_ASAP7_75t_L g469 ( .A(n_273), .B(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g321 ( .A(n_274), .B(n_322), .Y(n_321) );
OAI21xp5_ASAP7_75t_SL g341 ( .A1(n_275), .A2(n_342), .B(n_348), .Y(n_341) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_288), .Y(n_278) );
INVx1_ASAP7_75t_SL g395 ( .A(n_279), .Y(n_395) );
AND2x2_ASAP7_75t_L g425 ( .A(n_279), .B(n_335), .Y(n_425) );
AND2x4_ASAP7_75t_L g436 ( .A(n_279), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g302 ( .A(n_280), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g309 ( .A(n_280), .Y(n_309) );
AND2x4_ASAP7_75t_L g315 ( .A(n_280), .B(n_301), .Y(n_315) );
INVx2_ASAP7_75t_L g326 ( .A(n_280), .Y(n_326) );
INVx1_ASAP7_75t_L g375 ( .A(n_280), .Y(n_375) );
OR2x2_ASAP7_75t_L g396 ( .A(n_280), .B(n_380), .Y(n_396) );
OR2x2_ASAP7_75t_L g410 ( .A(n_280), .B(n_290), .Y(n_410) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_280), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_280), .B(n_332), .Y(n_482) );
OR2x6_ASAP7_75t_L g280 ( .A(n_281), .B(n_287), .Y(n_280) );
INVx1_ASAP7_75t_L g327 ( .A(n_288), .Y(n_327) );
AND2x2_ASAP7_75t_L g460 ( .A(n_288), .B(n_326), .Y(n_460) );
AND2x2_ASAP7_75t_L g485 ( .A(n_288), .B(n_315), .Y(n_485) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g303 ( .A(n_290), .Y(n_303) );
BUFx3_ASAP7_75t_L g345 ( .A(n_290), .Y(n_345) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_290), .Y(n_372) );
INVx1_ASAP7_75t_L g381 ( .A(n_290), .Y(n_381) );
AOI33xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_299), .A3(n_304), .B1(n_305), .B2(n_306), .B3(n_307), .Y(n_296) );
AOI21x1_ASAP7_75t_SL g399 ( .A1(n_297), .A2(n_321), .B(n_383), .Y(n_399) );
INVx2_ASAP7_75t_L g429 ( .A(n_297), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_297), .B(n_428), .Y(n_435) );
AND2x2_ASAP7_75t_L g383 ( .A(n_298), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g346 ( .A(n_301), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g447 ( .A(n_302), .Y(n_447) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_303), .Y(n_437) );
OAI32xp33_ASAP7_75t_L g486 ( .A1(n_304), .A2(n_306), .A3(n_482), .B1(n_487), .B2(n_489), .Y(n_486) );
AND2x2_ASAP7_75t_L g404 ( .A(n_305), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_SL g394 ( .A(n_306), .Y(n_394) );
AND2x2_ASAP7_75t_L g459 ( .A(n_306), .B(n_403), .Y(n_459) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI221xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_320), .B1(n_323), .B2(n_337), .C(n_341), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_314), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_315), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_315), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_315), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g364 ( .A(n_319), .Y(n_364) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR3xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_328), .C(n_333), .Y(n_323) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_325), .A2(n_387), .B1(n_427), .B2(n_430), .Y(n_426) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g330 ( .A(n_326), .Y(n_330) );
NOR2x1p5_ASAP7_75t_L g344 ( .A(n_326), .B(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_326), .Y(n_366) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI322xp33_ASAP7_75t_L g393 ( .A1(n_329), .A2(n_371), .A3(n_394), .B1(n_395), .B2(n_396), .C1(n_397), .C2(n_399), .Y(n_393) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_331), .A2(n_350), .B(n_351), .C(n_353), .Y(n_349) );
OR2x2_ASAP7_75t_L g441 ( .A(n_331), .B(n_395), .Y(n_441) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g348 ( .A(n_332), .B(n_336), .Y(n_348) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g354 ( .A(n_338), .B(n_355), .Y(n_354) );
INVx3_ASAP7_75t_SL g386 ( .A(n_339), .Y(n_386) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_343), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx1_ASAP7_75t_SL g390 ( .A(n_346), .Y(n_390) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_347), .Y(n_432) );
OR2x6_ASAP7_75t_SL g487 ( .A(n_350), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI211xp5_ASAP7_75t_L g477 ( .A1(n_355), .A2(n_478), .B(n_479), .C(n_486), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_359), .B(n_362), .C(n_366), .Y(n_356) );
OAI211xp5_ASAP7_75t_SL g368 ( .A1(n_357), .A2(n_369), .B(n_376), .C(n_400), .Y(n_368) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
NOR3xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_413), .C(n_457), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_373), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_372), .Y(n_464) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g419 ( .A(n_375), .Y(n_419) );
NOR3xp33_ASAP7_75t_SL g376 ( .A(n_377), .B(n_389), .C(n_393), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_382), .B1(n_385), .B2(n_388), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_381), .Y(n_488) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_SL g474 ( .A(n_387), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
OR2x2_ASAP7_75t_L g424 ( .A(n_390), .B(n_410), .Y(n_424) );
OR2x2_ASAP7_75t_L g475 ( .A(n_390), .B(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g473 ( .A(n_398), .Y(n_473) );
OR2x2_ASAP7_75t_L g489 ( .A(n_398), .B(n_428), .Y(n_489) );
OAI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_404), .B(n_406), .Y(n_400) );
OAI31xp33_ASAP7_75t_L g414 ( .A1(n_401), .A2(n_415), .A3(n_416), .B(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g446 ( .A(n_411), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND4xp25_ASAP7_75t_SL g413 ( .A(n_414), .B(n_422), .C(n_433), .D(n_438), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_421), .Y(n_456) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_442), .B1(n_446), .B2(n_448), .C(n_450), .Y(n_438) );
NAND2xp33_ASAP7_75t_SL g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx1_ASAP7_75t_L g483 ( .A(n_442), .Y(n_483) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_443), .B(n_445), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g478 ( .A(n_452), .Y(n_478) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_458), .B(n_477), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B1(n_461), .B2(n_463), .C(n_467), .Y(n_458) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
AOI21xp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_472), .B(n_475), .Y(n_467) );
INVxp33_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_482), .B1(n_483), .B2(n_484), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI222xp33_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B1(n_494), .B2(n_500), .C1(n_502), .C2(n_505), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_496), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
endmodule