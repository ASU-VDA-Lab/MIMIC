module fake_netlist_5_1650_n_1538 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_145, n_48, n_50, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_149, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1538);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_145;
input n_48;
input n_50;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_149;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1538;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_851;
wire n_615;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_980;
wire n_1115;
wire n_703;
wire n_698;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_175),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_159),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_191),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_106),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_56),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_7),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_298),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_235),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_230),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_324),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_61),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_243),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_132),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_118),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_234),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_239),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_219),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_196),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_141),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_102),
.Y(n_352)
);

BUFx2_ASAP7_75t_SL g353 ( 
.A(n_170),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_244),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_197),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_139),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_135),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_256),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_314),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_17),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_86),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_49),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_182),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_125),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_156),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_100),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_258),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_94),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_123),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_238),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_91),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_282),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_310),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_249),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_8),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_283),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_267),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_207),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_322),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_23),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_262),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_287),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_233),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_299),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_325),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_292),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_180),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_248),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_176),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_127),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_38),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_1),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_321),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_252),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_47),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_172),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_82),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_60),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_229),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_206),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_202),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_6),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_327),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_275),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_221),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_6),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_315),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_291),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_320),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_96),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_178),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_177),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_136),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_190),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_254),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_130),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_203),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_104),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_308),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_154),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_316),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_165),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_59),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_121),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_13),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_146),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_245),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_122),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_107),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_331),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_309),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_164),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_212),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_220),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_240),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_140),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_38),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_60),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_251),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_195),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_192),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_20),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_247),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_163),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_193),
.Y(n_445)
);

BUFx8_ASAP7_75t_SL g446 ( 
.A(n_297),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_168),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_73),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_128),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_40),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_306),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_242),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_278),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_72),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_37),
.Y(n_455)
);

BUFx10_ASAP7_75t_L g456 ( 
.A(n_25),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_46),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_41),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_208),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_32),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_31),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_44),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_2),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_200),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_185),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_41),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_83),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_63),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_27),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_276),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_289),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_183),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_305),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_15),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_120),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_270),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_255),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_259),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_326),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_300),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_79),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_209),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_26),
.Y(n_483)
);

BUFx2_ASAP7_75t_SL g484 ( 
.A(n_137),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_225),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_319),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_103),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_149),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_266),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_199),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_8),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_105),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_186),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_85),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_201),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_174),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_69),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_133),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_13),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_285),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_210),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_188),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_171),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_157),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_37),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_11),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_92),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_26),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_119),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_279),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_296),
.Y(n_511)
);

BUFx5_ASAP7_75t_L g512 ( 
.A(n_131),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_250),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_76),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_293),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_317),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_67),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_169),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_21),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_216),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_65),
.Y(n_521)
);

BUFx10_ASAP7_75t_L g522 ( 
.A(n_155),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_145),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_81),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_161),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_227),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_218),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_134),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_151),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_113),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_260),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_284),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_328),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_74),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_318),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_280),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_273),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_74),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_101),
.Y(n_539)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_286),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_48),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_263),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_246),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_126),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_45),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_265),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_281),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_49),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_269),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_116),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_187),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_40),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_179),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_14),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_15),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_152),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_112),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_129),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_261),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_78),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_68),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_194),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_142),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_514),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_372),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_372),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_372),
.Y(n_567)
);

AND2x6_ASAP7_75t_L g568 ( 
.A(n_372),
.B(n_84),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_514),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_402),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_514),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_349),
.B(n_0),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_370),
.B(n_0),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_400),
.B(n_87),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_370),
.B(n_1),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_420),
.B(n_2),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_421),
.B(n_3),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_436),
.B(n_3),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_400),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_373),
.B(n_4),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_451),
.B(n_4),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_514),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_373),
.B(n_5),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_451),
.B(n_5),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_402),
.B(n_7),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_336),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_511),
.B(n_9),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_400),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_551),
.B(n_9),
.Y(n_589)
);

CKINVDCx16_ASAP7_75t_R g590 ( 
.A(n_388),
.Y(n_590)
);

BUFx8_ASAP7_75t_SL g591 ( 
.A(n_446),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_496),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_553),
.B(n_10),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_435),
.B(n_10),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_332),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_464),
.B(n_11),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_531),
.B(n_12),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_384),
.Y(n_598)
);

BUFx8_ASAP7_75t_SL g599 ( 
.A(n_446),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_384),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_513),
.B(n_374),
.Y(n_601)
);

INVx5_ASAP7_75t_L g602 ( 
.A(n_537),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_337),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_384),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_537),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_540),
.B(n_12),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_374),
.B(n_14),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_474),
.B(n_16),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_456),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_474),
.B(n_16),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_537),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_537),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_387),
.B(n_17),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_561),
.Y(n_614)
);

INVx5_ASAP7_75t_L g615 ( 
.A(n_546),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_563),
.B(n_18),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_387),
.B(n_18),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_389),
.B(n_19),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_389),
.B(n_19),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_561),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_561),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_403),
.B(n_20),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_546),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_546),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_546),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_456),
.Y(n_626)
);

NOR2x1_ASAP7_75t_L g627 ( 
.A(n_506),
.B(n_88),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_403),
.B(n_21),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_522),
.Y(n_629)
);

INVx5_ASAP7_75t_L g630 ( 
.A(n_561),
.Y(n_630)
);

BUFx8_ASAP7_75t_SL g631 ( 
.A(n_460),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_417),
.B(n_22),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_506),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_517),
.B(n_360),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_417),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_517),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_538),
.Y(n_637)
);

BUFx8_ASAP7_75t_SL g638 ( 
.A(n_460),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_522),
.B(n_22),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_343),
.Y(n_640)
);

BUFx8_ASAP7_75t_SL g641 ( 
.A(n_481),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_456),
.B(n_23),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_441),
.B(n_24),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_522),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_563),
.B(n_24),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_441),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_333),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_375),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_444),
.B(n_89),
.Y(n_649)
);

NOR2x1_ASAP7_75t_L g650 ( 
.A(n_542),
.B(n_27),
.Y(n_650)
);

INVx5_ASAP7_75t_L g651 ( 
.A(n_512),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_512),
.B(n_28),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_512),
.B(n_29),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_338),
.B(n_29),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_512),
.B(n_30),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_340),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_380),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_334),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_391),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_335),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_512),
.B(n_30),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_341),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_362),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_512),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_346),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_369),
.B(n_31),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_512),
.B(n_32),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_353),
.Y(n_668)
);

INVx5_ASAP7_75t_L g669 ( 
.A(n_484),
.Y(n_669)
);

INVx5_ASAP7_75t_L g670 ( 
.A(n_398),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_355),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_357),
.B(n_33),
.Y(n_672)
);

BUFx8_ASAP7_75t_SL g673 ( 
.A(n_481),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_483),
.B(n_33),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_361),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_392),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_395),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_406),
.B(n_34),
.Y(n_678)
);

BUFx12f_ASAP7_75t_L g679 ( 
.A(n_425),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_454),
.Y(n_680)
);

BUFx12f_ASAP7_75t_L g681 ( 
.A(n_437),
.Y(n_681)
);

INVx5_ASAP7_75t_L g682 ( 
.A(n_442),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_448),
.B(n_34),
.Y(n_683)
);

INVx5_ASAP7_75t_L g684 ( 
.A(n_450),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_463),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_455),
.B(n_35),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_376),
.B(n_35),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_378),
.Y(n_688)
);

INVx5_ASAP7_75t_L g689 ( 
.A(n_457),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_469),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_385),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_386),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_458),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_401),
.Y(n_694)
);

INVx5_ASAP7_75t_L g695 ( 
.A(n_461),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_497),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_462),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_409),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_412),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_475),
.B(n_36),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_413),
.B(n_416),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_424),
.B(n_36),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_429),
.B(n_39),
.Y(n_703)
);

BUFx12f_ASAP7_75t_L g704 ( 
.A(n_466),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_430),
.B(n_39),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_432),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_521),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_339),
.Y(n_708)
);

INVx5_ASAP7_75t_L g709 ( 
.A(n_468),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_548),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_465),
.Y(n_711)
);

AND2x6_ASAP7_75t_L g712 ( 
.A(n_467),
.B(n_90),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_473),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_479),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_486),
.Y(n_715)
);

BUFx12f_ASAP7_75t_L g716 ( 
.A(n_491),
.Y(n_716)
);

AND2x6_ASAP7_75t_L g717 ( 
.A(n_490),
.B(n_93),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_586),
.B(n_344),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_603),
.B(n_345),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_648),
.B(n_347),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_564),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_657),
.B(n_348),
.Y(n_722)
);

BUFx10_ASAP7_75t_L g723 ( 
.A(n_601),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_659),
.B(n_350),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_581),
.A2(n_414),
.B1(n_516),
.B2(n_342),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_569),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_629),
.B(n_501),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_620),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_620),
.Y(n_729)
);

OAI22xp33_ASAP7_75t_L g730 ( 
.A1(n_606),
.A2(n_505),
.B1(n_508),
.B2(n_499),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_596),
.A2(n_545),
.B1(n_438),
.B2(n_423),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_566),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_647),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_566),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_SL g735 ( 
.A(n_584),
.B(n_342),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_SL g736 ( 
.A1(n_629),
.A2(n_545),
.B1(n_555),
.B2(n_414),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_566),
.Y(n_737)
);

AO22x2_ASAP7_75t_L g738 ( 
.A1(n_573),
.A2(n_515),
.B1(n_523),
.B2(n_504),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_571),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_567),
.Y(n_740)
);

AO22x2_ASAP7_75t_L g741 ( 
.A1(n_573),
.A2(n_575),
.B1(n_583),
.B2(n_580),
.Y(n_741)
);

AO22x2_ASAP7_75t_L g742 ( 
.A1(n_575),
.A2(n_532),
.B1(n_557),
.B2(n_526),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_SL g743 ( 
.A1(n_590),
.A2(n_516),
.B1(n_547),
.B2(n_525),
.Y(n_743)
);

AO22x2_ASAP7_75t_L g744 ( 
.A1(n_580),
.A2(n_559),
.B1(n_44),
.B2(n_42),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_594),
.A2(n_519),
.B1(n_534),
.B2(n_524),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_597),
.A2(n_552),
.B1(n_554),
.B2(n_541),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_590),
.A2(n_525),
.B1(n_556),
.B2(n_547),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_644),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_592),
.A2(n_556),
.B1(n_354),
.B2(n_560),
.Y(n_749)
);

OAI22xp33_ASAP7_75t_L g750 ( 
.A1(n_592),
.A2(n_352),
.B1(n_356),
.B2(n_351),
.Y(n_750)
);

OAI22xp33_ASAP7_75t_SL g751 ( 
.A1(n_639),
.A2(n_359),
.B1(n_363),
.B2(n_358),
.Y(n_751)
);

AO22x2_ASAP7_75t_L g752 ( 
.A1(n_583),
.A2(n_45),
.B1(n_42),
.B2(n_43),
.Y(n_752)
);

OAI22xp33_ASAP7_75t_R g753 ( 
.A1(n_609),
.A2(n_47),
.B1(n_43),
.B2(n_46),
.Y(n_753)
);

BUFx6f_ASAP7_75t_SL g754 ( 
.A(n_598),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_595),
.B(n_658),
.Y(n_755)
);

OAI22xp33_ASAP7_75t_L g756 ( 
.A1(n_626),
.A2(n_365),
.B1(n_366),
.B2(n_364),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_640),
.B(n_367),
.Y(n_757)
);

INVx4_ASAP7_75t_L g758 ( 
.A(n_708),
.Y(n_758)
);

OAI22xp33_ASAP7_75t_SL g759 ( 
.A1(n_572),
.A2(n_371),
.B1(n_377),
.B2(n_368),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_571),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_666),
.A2(n_381),
.B1(n_382),
.B2(n_379),
.Y(n_761)
);

AO22x2_ASAP7_75t_L g762 ( 
.A1(n_642),
.A2(n_51),
.B1(n_48),
.B2(n_50),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_600),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_700),
.A2(n_390),
.B1(n_393),
.B2(n_383),
.Y(n_764)
);

AOI22x1_ASAP7_75t_L g765 ( 
.A1(n_616),
.A2(n_396),
.B1(n_397),
.B2(n_394),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_697),
.B(n_399),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_679),
.A2(n_405),
.B1(n_407),
.B2(n_404),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_681),
.A2(n_410),
.B1(n_411),
.B2(n_408),
.Y(n_768)
);

AO22x2_ASAP7_75t_L g769 ( 
.A1(n_616),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_634),
.B(n_415),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_567),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_604),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_704),
.A2(n_485),
.B1(n_558),
.B2(n_550),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_582),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_582),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_SL g776 ( 
.A1(n_576),
.A2(n_562),
.B1(n_549),
.B2(n_544),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_570),
.B(n_52),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_L g778 ( 
.A1(n_644),
.A2(n_543),
.B1(n_539),
.B2(n_536),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_567),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_716),
.A2(n_535),
.B1(n_533),
.B2(n_530),
.Y(n_780)
);

INVx5_ASAP7_75t_L g781 ( 
.A(n_579),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_631),
.Y(n_782)
);

OR2x6_ASAP7_75t_L g783 ( 
.A(n_633),
.B(n_53),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_644),
.B(n_418),
.Y(n_784)
);

OA22x2_ASAP7_75t_L g785 ( 
.A1(n_707),
.A2(n_529),
.B1(n_528),
.B2(n_527),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_SL g786 ( 
.A1(n_702),
.A2(n_520),
.B1(n_518),
.B2(n_510),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_660),
.B(n_419),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_579),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_633),
.B(n_422),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_674),
.A2(n_472),
.B1(n_507),
.B2(n_503),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_678),
.A2(n_686),
.B1(n_683),
.B2(n_617),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_614),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_636),
.B(n_426),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_636),
.B(n_670),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_670),
.B(n_682),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_579),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_614),
.Y(n_797)
);

NAND2x1p5_ASAP7_75t_L g798 ( 
.A(n_670),
.B(n_427),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_621),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_621),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_613),
.A2(n_509),
.B1(n_502),
.B2(n_500),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_577),
.B(n_428),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_623),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_623),
.Y(n_804)
);

OAI22xp33_ASAP7_75t_SL g805 ( 
.A1(n_578),
.A2(n_498),
.B1(n_495),
.B2(n_494),
.Y(n_805)
);

BUFx6f_ASAP7_75t_SL g806 ( 
.A(n_591),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_682),
.B(n_431),
.Y(n_807)
);

OAI22xp33_ASAP7_75t_L g808 ( 
.A1(n_587),
.A2(n_493),
.B1(n_492),
.B2(n_489),
.Y(n_808)
);

OA22x2_ASAP7_75t_L g809 ( 
.A1(n_710),
.A2(n_488),
.B1(n_487),
.B2(n_482),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_682),
.B(n_433),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_623),
.Y(n_811)
);

AND2x2_ASAP7_75t_SL g812 ( 
.A(n_632),
.B(n_53),
.Y(n_812)
);

OR2x6_ASAP7_75t_L g813 ( 
.A(n_676),
.B(n_54),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_618),
.A2(n_480),
.B1(n_478),
.B2(n_477),
.Y(n_814)
);

NOR2x1p5_ASAP7_75t_L g815 ( 
.A(n_607),
.B(n_434),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_624),
.Y(n_816)
);

OAI22xp33_ASAP7_75t_L g817 ( 
.A1(n_589),
.A2(n_476),
.B1(n_471),
.B2(n_470),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_684),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_624),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_624),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_723),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_803),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_735),
.B(n_684),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_757),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_755),
.B(n_684),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_723),
.B(n_689),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_741),
.A2(n_701),
.B(n_628),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_747),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_803),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_791),
.B(n_668),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_741),
.A2(n_793),
.B(n_789),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_730),
.B(n_668),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_820),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_820),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_770),
.B(n_689),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_788),
.Y(n_836)
);

XNOR2xp5_ASAP7_75t_L g837 ( 
.A(n_743),
.B(n_599),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_788),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_732),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_734),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_781),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_739),
.B(n_664),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_737),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_740),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_771),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_779),
.Y(n_846)
);

AND2x6_ASAP7_75t_L g847 ( 
.A(n_727),
.B(n_632),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_796),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_758),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_802),
.B(n_689),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_804),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_811),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_816),
.Y(n_853)
);

XNOR2x2_ASAP7_75t_L g854 ( 
.A(n_769),
.B(n_650),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_819),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_766),
.B(n_693),
.Y(n_856)
);

XNOR2x2_ASAP7_75t_L g857 ( 
.A(n_769),
.B(n_650),
.Y(n_857)
);

AND2x2_ASAP7_75t_SL g858 ( 
.A(n_812),
.B(n_643),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_728),
.Y(n_859)
);

INVxp33_ASAP7_75t_L g860 ( 
.A(n_736),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_729),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_758),
.B(n_693),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_750),
.B(n_693),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_721),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_726),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_739),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_794),
.A2(n_645),
.B(n_619),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_733),
.Y(n_868)
);

XOR2x2_ASAP7_75t_L g869 ( 
.A(n_731),
.B(n_638),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_760),
.B(n_635),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_760),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_774),
.Y(n_872)
);

XNOR2xp5_ASAP7_75t_L g873 ( 
.A(n_725),
.B(n_731),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_756),
.B(n_761),
.Y(n_874)
);

INVxp67_ASAP7_75t_SL g875 ( 
.A(n_774),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_815),
.B(n_585),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_749),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_775),
.Y(n_878)
);

INVx4_ASAP7_75t_SL g879 ( 
.A(n_783),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_775),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_792),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_792),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_797),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_785),
.A2(n_809),
.B(n_765),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_797),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_718),
.B(n_695),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_801),
.B(n_668),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_719),
.B(n_720),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_799),
.Y(n_889)
);

XOR2xp5_ASAP7_75t_L g890 ( 
.A(n_782),
.B(n_439),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_799),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_800),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_722),
.B(n_695),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_800),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_777),
.B(n_763),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_764),
.B(n_695),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_781),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_781),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_783),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_787),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_772),
.Y(n_901)
);

AND2x2_ASAP7_75t_SL g902 ( 
.A(n_724),
.B(n_643),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_738),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_814),
.B(n_709),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_738),
.Y(n_905)
);

XOR2xp5_ASAP7_75t_L g906 ( 
.A(n_767),
.B(n_440),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_742),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_742),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_807),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_810),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_813),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_813),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_784),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_875),
.B(n_815),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_902),
.B(n_744),
.Y(n_915)
);

AND2x2_ASAP7_75t_SL g916 ( 
.A(n_858),
.B(n_654),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_888),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_875),
.B(n_765),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_870),
.Y(n_919)
);

AND2x6_ASAP7_75t_L g920 ( 
.A(n_903),
.B(n_627),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_866),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_909),
.B(n_654),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_871),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_872),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_895),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_878),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_870),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_910),
.B(n_744),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_880),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_868),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_867),
.B(n_790),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_852),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_913),
.B(n_752),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_867),
.B(n_808),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_831),
.B(n_817),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_821),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_830),
.B(n_752),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_847),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_852),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_821),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_881),
.Y(n_941)
);

OAI21x1_ASAP7_75t_L g942 ( 
.A1(n_827),
.A2(n_653),
.B(n_652),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_908),
.B(n_745),
.Y(n_943)
);

INVx4_ASAP7_75t_L g944 ( 
.A(n_847),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_882),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_852),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_847),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_843),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_905),
.B(n_907),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_830),
.B(n_762),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_864),
.Y(n_951)
);

NAND2x1p5_ASAP7_75t_L g952 ( 
.A(n_824),
.B(n_795),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_827),
.B(n_669),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_R g954 ( 
.A(n_849),
.B(n_806),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_883),
.Y(n_955)
);

AND2x2_ASAP7_75t_SL g956 ( 
.A(n_874),
.B(n_655),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_865),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_847),
.B(n_669),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_900),
.B(n_762),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_885),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_876),
.B(n_884),
.Y(n_961)
);

INVxp67_ASAP7_75t_SL g962 ( 
.A(n_842),
.Y(n_962)
);

NAND2x1p5_ASAP7_75t_L g963 ( 
.A(n_823),
.B(n_818),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_841),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_889),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_884),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_891),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_892),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_894),
.Y(n_969)
);

INVxp67_ASAP7_75t_SL g970 ( 
.A(n_842),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_R g971 ( 
.A(n_877),
.B(n_806),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_854),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_839),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_822),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_876),
.B(n_712),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_856),
.B(n_712),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_886),
.B(n_608),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_893),
.B(n_610),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_840),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_832),
.B(n_714),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_829),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_833),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_832),
.A2(n_717),
.B(n_712),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_857),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_850),
.B(n_669),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_859),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_834),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_826),
.B(n_663),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_835),
.B(n_663),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_844),
.B(n_712),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_825),
.B(n_887),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_887),
.B(n_717),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_896),
.B(n_685),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_861),
.B(n_685),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_845),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_904),
.B(n_690),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_846),
.Y(n_997)
);

AND2x2_ASAP7_75t_SL g998 ( 
.A(n_863),
.B(n_661),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_848),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_879),
.B(n_751),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_851),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_853),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_841),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_855),
.B(n_717),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_901),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_899),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_911),
.B(n_786),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_879),
.B(n_676),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_879),
.B(n_677),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_921),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_939),
.Y(n_1011)
);

NAND2x1_ASAP7_75t_SL g1012 ( 
.A(n_915),
.B(n_912),
.Y(n_1012)
);

OR2x6_ASAP7_75t_L g1013 ( 
.A(n_930),
.B(n_862),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_924),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_949),
.B(n_1008),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_924),
.Y(n_1016)
);

INVxp67_ASAP7_75t_SL g1017 ( 
.A(n_939),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_1008),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_949),
.B(n_836),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_917),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_939),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_966),
.B(n_746),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_949),
.B(n_838),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_945),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_962),
.B(n_759),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_921),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_1008),
.B(n_768),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_945),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_925),
.Y(n_1029)
);

AND2x6_ASAP7_75t_L g1030 ( 
.A(n_947),
.B(n_667),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_939),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_1009),
.B(n_961),
.Y(n_1032)
);

NAND2x1p5_ASAP7_75t_L g1033 ( 
.A(n_947),
.B(n_748),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_923),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_980),
.B(n_873),
.Y(n_1035)
);

OR2x6_ASAP7_75t_L g1036 ( 
.A(n_930),
.B(n_677),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_970),
.B(n_776),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_980),
.B(n_860),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_961),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_936),
.B(n_940),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_988),
.B(n_906),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_1006),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_1005),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_919),
.B(n_805),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_939),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_927),
.B(n_635),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_991),
.B(n_828),
.Y(n_1047)
);

INVx5_ASAP7_75t_L g1048 ( 
.A(n_975),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_1009),
.B(n_773),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_914),
.B(n_641),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_915),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_1009),
.B(n_780),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_968),
.B(n_680),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_943),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_975),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_975),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_965),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_923),
.B(n_680),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_956),
.B(n_635),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_926),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_956),
.B(n_646),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_1005),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_943),
.B(n_890),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_994),
.Y(n_1064)
);

NAND2x1p5_ASAP7_75t_L g1065 ( 
.A(n_938),
.B(n_897),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_981),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_955),
.B(n_646),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_988),
.B(n_869),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_SL g1069 ( 
.A(n_916),
.B(n_568),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_965),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_974),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_926),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_955),
.B(n_646),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_916),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_972),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_972),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_981),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_938),
.B(n_898),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_955),
.B(n_778),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_981),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_974),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_929),
.B(n_696),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_984),
.B(n_837),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_977),
.B(n_709),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_984),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_994),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_929),
.B(n_696),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_969),
.B(n_649),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_977),
.B(n_690),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_969),
.B(n_649),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_941),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1039),
.B(n_998),
.Y(n_1092)
);

BUFx12f_ASAP7_75t_L g1093 ( 
.A(n_1036),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1014),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1016),
.Y(n_1095)
);

INVx5_ASAP7_75t_L g1096 ( 
.A(n_1055),
.Y(n_1096)
);

INVx5_ASAP7_75t_SL g1097 ( 
.A(n_1055),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_1040),
.Y(n_1098)
);

INVx3_ASAP7_75t_SL g1099 ( 
.A(n_1029),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1024),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_1043),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_1036),
.Y(n_1102)
);

BUFx2_ASAP7_75t_R g1103 ( 
.A(n_1083),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1028),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_1029),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1057),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1038),
.B(n_998),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1055),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_1056),
.Y(n_1109)
);

INVx6_ASAP7_75t_L g1110 ( 
.A(n_1048),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_1018),
.Y(n_1111)
);

BUFx12f_ASAP7_75t_L g1112 ( 
.A(n_1036),
.Y(n_1112)
);

INVx5_ASAP7_75t_L g1113 ( 
.A(n_1056),
.Y(n_1113)
);

BUFx2_ASAP7_75t_SL g1114 ( 
.A(n_1048),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1035),
.B(n_1007),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_1054),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_1042),
.Y(n_1117)
);

BUFx12f_ASAP7_75t_L g1118 ( 
.A(n_1013),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1010),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_1056),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1011),
.Y(n_1121)
);

INVx4_ASAP7_75t_L g1122 ( 
.A(n_1066),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1066),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1026),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_1051),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_1064),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1066),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1032),
.B(n_941),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1077),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_1032),
.B(n_960),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_1075),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1086),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_1015),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_1015),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1070),
.B(n_978),
.Y(n_1135)
);

BUFx8_ASAP7_75t_L g1136 ( 
.A(n_1076),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1034),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1060),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_1085),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1071),
.B(n_978),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_1077),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1077),
.Y(n_1142)
);

BUFx12f_ASAP7_75t_L g1143 ( 
.A(n_1013),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_1012),
.Y(n_1144)
);

BUFx2_ASAP7_75t_SL g1145 ( 
.A(n_1048),
.Y(n_1145)
);

NAND2xp33_ASAP7_75t_L g1146 ( 
.A(n_1080),
.B(n_947),
.Y(n_1146)
);

INVx3_ASAP7_75t_SL g1147 ( 
.A(n_1013),
.Y(n_1147)
);

BUFx2_ASAP7_75t_SL g1148 ( 
.A(n_1080),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1020),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_1041),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1072),
.Y(n_1151)
);

INVx5_ASAP7_75t_L g1152 ( 
.A(n_1080),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1011),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_1011),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_1031),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_SL g1156 ( 
.A(n_1047),
.B(n_673),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1081),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1063),
.B(n_950),
.Y(n_1158)
);

BUFx10_ASAP7_75t_L g1159 ( 
.A(n_1050),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1019),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1019),
.Y(n_1161)
);

BUFx12f_ASAP7_75t_L g1162 ( 
.A(n_1027),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1022),
.B(n_993),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1163),
.A2(n_1061),
.B(n_1059),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1094),
.Y(n_1165)
);

CKINVDCx11_ASAP7_75t_R g1166 ( 
.A(n_1099),
.Y(n_1166)
);

CKINVDCx6p67_ASAP7_75t_R g1167 ( 
.A(n_1099),
.Y(n_1167)
);

BUFx4f_ASAP7_75t_SL g1168 ( 
.A(n_1099),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1107),
.A2(n_950),
.B1(n_937),
.B2(n_931),
.Y(n_1169)
);

BUFx8_ASAP7_75t_L g1170 ( 
.A(n_1093),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1149),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1101),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1157),
.Y(n_1173)
);

BUFx12f_ASAP7_75t_L g1174 ( 
.A(n_1093),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1107),
.B(n_1022),
.Y(n_1175)
);

INVx6_ASAP7_75t_L g1176 ( 
.A(n_1136),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1157),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1094),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1115),
.B(n_1068),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1095),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1095),
.Y(n_1181)
);

INVx6_ASAP7_75t_L g1182 ( 
.A(n_1136),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1100),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_1150),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1100),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_1150),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1119),
.Y(n_1187)
);

BUFx12f_ASAP7_75t_L g1188 ( 
.A(n_1102),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1092),
.A2(n_937),
.B1(n_934),
.B2(n_1058),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1119),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1135),
.B(n_1089),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_SL g1192 ( 
.A1(n_1156),
.A2(n_1102),
.B1(n_1112),
.B2(n_1158),
.Y(n_1192)
);

OAI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1140),
.A2(n_1069),
.B1(n_1074),
.B2(n_1044),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_1116),
.Y(n_1194)
);

BUFx2_ASAP7_75t_SL g1195 ( 
.A(n_1101),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1104),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1106),
.A2(n_1037),
.B1(n_1025),
.B2(n_1062),
.Y(n_1197)
);

OAI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1106),
.A2(n_1069),
.B1(n_1044),
.B2(n_1025),
.Y(n_1198)
);

BUFx12f_ASAP7_75t_L g1199 ( 
.A(n_1112),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1124),
.Y(n_1200)
);

CKINVDCx11_ASAP7_75t_R g1201 ( 
.A(n_1147),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1149),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_SL g1203 ( 
.A1(n_1162),
.A2(n_971),
.B1(n_954),
.B2(n_754),
.Y(n_1203)
);

OAI21xp33_ASAP7_75t_L g1204 ( 
.A1(n_1105),
.A2(n_1037),
.B(n_959),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1124),
.Y(n_1205)
);

OAI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1131),
.A2(n_1079),
.B1(n_1091),
.B2(n_935),
.Y(n_1206)
);

CKINVDCx6p67_ASAP7_75t_R g1207 ( 
.A(n_1111),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_SL g1208 ( 
.A1(n_1162),
.A2(n_754),
.B1(n_1052),
.B2(n_1049),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1125),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1137),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1137),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1128),
.A2(n_1079),
.B1(n_992),
.B2(n_1017),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1110),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1128),
.A2(n_1058),
.B1(n_1087),
.B2(n_1082),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1138),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1128),
.A2(n_1082),
.B1(n_1087),
.B2(n_753),
.Y(n_1216)
);

OAI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1147),
.A2(n_1061),
.B1(n_1059),
.B2(n_918),
.Y(n_1217)
);

BUFx4f_ASAP7_75t_SL g1218 ( 
.A(n_1118),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_1139),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1116),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1130),
.A2(n_753),
.B1(n_622),
.B2(n_920),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1130),
.A2(n_920),
.B1(n_1053),
.B2(n_967),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1159),
.A2(n_920),
.B1(n_983),
.B2(n_993),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1151),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1151),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1096),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1121),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_SL g1228 ( 
.A1(n_1144),
.A2(n_1000),
.B(n_959),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1130),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1108),
.Y(n_1230)
);

OAI22xp33_ASAP7_75t_SL g1231 ( 
.A1(n_1139),
.A2(n_1000),
.B1(n_593),
.B2(n_1046),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1144),
.A2(n_944),
.B1(n_938),
.B2(n_969),
.Y(n_1232)
);

OR2x2_ASAP7_75t_SL g1233 ( 
.A(n_1176),
.B(n_1103),
.Y(n_1233)
);

AOI222xp33_ASAP7_75t_L g1234 ( 
.A1(n_1221),
.A2(n_1216),
.B1(n_1175),
.B2(n_1169),
.C1(n_1189),
.C2(n_1191),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1227),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1165),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1171),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_SL g1238 ( 
.A1(n_1168),
.A2(n_1159),
.B1(n_1143),
.B2(n_1125),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1221),
.A2(n_1143),
.B1(n_1147),
.B2(n_687),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1219),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1179),
.B(n_1098),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1204),
.A2(n_703),
.B1(n_705),
.B2(n_672),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_SL g1243 ( 
.A1(n_1208),
.A2(n_963),
.B(n_952),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1169),
.B(n_1098),
.Y(n_1244)
);

OAI21xp33_ASAP7_75t_L g1245 ( 
.A1(n_1189),
.A2(n_996),
.B(n_989),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1178),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1185),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1197),
.A2(n_920),
.B1(n_1053),
.B2(n_1084),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1192),
.A2(n_920),
.B1(n_1134),
.B2(n_1133),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1206),
.A2(n_1134),
.B1(n_1133),
.B2(n_967),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1206),
.A2(n_960),
.B1(n_928),
.B2(n_933),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1168),
.A2(n_963),
.B1(n_1132),
.B2(n_1126),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1214),
.A2(n_1117),
.B1(n_1132),
.B2(n_1126),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1227),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1193),
.A2(n_982),
.B1(n_987),
.B2(n_922),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1228),
.B(n_1160),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1196),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1214),
.A2(n_1160),
.B1(n_1161),
.B2(n_952),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1231),
.B(n_1161),
.Y(n_1259)
);

BUFx4f_ASAP7_75t_SL g1260 ( 
.A(n_1194),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1198),
.A2(n_922),
.B1(n_1002),
.B2(n_1046),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1198),
.A2(n_1002),
.B1(n_951),
.B2(n_957),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1164),
.A2(n_986),
.B1(n_999),
.B2(n_995),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1202),
.B(n_989),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1223),
.A2(n_1001),
.B1(n_942),
.B2(n_1030),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1229),
.B(n_1108),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1166),
.A2(n_1030),
.B1(n_981),
.B2(n_1111),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1176),
.A2(n_947),
.B1(n_1030),
.B2(n_944),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1180),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1184),
.B(n_1023),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1176),
.A2(n_947),
.B1(n_1030),
.B2(n_944),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1180),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1222),
.A2(n_1097),
.B1(n_1110),
.B2(n_1109),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1166),
.A2(n_981),
.B1(n_979),
.B2(n_973),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1181),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_SL g1276 ( 
.A1(n_1203),
.A2(n_976),
.B(n_958),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1209),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1181),
.Y(n_1278)
);

BUFx12f_ASAP7_75t_L g1279 ( 
.A(n_1201),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1201),
.A2(n_942),
.B1(n_656),
.B2(n_665),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1172),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1173),
.A2(n_656),
.B1(n_665),
.B2(n_662),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1186),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1167),
.A2(n_1097),
.B1(n_1110),
.B2(n_1109),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_SL g1285 ( 
.A1(n_1217),
.A2(n_976),
.B(n_798),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_1220),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1177),
.A2(n_656),
.B1(n_665),
.B2(n_662),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1183),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1183),
.B(n_1108),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_SL g1290 ( 
.A1(n_1182),
.A2(n_1145),
.B1(n_1114),
.B2(n_1146),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1195),
.A2(n_1097),
.B1(n_1120),
.B2(n_1113),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1172),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1213),
.B(n_1023),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1182),
.A2(n_1114),
.B1(n_1145),
.B2(n_1146),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1239),
.A2(n_1218),
.B1(n_1182),
.B2(n_1207),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1234),
.A2(n_1188),
.B1(n_1199),
.B2(n_1174),
.Y(n_1296)
);

OAI222xp33_ASAP7_75t_L g1297 ( 
.A1(n_1239),
.A2(n_1212),
.B1(n_1200),
.B2(n_1225),
.C1(n_1218),
.C2(n_1187),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1242),
.B(n_953),
.C(n_985),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1252),
.A2(n_1213),
.B1(n_1232),
.B2(n_1120),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1245),
.A2(n_1170),
.B1(n_649),
.B2(n_574),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1241),
.B(n_1240),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1243),
.A2(n_1226),
.B1(n_1230),
.B2(n_1211),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1256),
.A2(n_1170),
.B1(n_1226),
.B2(n_1148),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1244),
.A2(n_649),
.B1(n_574),
.B2(n_568),
.Y(n_1304)
);

INVxp67_ASAP7_75t_SL g1305 ( 
.A(n_1237),
.Y(n_1305)
);

NAND3xp33_ASAP7_75t_L g1306 ( 
.A(n_1242),
.B(n_671),
.C(n_662),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1259),
.A2(n_574),
.B1(n_568),
.B2(n_973),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1258),
.A2(n_1148),
.B1(n_976),
.B2(n_1113),
.Y(n_1308)
);

AOI21xp33_ASAP7_75t_L g1309 ( 
.A1(n_1248),
.A2(n_1210),
.B(n_1205),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1264),
.A2(n_574),
.B1(n_568),
.B2(n_973),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1281),
.Y(n_1311)
);

NAND3xp33_ASAP7_75t_L g1312 ( 
.A(n_1263),
.B(n_445),
.C(n_443),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1279),
.A2(n_997),
.B1(n_979),
.B2(n_1190),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1255),
.A2(n_997),
.B1(n_979),
.B2(n_1215),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1255),
.B(n_1210),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1249),
.A2(n_948),
.B1(n_1224),
.B2(n_932),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1251),
.A2(n_1096),
.B1(n_1113),
.B2(n_1078),
.Y(n_1317)
);

OAI221xp5_ASAP7_75t_L g1318 ( 
.A1(n_1285),
.A2(n_1276),
.B1(n_1238),
.B2(n_1267),
.C(n_1250),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1270),
.A2(n_1004),
.B1(n_990),
.B2(n_452),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1233),
.A2(n_1096),
.B1(n_1113),
.B2(n_1078),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1261),
.A2(n_1073),
.B(n_1067),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1253),
.A2(n_447),
.B1(n_449),
.B2(n_459),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1260),
.A2(n_1113),
.B1(n_1096),
.B2(n_1227),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1269),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1277),
.A2(n_990),
.B1(n_1004),
.B2(n_453),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1272),
.B(n_1227),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1278),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1273),
.A2(n_1096),
.B1(n_1113),
.B2(n_1152),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1293),
.A2(n_1261),
.B1(n_1263),
.B2(n_1262),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1288),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1262),
.A2(n_1123),
.B1(n_1127),
.B2(n_1129),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1275),
.B(n_1123),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1280),
.A2(n_1073),
.B(n_1067),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1274),
.A2(n_1096),
.B1(n_1065),
.B2(n_1152),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1236),
.B(n_1129),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1265),
.A2(n_1142),
.B1(n_699),
.B2(n_691),
.Y(n_1336)
);

OAI222xp33_ASAP7_75t_L g1337 ( 
.A1(n_1290),
.A2(n_1141),
.B1(n_1122),
.B2(n_637),
.C1(n_1090),
.C2(n_1088),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1283),
.A2(n_706),
.B1(n_713),
.B2(n_671),
.Y(n_1338)
);

OAI222xp33_ASAP7_75t_L g1339 ( 
.A1(n_1294),
.A2(n_1141),
.B1(n_1122),
.B2(n_1090),
.C1(n_1088),
.C2(n_1154),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1286),
.A2(n_699),
.B1(n_711),
.B2(n_671),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1280),
.A2(n_706),
.B1(n_713),
.B2(n_675),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1246),
.A2(n_1257),
.B(n_1247),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1292),
.A2(n_698),
.B1(n_715),
.B2(n_675),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1266),
.B(n_1121),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1268),
.A2(n_711),
.B1(n_715),
.B2(n_688),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1271),
.A2(n_1065),
.B1(n_1152),
.B2(n_1033),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1284),
.A2(n_698),
.B1(n_713),
.B2(n_688),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1291),
.A2(n_1152),
.B1(n_1122),
.B2(n_1153),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1289),
.B(n_1121),
.Y(n_1349)
);

NOR3xp33_ASAP7_75t_L g1350 ( 
.A(n_1282),
.B(n_1154),
.C(n_946),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1282),
.A2(n_692),
.B1(n_711),
.B2(n_691),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1287),
.A2(n_692),
.B1(n_694),
.B2(n_715),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1287),
.A2(n_694),
.B1(n_1045),
.B2(n_1021),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1301),
.B(n_1235),
.Y(n_1354)
);

AOI21xp33_ASAP7_75t_L g1355 ( 
.A1(n_1322),
.A2(n_1296),
.B(n_1312),
.Y(n_1355)
);

AOI221xp5_ASAP7_75t_L g1356 ( 
.A1(n_1306),
.A2(n_1318),
.B1(n_1297),
.B2(n_1302),
.C(n_1340),
.Y(n_1356)
);

NOR3xp33_ASAP7_75t_SL g1357 ( 
.A(n_1295),
.B(n_54),
.C(n_55),
.Y(n_1357)
);

OAI21xp33_ASAP7_75t_L g1358 ( 
.A1(n_1322),
.A2(n_1254),
.B(n_1235),
.Y(n_1358)
);

NOR3xp33_ASAP7_75t_SL g1359 ( 
.A(n_1320),
.B(n_1254),
.C(n_1235),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1303),
.A2(n_1254),
.B(n_55),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_SL g1361 ( 
.A(n_1299),
.B(n_1154),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1305),
.B(n_56),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1329),
.A2(n_1155),
.B1(n_1153),
.B2(n_1121),
.Y(n_1363)
);

NOR3xp33_ASAP7_75t_L g1364 ( 
.A(n_1298),
.B(n_1045),
.C(n_1021),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1311),
.B(n_57),
.Y(n_1365)
);

OAI221xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1338),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.C(n_61),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1311),
.B(n_625),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1327),
.B(n_58),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1330),
.B(n_62),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1326),
.B(n_64),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1319),
.A2(n_64),
.B(n_65),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1324),
.B(n_66),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1308),
.A2(n_1155),
.B1(n_1153),
.B2(n_1121),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1324),
.B(n_66),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1335),
.B(n_67),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1317),
.A2(n_651),
.B1(n_1155),
.B2(n_1153),
.Y(n_1376)
);

AOI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1349),
.A2(n_1344),
.B(n_1315),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_SL g1378 ( 
.A1(n_1325),
.A2(n_69),
.B(n_70),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1332),
.B(n_70),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1332),
.B(n_71),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1342),
.B(n_1315),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1350),
.A2(n_1155),
.B1(n_1153),
.B2(n_1031),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1313),
.A2(n_1155),
.B1(n_1031),
.B2(n_565),
.Y(n_1383)
);

OAI21xp33_ASAP7_75t_L g1384 ( 
.A1(n_1336),
.A2(n_1341),
.B(n_1343),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1307),
.A2(n_1323),
.B(n_1348),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1342),
.B(n_71),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1342),
.B(n_72),
.Y(n_1387)
);

OAI21xp33_ASAP7_75t_L g1388 ( 
.A1(n_1347),
.A2(n_625),
.B(n_75),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1328),
.B(n_73),
.Y(n_1389)
);

AOI21xp33_ASAP7_75t_L g1390 ( 
.A1(n_1298),
.A2(n_75),
.B(n_76),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1309),
.B(n_77),
.Y(n_1391)
);

NAND3xp33_ASAP7_75t_L g1392 ( 
.A(n_1300),
.B(n_630),
.C(n_588),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1334),
.B(n_588),
.Y(n_1393)
);

AO22x1_ASAP7_75t_L g1394 ( 
.A1(n_1346),
.A2(n_1321),
.B1(n_1333),
.B2(n_1337),
.Y(n_1394)
);

NAND3xp33_ASAP7_75t_L g1395 ( 
.A(n_1316),
.B(n_630),
.C(n_588),
.Y(n_1395)
);

AOI221xp5_ASAP7_75t_L g1396 ( 
.A1(n_1339),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.C(n_615),
.Y(n_1396)
);

OAI221xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1345),
.A2(n_80),
.B1(n_95),
.B2(n_97),
.C(n_98),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1354),
.B(n_1331),
.Y(n_1398)
);

OAI211xp5_ASAP7_75t_L g1399 ( 
.A1(n_1357),
.A2(n_1304),
.B(n_1352),
.C(n_1351),
.Y(n_1399)
);

OAI211xp5_ASAP7_75t_L g1400 ( 
.A1(n_1357),
.A2(n_1353),
.B(n_1310),
.C(n_1314),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_L g1401 ( 
.A(n_1371),
.B(n_99),
.C(n_108),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1370),
.B(n_109),
.Y(n_1402)
);

NOR3xp33_ASAP7_75t_L g1403 ( 
.A(n_1378),
.B(n_110),
.C(n_111),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1386),
.B(n_114),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1387),
.B(n_115),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1381),
.B(n_117),
.Y(n_1406)
);

INVx5_ASAP7_75t_L g1407 ( 
.A(n_1372),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1377),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1365),
.B(n_124),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1367),
.Y(n_1410)
);

NOR3xp33_ASAP7_75t_L g1411 ( 
.A(n_1355),
.B(n_138),
.C(n_143),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1362),
.B(n_1375),
.Y(n_1412)
);

BUFx12f_ASAP7_75t_L g1413 ( 
.A(n_1389),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1368),
.B(n_144),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1390),
.A2(n_612),
.B(n_611),
.Y(n_1415)
);

NAND3xp33_ASAP7_75t_L g1416 ( 
.A(n_1356),
.B(n_612),
.C(n_611),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1374),
.Y(n_1417)
);

INVx3_ASAP7_75t_SL g1418 ( 
.A(n_1393),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1369),
.B(n_1379),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1380),
.B(n_147),
.Y(n_1420)
);

INVxp67_ASAP7_75t_SL g1421 ( 
.A(n_1364),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1391),
.Y(n_1422)
);

NAND4xp75_ASAP7_75t_L g1423 ( 
.A(n_1396),
.B(n_148),
.C(n_150),
.D(n_153),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1359),
.B(n_158),
.Y(n_1424)
);

AOI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1366),
.A2(n_605),
.B1(n_602),
.B2(n_166),
.C(n_167),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1394),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1358),
.B(n_1363),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1407),
.B(n_1376),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1407),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1408),
.B(n_1364),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1407),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1407),
.B(n_1412),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_SL g1433 ( 
.A1(n_1426),
.A2(n_1376),
.B1(n_1382),
.B2(n_1373),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1410),
.B(n_1385),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1417),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1422),
.B(n_1361),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1419),
.B(n_1360),
.Y(n_1437)
);

XOR2x2_ASAP7_75t_L g1438 ( 
.A(n_1403),
.B(n_1366),
.Y(n_1438)
);

NAND4xp25_ASAP7_75t_L g1439 ( 
.A(n_1425),
.B(n_1397),
.C(n_1388),
.D(n_1384),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1406),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1421),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1427),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1398),
.Y(n_1443)
);

OAI31xp33_ASAP7_75t_L g1444 ( 
.A1(n_1403),
.A2(n_1392),
.A3(n_1395),
.B(n_1383),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1405),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1404),
.Y(n_1446)
);

NAND4xp75_ASAP7_75t_L g1447 ( 
.A(n_1425),
.B(n_160),
.C(n_162),
.D(n_173),
.Y(n_1447)
);

XOR2x2_ASAP7_75t_L g1448 ( 
.A(n_1401),
.B(n_181),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1435),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1432),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1441),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1443),
.B(n_1418),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1429),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1430),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1429),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1438),
.A2(n_1401),
.B1(n_1416),
.B2(n_1423),
.Y(n_1456)
);

XNOR2x1_ASAP7_75t_L g1457 ( 
.A(n_1448),
.B(n_1420),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1430),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1440),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1432),
.B(n_1440),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1431),
.B(n_1404),
.Y(n_1461)
);

XOR2x2_ASAP7_75t_L g1462 ( 
.A(n_1437),
.B(n_1447),
.Y(n_1462)
);

XNOR2x1_ASAP7_75t_L g1463 ( 
.A(n_1437),
.B(n_1414),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1431),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_R g1465 ( 
.A(n_1436),
.B(n_1413),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1434),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1428),
.B(n_1424),
.Y(n_1467)
);

AO22x2_ASAP7_75t_L g1468 ( 
.A1(n_1436),
.A2(n_1411),
.B1(n_1424),
.B2(n_1415),
.Y(n_1468)
);

INVx1_ASAP7_75t_SL g1469 ( 
.A(n_1434),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1456),
.A2(n_1439),
.B1(n_1433),
.B2(n_1442),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1458),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1458),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1452),
.Y(n_1473)
);

AO22x2_ASAP7_75t_L g1474 ( 
.A1(n_1453),
.A2(n_1428),
.B1(n_1445),
.B2(n_1446),
.Y(n_1474)
);

AOI22x1_ASAP7_75t_L g1475 ( 
.A1(n_1468),
.A2(n_1446),
.B1(n_1409),
.B2(n_1402),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1449),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1454),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1459),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1451),
.Y(n_1479)
);

OA22x2_ASAP7_75t_L g1480 ( 
.A1(n_1467),
.A2(n_1400),
.B1(n_1399),
.B2(n_1444),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1460),
.Y(n_1481)
);

AO22x2_ASAP7_75t_L g1482 ( 
.A1(n_1453),
.A2(n_1399),
.B1(n_189),
.B2(n_198),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1471),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1479),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1478),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1472),
.Y(n_1486)
);

OAI322xp33_ASAP7_75t_L g1487 ( 
.A1(n_1480),
.A2(n_1463),
.A3(n_1457),
.B1(n_1469),
.B2(n_1466),
.C1(n_1450),
.C2(n_1455),
.Y(n_1487)
);

XOR2x2_ASAP7_75t_L g1488 ( 
.A(n_1470),
.B(n_1462),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1481),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1473),
.B(n_1463),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1476),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1477),
.Y(n_1492)
);

AOI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1487),
.A2(n_1482),
.B1(n_1474),
.B2(n_1455),
.C(n_1467),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_SL g1494 ( 
.A1(n_1490),
.A2(n_1457),
.B1(n_1465),
.B2(n_1475),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1484),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1489),
.A2(n_1461),
.B1(n_1464),
.B2(n_605),
.Y(n_1496)
);

AND4x1_ASAP7_75t_L g1497 ( 
.A(n_1488),
.B(n_1461),
.C(n_204),
.D(n_205),
.Y(n_1497)
);

OAI322xp33_ASAP7_75t_L g1498 ( 
.A1(n_1483),
.A2(n_184),
.A3(n_211),
.B1(n_213),
.B2(n_214),
.C1(n_215),
.C2(n_217),
.Y(n_1498)
);

AOI221xp5_ASAP7_75t_L g1499 ( 
.A1(n_1493),
.A2(n_1485),
.B1(n_1486),
.B2(n_1492),
.C(n_1491),
.Y(n_1499)
);

OAI22x1_ASAP7_75t_L g1500 ( 
.A1(n_1497),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1495),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1496),
.Y(n_1502)
);

O2A1O1Ixp33_ASAP7_75t_SL g1503 ( 
.A1(n_1498),
.A2(n_226),
.B(n_228),
.C(n_231),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1494),
.A2(n_232),
.B1(n_236),
.B2(n_237),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1501),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1499),
.B(n_241),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1502),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1504),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1500),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1505),
.B(n_1503),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1509),
.B(n_1003),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1507),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1506),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1512),
.Y(n_1514)
);

NOR2x1_ASAP7_75t_L g1515 ( 
.A(n_1510),
.B(n_1508),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1511),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1514),
.B(n_1513),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1515),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1515),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1516),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1518),
.Y(n_1521)
);

OAI22x1_ASAP7_75t_L g1522 ( 
.A1(n_1520),
.A2(n_253),
.B1(n_257),
.B2(n_264),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1519),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1520),
.A2(n_964),
.B1(n_271),
.B2(n_272),
.Y(n_1524)
);

OAI22x1_ASAP7_75t_L g1525 ( 
.A1(n_1517),
.A2(n_268),
.B1(n_274),
.B2(n_277),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1521),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1523),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1522),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1525),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1528),
.A2(n_1524),
.B1(n_964),
.B2(n_288),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1526),
.A2(n_290),
.B1(n_294),
.B2(n_295),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1529),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1532),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1530),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1533),
.A2(n_1527),
.B1(n_1531),
.B2(n_307),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1535),
.Y(n_1536)
);

AOI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1536),
.A2(n_1534),
.B1(n_311),
.B2(n_312),
.C(n_313),
.Y(n_1537)
);

AOI211xp5_ASAP7_75t_L g1538 ( 
.A1(n_1537),
.A2(n_323),
.B(n_329),
.C(n_330),
.Y(n_1538)
);


endmodule