module real_jpeg_17080_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_611, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_611;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_372;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_431;
wire n_357;
wire n_420;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_608;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_0),
.A2(n_21),
.B(n_607),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_0),
.B(n_608),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_1),
.A2(n_109),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_1),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_1),
.A2(n_360),
.B1(n_391),
.B2(n_394),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_1),
.A2(n_360),
.B1(n_531),
.B2(n_534),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_SL g541 ( 
.A1(n_1),
.A2(n_360),
.B1(n_542),
.B2(n_544),
.Y(n_541)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_2),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_2),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_2),
.A2(n_63),
.B1(n_94),
.B2(n_119),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_2),
.A2(n_94),
.B1(n_234),
.B2(n_239),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_2),
.A2(n_94),
.B1(n_344),
.B2(n_348),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_3),
.A2(n_352),
.B1(n_353),
.B2(n_355),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_3),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_3),
.A2(n_352),
.B1(n_416),
.B2(n_419),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_3),
.A2(n_352),
.B1(n_508),
.B2(n_513),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_3),
.A2(n_349),
.B1(n_352),
.B2(n_564),
.Y(n_563)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_4),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_4),
.Y(n_222)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_4),
.Y(n_379)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_5),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_6),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_6),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_6),
.A2(n_292),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_6),
.A2(n_292),
.B1(n_461),
.B2(n_462),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_6),
.A2(n_292),
.B1(n_518),
.B2(n_520),
.Y(n_517)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_7),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_7),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_7),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_7),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_8),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_8),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_8),
.A2(n_250),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_8),
.A2(n_250),
.B1(n_399),
.B2(n_402),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_8),
.A2(n_250),
.B1(n_478),
.B2(n_483),
.Y(n_477)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_9),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_9),
.B(n_101),
.Y(n_429)
);

OAI32xp33_ASAP7_75t_L g469 ( 
.A1(n_9),
.A2(n_29),
.A3(n_399),
.B1(n_470),
.B2(n_473),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_9),
.B(n_53),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_9),
.A2(n_216),
.B1(n_376),
.B2(n_563),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_SL g581 ( 
.A1(n_9),
.A2(n_326),
.B1(n_582),
.B2(n_583),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_10),
.A2(n_56),
.B1(n_62),
.B2(n_63),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_10),
.A2(n_62),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_10),
.A2(n_62),
.B1(n_224),
.B2(n_229),
.Y(n_223)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_11),
.Y(n_608)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_12),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_12),
.Y(n_146)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_12),
.Y(n_228)
);

BUFx4f_ASAP7_75t_L g347 ( 
.A(n_12),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_13),
.A2(n_103),
.B1(n_108),
.B2(n_112),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_13),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_13),
.A2(n_112),
.B1(n_117),
.B2(n_122),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_13),
.A2(n_112),
.B1(n_199),
.B2(n_202),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_13),
.A2(n_112),
.B1(n_277),
.B2(n_280),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_14),
.A2(n_130),
.B1(n_132),
.B2(n_134),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_14),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_14),
.A2(n_134),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_14),
.A2(n_134),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_L g337 ( 
.A1(n_14),
.A2(n_134),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_16),
.A2(n_92),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_16),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_16),
.A2(n_176),
.B1(n_297),
.B2(n_299),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_16),
.A2(n_176),
.B1(n_370),
.B2(n_372),
.Y(n_369)
);

OAI22x1_ASAP7_75t_SL g421 ( 
.A1(n_16),
.A2(n_176),
.B1(n_422),
.B2(n_424),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_17),
.Y(n_154)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_17),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_17),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_17),
.Y(n_374)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_17),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_19),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g354 ( 
.A(n_19),
.Y(n_354)
);

BUFx5_ASAP7_75t_L g357 ( 
.A(n_19),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_182),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_181),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_166),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_25),
.B(n_166),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g610 ( 
.A(n_25),
.Y(n_610)
);

FAx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_67),
.CI(n_113),
.CON(n_25),
.SN(n_25)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_53),
.B(n_54),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_27),
.A2(n_53),
.B1(n_205),
.B2(n_211),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_27),
.A2(n_53),
.B1(n_311),
.B2(n_390),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_27),
.A2(n_53),
.B1(n_390),
.B2(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_28),
.A2(n_55),
.B1(n_116),
.B2(n_126),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_28),
.A2(n_116),
.B1(n_126),
.B2(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_28),
.A2(n_126),
.B1(n_206),
.B2(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_28),
.A2(n_126),
.B1(n_310),
.B2(n_316),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_28),
.A2(n_126),
.B1(n_296),
.B2(n_316),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_28),
.A2(n_126),
.B1(n_415),
.B2(n_581),
.Y(n_580)
);

AO21x2_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_38),
.B(n_46),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_35),
.Y(n_312)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_37),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_43),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_45),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_47),
.Y(n_165)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_47),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_47),
.Y(n_371)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_51),
.Y(n_203)
);

INVx6_ASAP7_75t_L g491 ( 
.A(n_51),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_52),
.Y(n_401)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_66),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_66),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_90),
.B1(n_100),
.B2(n_102),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_68),
.A2(n_100),
.B1(n_129),
.B2(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_68),
.A2(n_80),
.B1(n_173),
.B2(n_248),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_L g288 ( 
.A1(n_68),
.A2(n_80),
.B1(n_248),
.B2(n_289),
.Y(n_288)
);

OAI22x1_ASAP7_75t_SL g381 ( 
.A1(n_68),
.A2(n_100),
.B1(n_289),
.B2(n_359),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_69),
.A2(n_91),
.B1(n_101),
.B2(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_69),
.A2(n_101),
.B1(n_351),
.B2(n_358),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_69),
.A2(n_101),
.B1(n_351),
.B2(n_396),
.Y(n_395)
);

OA21x2_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_77),
.B(n_80),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_77),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_78),
.Y(n_328)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

AOI22x1_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_87),
.Y(n_210)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_92),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_108),
.B(n_326),
.Y(n_325)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g291 ( 
.A(n_111),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_127),
.C(n_135),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_114),
.A2(n_115),
.B1(n_135),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_119),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_119),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_120),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_121),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_124),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_124),
.Y(n_394)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_125),
.Y(n_393)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_125),
.Y(n_587)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_135),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_171),
.C(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_135),
.B(n_179),
.Y(n_193)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_149),
.B(n_161),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_136),
.A2(n_149),
.B1(n_161),
.B2(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_136),
.B(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_136),
.A2(n_149),
.B1(n_398),
.B2(n_406),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_136),
.A2(n_149),
.B1(n_505),
.B2(n_507),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_136),
.A2(n_149),
.B1(n_507),
.B2(n_530),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_136),
.A2(n_149),
.B1(n_460),
.B2(n_530),
.Y(n_589)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_137),
.A2(n_198),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_137),
.A2(n_232),
.B1(n_265),
.B2(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_137),
.A2(n_232),
.B1(n_459),
.B2(n_466),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_137),
.B(n_326),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_138),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_142),
.B1(n_144),
.B2(n_147),
.Y(n_138)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_143),
.Y(n_220)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_143),
.Y(n_230)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_143),
.Y(n_279)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_143),
.Y(n_349)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_143),
.Y(n_423)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_143),
.Y(n_482)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_146),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_146),
.Y(n_543)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_146),
.Y(n_560)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_148),
.Y(n_499)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_149),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_149),
.B(n_264),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_155),
.B1(n_158),
.B2(n_160),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_154),
.Y(n_465)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_158),
.Y(n_493)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_165),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_177),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_170),
.B1(n_171),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_303),
.B(n_604),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_253),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g604 ( 
.A1(n_187),
.A2(n_605),
.B(n_606),
.Y(n_604)
);

NOR2x1_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_188),
.B(n_191),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_212),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_192),
.A2(n_194),
.B1(n_195),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_192),
.Y(n_302)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_195),
.A2(n_196),
.B(n_204),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_204),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_199),
.Y(n_506)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_201),
.Y(n_461)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_212),
.B(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_244),
.B1(n_252),
.B2(n_611),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_213),
.A2(n_214),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_231),
.Y(n_214)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_215),
.A2(n_246),
.B1(n_247),
.B2(n_252),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_215),
.A2(n_231),
.B1(n_252),
.B2(n_441),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_221),
.B(n_223),
.Y(n_215)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_216),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_216),
.A2(n_336),
.B1(n_341),
.B2(n_343),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_216),
.A2(n_276),
.B1(n_343),
.B2(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_216),
.A2(n_285),
.B1(n_517),
.B2(n_525),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_216),
.A2(n_541),
.B1(n_563),
.B2(n_567),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_219),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_219),
.Y(n_342)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_220),
.Y(n_338)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_220),
.Y(n_492)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g568 ( 
.A(n_222),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_223),
.Y(n_286)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_226),
.Y(n_340)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_226),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_227),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_228),
.Y(n_283)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_231),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_233),
.Y(n_272)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_238),
.Y(n_243)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_238),
.Y(n_405)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_249),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_300),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_254),
.B(n_300),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_259),
.C(n_261),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_256),
.B(n_260),
.Y(n_435)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_261),
.B(n_435),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_287),
.C(n_295),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_262),
.B(n_439),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_271),
.B(n_273),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_263),
.B(n_271),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_273),
.B(n_365),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_284),
.B2(n_286),
.Y(n_273)
);

AOI22x1_ASAP7_75t_SL g420 ( 
.A1(n_274),
.A2(n_337),
.B1(n_421),
.B2(n_427),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_274),
.A2(n_377),
.B1(n_421),
.B2(n_477),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_274),
.A2(n_540),
.B1(n_547),
.B2(n_548),
.Y(n_539)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_288),
.B(n_295),
.Y(n_439)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_291),
.Y(n_294)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_450),
.B(n_599),
.Y(n_303)
);

NAND3xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_433),
.C(n_445),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_383),
.B(n_407),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_306),
.B(n_383),
.C(n_601),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_363),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_307),
.B(n_364),
.C(n_366),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_323),
.C(n_350),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_309),
.B(n_350),
.Y(n_386)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx6_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_321),
.Y(n_333)
);

INVx8_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_323),
.B(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_335),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_324),
.B(n_335),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_327),
.B1(n_333),
.B2(n_334),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_SL g396 ( 
.A1(n_325),
.A2(n_326),
.B(n_353),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_326),
.B(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_326),
.B(n_495),
.Y(n_494)
);

OAI21xp33_ASAP7_75t_SL g505 ( 
.A1(n_326),
.A2(n_494),
.B(n_506),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_326),
.B(n_428),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_346),
.Y(n_483)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_347),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_347),
.Y(n_519)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx12f_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_357),
.Y(n_362)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_380),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_367),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_375),
.Y(n_367)
);

XOR2x2_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_375),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_369),
.Y(n_406)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_373),
.Y(n_535)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_376),
.Y(n_547)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_378),
.Y(n_428)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_382),
.C(n_444),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_387),
.C(n_388),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_384),
.A2(n_385),
.B1(n_431),
.B2(n_432),
.Y(n_430)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_387),
.B(n_388),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_395),
.C(n_397),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_397),
.Y(n_410)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_410),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_398),
.Y(n_466)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_404),
.Y(n_474)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_430),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_408),
.B(n_430),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.C(n_412),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_409),
.B(n_453),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_411),
.B(n_412),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_420),
.C(n_429),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_413),
.B(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx2_ASAP7_75t_SL g417 ( 
.A(n_418),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_420),
.B(n_429),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_422),
.Y(n_564)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx6_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_431),
.Y(n_432)
);

A2O1A1O1Ixp25_ASAP7_75t_L g599 ( 
.A1(n_433),
.A2(n_445),
.B(n_600),
.C(n_602),
.D(n_603),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_436),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_434),
.B(n_436),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_440),
.C(n_442),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_437),
.A2(n_438),
.B1(n_440),
.B2(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_440),
.Y(n_448)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_443),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_449),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_446),
.B(n_449),
.Y(n_602)
);

AOI21x1_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_484),
.B(n_598),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_454),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_452),
.B(n_454),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_458),
.C(n_467),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_455),
.A2(n_456),
.B1(n_593),
.B2(n_594),
.Y(n_592)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_458),
.A2(n_467),
.B1(n_468),
.B2(n_595),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_458),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx5_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_475),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_469),
.A2(n_475),
.B1(n_476),
.B2(n_577),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_469),
.Y(n_577)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_474),
.Y(n_495)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_477),
.Y(n_525)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_591),
.B(n_597),
.Y(n_484)
);

AOI21x1_ASAP7_75t_SL g485 ( 
.A1(n_486),
.A2(n_573),
.B(n_590),
.Y(n_485)
);

OAI21x1_ASAP7_75t_L g486 ( 
.A1(n_487),
.A2(n_537),
.B(n_572),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_515),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_488),
.B(n_515),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_503),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_489),
.A2(n_503),
.B1(n_504),
.B2(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_489),
.Y(n_550)
);

OAI32xp33_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_492),
.A3(n_493),
.B1(n_494),
.B2(n_496),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_500),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_512),
.Y(n_514)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_512),
.Y(n_533)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_526),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_516),
.B(n_528),
.C(n_536),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_517),
.Y(n_548)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_528),
.B1(n_529),
.B2(n_536),
.Y(n_526)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_527),
.Y(n_536)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_538),
.A2(n_551),
.B(n_571),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_549),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_539),
.B(n_549),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_546),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_552),
.A2(n_565),
.B(n_570),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_562),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_561),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_566),
.B(n_569),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_566),
.B(n_569),
.Y(n_570)
);

INVx6_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_574),
.B(n_575),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_574),
.B(n_575),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_578),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_576),
.B(n_579),
.C(n_589),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_579),
.A2(n_580),
.B1(n_588),
.B2(n_589),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

NOR2xp67_ASAP7_75t_SL g591 ( 
.A(n_592),
.B(n_596),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_592),
.B(n_596),
.Y(n_597)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);


endmodule