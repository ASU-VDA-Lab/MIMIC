module real_jpeg_29404_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_0),
.A2(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_105)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_2),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_2),
.A2(n_58),
.B1(n_67),
.B2(n_68),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_2),
.A2(n_25),
.B1(n_29),
.B2(n_58),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_3),
.A2(n_25),
.B1(n_29),
.B2(n_41),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_4),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_5),
.A2(n_25),
.B1(n_29),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_8),
.A2(n_67),
.B1(n_68),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_8),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_8),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_72),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_8),
.A2(n_25),
.B1(n_29),
.B2(n_72),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_9),
.A2(n_67),
.B1(n_68),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_9),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_74),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_9),
.A2(n_25),
.B1(n_29),
.B2(n_74),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_10),
.A2(n_77),
.B1(n_78),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_10),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_10),
.A2(n_67),
.B1(n_68),
.B2(n_86),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_86),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_10),
.A2(n_25),
.B1(n_29),
.B2(n_86),
.Y(n_184)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_12),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_12),
.B(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_12),
.B(n_67),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g137 ( 
.A1(n_12),
.A2(n_67),
.B(n_133),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_79),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_12),
.A2(n_25),
.B(n_30),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_12),
.B(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_12),
.A2(n_43),
.B1(n_51),
.B2(n_184),
.Y(n_186)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_15),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_123),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_106),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_87),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_42),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_36),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_24),
.A2(n_38),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_24),
.A2(n_38),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_24),
.A2(n_38),
.B1(n_140),
.B2(n_159),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_24),
.B(n_79),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_24)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_28),
.A2(n_33),
.B(n_79),
.C(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_29),
.B(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_32),
.A2(n_33),
.B1(n_65),
.B2(n_66),
.Y(n_70)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_32),
.A2(n_68),
.A3(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_131)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g134 ( 
.A(n_33),
.B(n_65),
.Y(n_134)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_56),
.B(n_59),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_38),
.A2(n_141),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_47),
.B(n_49),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_43),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_43),
.A2(n_118),
.B1(n_176),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_44),
.B(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_44),
.A2(n_50),
.B(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_44),
.A2(n_45),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_45),
.B(n_130),
.Y(n_171)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_51),
.B(n_79),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.C(n_75),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_57),
.B(n_60),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_62)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_63),
.A2(n_70),
.B1(n_71),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_63),
.A2(n_70),
.B1(n_114),
.B2(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_64)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_68),
.B1(n_81),
.B2(n_82),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_81),
.Y(n_103)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_76),
.B1(n_83),
.B2(n_103),
.Y(n_102)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_75),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.CON(n_76),
.SN(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_81),
.B(n_83),
.C(n_84),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_81),
.Y(n_83)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_101),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_104),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_112),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_107),
.A2(n_108),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_112),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.C(n_117),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_117),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_199),
.B(n_205),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_152),
.B(n_198),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_142),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_126),
.B(n_142),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_135),
.C(n_138),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_127),
.A2(n_128),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_131),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_149),
.C(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_192),
.B(n_197),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_172),
.B(n_191),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_162),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_155),
.B(n_162),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_179),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_169),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_168),
.C(n_169),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_170),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_180),
.B(n_190),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_178),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_185),
.B(n_189),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_183),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_193),
.B(n_194),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_200),
.B(n_201),
.Y(n_205)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);


endmodule