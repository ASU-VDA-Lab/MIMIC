module real_jpeg_15409_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OA22x2_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_4),
.B1(n_15),
.B2(n_16),
.Y(n_14)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_0),
.B(n_3),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g9 ( 
.A(n_1),
.B(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

OAI322xp33_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_15),
.A3(n_20),
.B1(n_21),
.B2(n_22),
.C1(n_23),
.C2(n_24),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_3),
.B(n_15),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_3),
.A2(n_11),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

AOI321xp33_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_13),
.A3(n_17),
.B1(n_18),
.B2(n_19),
.C(n_25),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

AND2x2_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_12),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_14),
.Y(n_13)
);

INVx2_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_18),
.B(n_33),
.Y(n_32)
);

OAI221xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.C(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);


endmodule