module fake_netlist_6_3092_n_2678 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_533, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_546, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2678);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_533;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_546;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2678;

wire n_992;
wire n_2542;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_558;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_622;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_2307;
wire n_2069;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_683;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2545;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2511;
wire n_2475;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2617;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2420;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_1332;
wire n_2670;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_2671;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_752;
wire n_2649;
wire n_944;
wire n_2034;
wire n_1028;
wire n_576;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2471;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_241),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_70),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_543),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_420),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_168),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_422),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_332),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_445),
.Y(n_556)
);

BUFx8_ASAP7_75t_SL g557 ( 
.A(n_90),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_528),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_342),
.Y(n_559)
);

BUFx10_ASAP7_75t_L g560 ( 
.A(n_34),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_449),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_33),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_108),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_353),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_489),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_110),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_248),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_328),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_139),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_268),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_271),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_446),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_546),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_57),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_320),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_330),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_204),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_458),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_132),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_515),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_2),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_202),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_510),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_339),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_434),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_44),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_188),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_17),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_259),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_481),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_394),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_540),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_397),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_15),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_128),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_490),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_545),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_433),
.Y(n_598)
);

BUFx5_ASAP7_75t_L g599 ( 
.A(n_75),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_313),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_379),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_488),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_268),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_415),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_453),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_512),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_15),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_243),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_330),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_177),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_236),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_361),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_313),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_262),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_7),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_343),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_301),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_288),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_226),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_389),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_537),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_95),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_76),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_542),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_322),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_269),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_16),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_127),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_279),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_466),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_436),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_526),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_401),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_426),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_60),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_531),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_346),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_3),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_30),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_133),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_108),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_432),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_202),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_370),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_118),
.Y(n_645)
);

BUFx5_ASAP7_75t_L g646 ( 
.A(n_460),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_388),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_544),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_156),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_141),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_500),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_412),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_344),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_497),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_100),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_413),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_310),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_465),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_398),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_456),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_338),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_145),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_511),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_354),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_476),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_211),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_498),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_509),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_532),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_10),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_333),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_533),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_307),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_381),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_522),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_144),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_93),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_505),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_345),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_301),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_117),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_539),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_373),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_410),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_85),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_201),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_424),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_494),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_152),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_502),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_78),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_442),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_255),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_326),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_455),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_159),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_469),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_471),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_486),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_81),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_285),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_260),
.Y(n_702)
);

BUFx10_ASAP7_75t_L g703 ( 
.A(n_487),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_37),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_463),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_54),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_479),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_470),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_506),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_495),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_294),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_480),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_232),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_97),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_356),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_337),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_255),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_419),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_452),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_541),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_318),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_414),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_100),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_253),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_22),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_31),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_201),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_536),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_277),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_9),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_369),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_180),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_357),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_341),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_99),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_477),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_193),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_54),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_145),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_350),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_270),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_457),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_212),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_416),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_295),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_72),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_402),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_314),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_28),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_1),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_274),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_523),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_41),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_535),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_437),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_474),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_58),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_530),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_170),
.Y(n_759)
);

BUFx10_ASAP7_75t_L g760 ( 
.A(n_529),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_137),
.Y(n_761)
);

CKINVDCx14_ASAP7_75t_R g762 ( 
.A(n_125),
.Y(n_762)
);

BUFx10_ASAP7_75t_L g763 ( 
.A(n_79),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_309),
.Y(n_764)
);

BUFx2_ASAP7_75t_SL g765 ( 
.A(n_146),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_339),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_24),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_85),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_411),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_336),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_325),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_122),
.Y(n_772)
);

CKINVDCx6p67_ASAP7_75t_R g773 ( 
.A(n_97),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_538),
.Y(n_774)
);

BUFx10_ASAP7_75t_L g775 ( 
.A(n_84),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_326),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_150),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_340),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_322),
.Y(n_779)
);

BUFx5_ASAP7_75t_L g780 ( 
.A(n_69),
.Y(n_780)
);

CKINVDCx16_ASAP7_75t_R g781 ( 
.A(n_104),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_534),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_491),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_165),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_266),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_296),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_165),
.Y(n_787)
);

BUFx10_ASAP7_75t_L g788 ( 
.A(n_362),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_69),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_429),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_516),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_599),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_599),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_599),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_577),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_557),
.Y(n_796)
);

INVxp33_ASAP7_75t_L g797 ( 
.A(n_768),
.Y(n_797)
);

CKINVDCx14_ASAP7_75t_R g798 ( 
.A(n_762),
.Y(n_798)
);

INVxp67_ASAP7_75t_SL g799 ( 
.A(n_705),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_599),
.Y(n_800)
);

INVxp67_ASAP7_75t_SL g801 ( 
.A(n_596),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_599),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_557),
.Y(n_803)
);

CKINVDCx14_ASAP7_75t_R g804 ( 
.A(n_762),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_599),
.Y(n_805)
);

CKINVDCx16_ASAP7_75t_R g806 ( 
.A(n_781),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_780),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_552),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_556),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_558),
.Y(n_810)
);

INVxp33_ASAP7_75t_SL g811 ( 
.A(n_574),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_780),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_780),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_586),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_561),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_780),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_623),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_780),
.Y(n_818)
);

INVxp33_ASAP7_75t_SL g819 ( 
.A(n_694),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_620),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_780),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_577),
.Y(n_822)
);

CKINVDCx16_ASAP7_75t_R g823 ( 
.A(n_699),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_585),
.Y(n_824)
);

CKINVDCx16_ASAP7_75t_R g825 ( 
.A(n_699),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_646),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_683),
.B(n_0),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_771),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_587),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_587),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_614),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_635),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_611),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_646),
.Y(n_834)
);

INVxp33_ASAP7_75t_SL g835 ( 
.A(n_549),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_611),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_693),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_693),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_711),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_711),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_646),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_735),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_735),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_745),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_745),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_680),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_550),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_579),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_579),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_591),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_560),
.Y(n_851)
);

INVxp33_ASAP7_75t_SL g852 ( 
.A(n_563),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_686),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_579),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_592),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_620),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_560),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_696),
.Y(n_858)
);

INVxp33_ASAP7_75t_L g859 ( 
.A(n_562),
.Y(n_859)
);

INVxp33_ASAP7_75t_SL g860 ( 
.A(n_765),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_579),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_641),
.Y(n_862)
);

CKINVDCx16_ASAP7_75t_R g863 ( 
.A(n_560),
.Y(n_863)
);

BUFx8_ASAP7_75t_SL g864 ( 
.A(n_717),
.Y(n_864)
);

INVxp33_ASAP7_75t_SL g865 ( 
.A(n_570),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_641),
.Y(n_866)
);

INVxp67_ASAP7_75t_L g867 ( 
.A(n_575),
.Y(n_867)
);

INVxp33_ASAP7_75t_SL g868 ( 
.A(n_571),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_575),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_641),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_748),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_646),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_581),
.Y(n_873)
);

CKINVDCx14_ASAP7_75t_R g874 ( 
.A(n_551),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_641),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_726),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_575),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_582),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_726),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_654),
.Y(n_880)
);

CKINVDCx14_ASAP7_75t_R g881 ( 
.A(n_551),
.Y(n_881)
);

INVxp67_ASAP7_75t_SL g882 ( 
.A(n_654),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_726),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_726),
.Y(n_884)
);

INVxp67_ASAP7_75t_SL g885 ( 
.A(n_774),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_733),
.Y(n_886)
);

INVxp33_ASAP7_75t_SL g887 ( 
.A(n_584),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_751),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_757),
.Y(n_889)
);

INVxp33_ASAP7_75t_SL g890 ( 
.A(n_588),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_751),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_751),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_751),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_848),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_849),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_820),
.B(n_774),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_808),
.B(n_554),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_882),
.B(n_683),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_886),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_886),
.Y(n_900)
);

AOI22x1_ASAP7_75t_SL g901 ( 
.A1(n_814),
.A2(n_789),
.B1(n_778),
.B2(n_594),
.Y(n_901)
);

BUFx8_ASAP7_75t_L g902 ( 
.A(n_817),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_809),
.B(n_583),
.Y(n_903)
);

NOR2x1_ASAP7_75t_L g904 ( 
.A(n_827),
.B(n_564),
.Y(n_904)
);

CKINVDCx11_ASAP7_75t_R g905 ( 
.A(n_814),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_854),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_886),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_798),
.B(n_551),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_886),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_810),
.B(n_756),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_861),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_815),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_885),
.B(n_756),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_856),
.Y(n_914)
);

BUFx12f_ASAP7_75t_L g915 ( 
.A(n_796),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_811),
.A2(n_819),
.B1(n_806),
.B2(n_801),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_793),
.A2(n_572),
.B(n_565),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_824),
.B(n_573),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_798),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_839),
.Y(n_920)
);

AND2x2_ASAP7_75t_SL g921 ( 
.A(n_823),
.B(n_733),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_856),
.B(n_880),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_850),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_862),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_811),
.A2(n_589),
.B1(n_603),
.B2(n_595),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_855),
.B(n_578),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_880),
.B(n_580),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_793),
.Y(n_928)
);

BUFx8_ASAP7_75t_L g929 ( 
.A(n_877),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_822),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_866),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_870),
.Y(n_932)
);

NOR2x1_ASAP7_75t_L g933 ( 
.A(n_875),
.B(n_590),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_876),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_879),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_799),
.B(n_597),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_883),
.Y(n_937)
);

BUFx8_ASAP7_75t_L g938 ( 
.A(n_877),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_884),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_888),
.Y(n_940)
);

INVx5_ASAP7_75t_L g941 ( 
.A(n_826),
.Y(n_941)
);

INVx5_ASAP7_75t_L g942 ( 
.A(n_826),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_891),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_892),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_864),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_893),
.Y(n_946)
);

INVx5_ASAP7_75t_L g947 ( 
.A(n_834),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_792),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_804),
.B(n_874),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_819),
.A2(n_608),
.B1(n_613),
.B2(n_610),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_794),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_800),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_802),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_805),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_807),
.Y(n_955)
);

OA21x2_ASAP7_75t_L g956 ( 
.A1(n_812),
.A2(n_606),
.B(n_604),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_813),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_834),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_816),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_898),
.B(n_804),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_928),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_928),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_948),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_952),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_917),
.A2(n_904),
.B(n_956),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_929),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_920),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_929),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_948),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_953),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_929),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_898),
.B(n_874),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_952),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_953),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_902),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_952),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_957),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_952),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_913),
.B(n_859),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_954),
.Y(n_980)
);

INVx4_ASAP7_75t_SL g981 ( 
.A(n_954),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_954),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_954),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_958),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_913),
.B(n_859),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_955),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_914),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_902),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_913),
.B(n_795),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_R g990 ( 
.A(n_912),
.B(n_881),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_905),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_955),
.Y(n_992)
);

NOR2xp67_ASAP7_75t_L g993 ( 
.A(n_912),
.B(n_847),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_955),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_955),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_938),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_951),
.Y(n_997)
);

CKINVDCx16_ASAP7_75t_R g998 ( 
.A(n_919),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_957),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_938),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_959),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_938),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_959),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_905),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_898),
.B(n_881),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_930),
.Y(n_1006)
);

CKINVDCx8_ASAP7_75t_R g1007 ( 
.A(n_923),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_899),
.Y(n_1008)
);

INVxp67_ASAP7_75t_L g1009 ( 
.A(n_914),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_910),
.B(n_835),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_923),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_899),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_900),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_945),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_900),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_945),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_930),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_922),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_902),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_932),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_907),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_894),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_895),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_918),
.B(n_852),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_906),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_932),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_911),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_919),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_915),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_924),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_932),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_931),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_935),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_946),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_907),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_922),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_922),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_932),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_915),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_909),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_909),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_934),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_896),
.B(n_795),
.Y(n_1043)
);

NAND2xp33_ASAP7_75t_R g1044 ( 
.A(n_908),
.B(n_890),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_896),
.B(n_829),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_934),
.Y(n_1046)
);

OA21x2_ASAP7_75t_L g1047 ( 
.A1(n_927),
.A2(n_821),
.B(n_818),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_896),
.B(n_933),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_921),
.B(n_865),
.Y(n_1049)
);

OR2x6_ASAP7_75t_L g1050 ( 
.A(n_975),
.B(n_803),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_979),
.B(n_949),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1045),
.A2(n_979),
.B1(n_985),
.B2(n_1043),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_1024),
.B(n_868),
.Y(n_1053)
);

INVx4_ASAP7_75t_L g1054 ( 
.A(n_973),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_985),
.B(n_921),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_962),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_1010),
.B(n_887),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_962),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1036),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1037),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_1045),
.B(n_936),
.C(n_926),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1018),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1047),
.A2(n_956),
.B1(n_958),
.B2(n_860),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_962),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_989),
.B(n_956),
.C(n_903),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_1008),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_961),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1022),
.Y(n_1068)
);

AND2x6_ASAP7_75t_L g1069 ( 
.A(n_1043),
.B(n_733),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_984),
.B(n_897),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_973),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_L g1072 ( 
.A(n_1049),
.B(n_950),
.C(n_925),
.Y(n_1072)
);

INVx4_ASAP7_75t_L g1073 ( 
.A(n_973),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_967),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_963),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_963),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_969),
.Y(n_1077)
);

INVxp67_ASAP7_75t_SL g1078 ( 
.A(n_984),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_984),
.B(n_860),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_989),
.B(n_841),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_973),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_969),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_1009),
.B(n_890),
.Y(n_1083)
);

AND2x6_ASAP7_75t_L g1084 ( 
.A(n_1048),
.B(n_733),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_998),
.B(n_825),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_1048),
.B(n_916),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_972),
.A2(n_828),
.B1(n_637),
.B2(n_779),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_1048),
.B(n_863),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_993),
.B(n_602),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1023),
.Y(n_1090)
);

OR2x6_ASAP7_75t_L g1091 ( 
.A(n_988),
.B(n_960),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_970),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1025),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_970),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1027),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1030),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1032),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_987),
.B(n_873),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1033),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_974),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_1005),
.B(n_1006),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1047),
.A2(n_637),
.B1(n_779),
.B2(n_562),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_990),
.B(n_630),
.Y(n_1103)
);

CKINVDCx16_ASAP7_75t_R g1104 ( 
.A(n_1028),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1047),
.B(n_841),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1034),
.Y(n_1106)
);

NAND2xp33_ASAP7_75t_L g1107 ( 
.A(n_997),
.B(n_646),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1017),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_1044),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_1007),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_977),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_977),
.B(n_872),
.Y(n_1112)
);

INVxp67_ASAP7_75t_L g1113 ( 
.A(n_999),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1003),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_980),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1003),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1008),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_1028),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_1011),
.B(n_878),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_1012),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1001),
.A2(n_787),
.B1(n_555),
.B2(n_559),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_1012),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_1011),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1013),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1013),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_964),
.B(n_872),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1007),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1015),
.Y(n_1128)
);

BUFx10_ASAP7_75t_L g1129 ( 
.A(n_1014),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_991),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1015),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1021),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1021),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1035),
.Y(n_1134)
);

XNOR2xp5_ASAP7_75t_L g1135 ( 
.A(n_991),
.B(n_831),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_1035),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_966),
.B(n_797),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_966),
.B(n_797),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1040),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_976),
.A2(n_621),
.B1(n_642),
.B2(n_636),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_968),
.B(n_831),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1040),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1041),
.Y(n_1143)
);

BUFx10_ASAP7_75t_L g1144 ( 
.A(n_1014),
.Y(n_1144)
);

AND2x6_ASAP7_75t_L g1145 ( 
.A(n_1041),
.B(n_644),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1046),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_968),
.B(n_782),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_1046),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_980),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_971),
.B(n_783),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_971),
.B(n_832),
.Y(n_1151)
);

OAI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_996),
.A2(n_691),
.B1(n_770),
.B2(n_689),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_978),
.B(n_941),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_980),
.Y(n_1154)
);

CKINVDCx6p67_ASAP7_75t_R g1155 ( 
.A(n_1004),
.Y(n_1155)
);

BUFx4f_ASAP7_75t_L g1156 ( 
.A(n_986),
.Y(n_1156)
);

AO22x2_ASAP7_75t_L g1157 ( 
.A1(n_992),
.A2(n_901),
.B1(n_628),
.B2(n_649),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_994),
.B(n_941),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1000),
.B(n_846),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_980),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_982),
.Y(n_1161)
);

AND2x2_ASAP7_75t_SL g1162 ( 
.A(n_1000),
.B(n_787),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_965),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1002),
.B(n_624),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_965),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1038),
.Y(n_1166)
);

INVxp33_ASAP7_75t_L g1167 ( 
.A(n_1004),
.Y(n_1167)
);

NAND2xp33_ASAP7_75t_SL g1168 ( 
.A(n_1002),
.B(n_618),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1042),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_982),
.B(n_658),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_982),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_995),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_982),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1016),
.B(n_851),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1016),
.B(n_857),
.Y(n_1175)
);

INVxp67_ASAP7_75t_SL g1176 ( 
.A(n_983),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_983),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_983),
.Y(n_1178)
);

INVx5_ASAP7_75t_L g1179 ( 
.A(n_983),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1019),
.A2(n_566),
.B1(n_567),
.B2(n_553),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_1029),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_1019),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_SL g1183 ( 
.A(n_1029),
.B(n_626),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1039),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_1039),
.B(n_867),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1059),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1114),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1116),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1078),
.B(n_1020),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1067),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1072),
.A2(n_675),
.B1(n_682),
.B2(n_672),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1066),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1053),
.B(n_869),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1062),
.B(n_830),
.Y(n_1194)
);

NAND2x1p5_ASAP7_75t_L g1195 ( 
.A(n_1110),
.B(n_1020),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1060),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1181),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1057),
.B(n_846),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_L g1199 ( 
.A(n_1119),
.B(n_616),
.C(n_615),
.Y(n_1199)
);

CKINVDCx16_ASAP7_75t_R g1200 ( 
.A(n_1104),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1075),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1078),
.B(n_1020),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1076),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1074),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_1127),
.B(n_1020),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1077),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1071),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1070),
.B(n_1026),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1082),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1092),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1094),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1070),
.B(n_1026),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1100),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1051),
.B(n_833),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1066),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1098),
.Y(n_1216)
);

INVx5_ASAP7_75t_L g1217 ( 
.A(n_1091),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1108),
.B(n_836),
.Y(n_1218)
);

CKINVDCx8_ASAP7_75t_R g1219 ( 
.A(n_1123),
.Y(n_1219)
);

INVxp33_ASAP7_75t_SL g1220 ( 
.A(n_1135),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1155),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1109),
.B(n_853),
.Y(n_1222)
);

BUFx4f_ASAP7_75t_L g1223 ( 
.A(n_1091),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1129),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1055),
.B(n_853),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1068),
.B(n_837),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1090),
.B(n_838),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1052),
.B(n_858),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1111),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1093),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1120),
.Y(n_1231)
);

INVx4_ASAP7_75t_SL g1232 ( 
.A(n_1084),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1085),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1079),
.B(n_1026),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1071),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1095),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1096),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1097),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1099),
.B(n_840),
.Y(n_1239)
);

AND2x6_ASAP7_75t_L g1240 ( 
.A(n_1163),
.B(n_684),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1052),
.B(n_858),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1106),
.B(n_842),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_SL g1243 ( 
.A1(n_1162),
.A2(n_871),
.B1(n_889),
.B2(n_864),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_L g1244 ( 
.A(n_1072),
.B(n_619),
.C(n_617),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1117),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_1071),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1124),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1174),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1134),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1142),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1113),
.B(n_843),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1120),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1081),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1122),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1136),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1125),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1083),
.B(n_871),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1065),
.A2(n_690),
.B1(n_692),
.B2(n_687),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1128),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1109),
.B(n_889),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1137),
.A2(n_760),
.B1(n_788),
.B2(n_703),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_1118),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1148),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1113),
.B(n_844),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1081),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1079),
.B(n_1026),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1146),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1131),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1130),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1132),
.Y(n_1270)
);

AND2x6_ASAP7_75t_L g1271 ( 
.A(n_1165),
.B(n_697),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1086),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1089),
.B(n_773),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1091),
.B(n_845),
.Y(n_1274)
);

AO22x2_ASAP7_75t_L g1275 ( 
.A1(n_1180),
.A2(n_568),
.B1(n_576),
.B2(n_569),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1133),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1139),
.Y(n_1277)
);

AO22x2_ASAP7_75t_L g1278 ( 
.A1(n_1180),
.A2(n_607),
.B1(n_609),
.B2(n_600),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1129),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1143),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1061),
.B(n_981),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1126),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1081),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1175),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1148),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1126),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1061),
.B(n_981),
.Y(n_1287)
);

AO22x2_ASAP7_75t_L g1288 ( 
.A1(n_1087),
.A2(n_627),
.B1(n_643),
.B2(n_625),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1161),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1144),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1056),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1101),
.B(n_1031),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1166),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1169),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1080),
.B(n_1031),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1149),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1138),
.B(n_763),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1050),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1172),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1080),
.B(n_1031),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1156),
.B(n_981),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1112),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1058),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1112),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1064),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_SL g1306 ( 
.A1(n_1141),
.A2(n_676),
.B1(n_737),
.B2(n_657),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1171),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_1144),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1173),
.Y(n_1309)
);

NAND2x1p5_ASAP7_75t_L g1310 ( 
.A(n_1179),
.B(n_1031),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1178),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1184),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1160),
.Y(n_1313)
);

AND2x6_ASAP7_75t_L g1314 ( 
.A(n_1105),
.B(n_698),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1161),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1176),
.B(n_981),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1088),
.B(n_1176),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1161),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1182),
.B(n_666),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1105),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1065),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1063),
.B(n_709),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1087),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1145),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1145),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1145),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1183),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1145),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1151),
.A2(n_714),
.B1(n_743),
.B2(n_679),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1164),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1156),
.B(n_593),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1054),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1153),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1054),
.Y(n_1334)
);

NAND2x1p5_ASAP7_75t_L g1335 ( 
.A(n_1179),
.B(n_934),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1170),
.A2(n_712),
.B1(n_715),
.B2(n_710),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1073),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1103),
.B(n_622),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1073),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1050),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1102),
.B(n_740),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1102),
.B(n_754),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1115),
.B(n_755),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1179),
.Y(n_1344)
);

INVx4_ASAP7_75t_L g1345 ( 
.A(n_1115),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1153),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1154),
.B(n_598),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1154),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1158),
.Y(n_1349)
);

INVx6_ASAP7_75t_L g1350 ( 
.A(n_1050),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1177),
.B(n_601),
.Y(n_1351)
);

NAND3xp33_ASAP7_75t_L g1352 ( 
.A(n_1168),
.B(n_638),
.C(n_629),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1177),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1158),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1084),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1147),
.B(n_677),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1084),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1107),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1084),
.B(n_758),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1150),
.B(n_1159),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1069),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1069),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1152),
.B(n_639),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1069),
.B(n_769),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1157),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1185),
.Y(n_1366)
);

NAND2xp33_ASAP7_75t_L g1367 ( 
.A(n_1140),
.B(n_646),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1152),
.B(n_640),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_SL g1369 ( 
.A(n_1167),
.B(n_703),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1121),
.B(n_605),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1121),
.B(n_612),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1157),
.Y(n_1372)
);

OR2x6_ASAP7_75t_L g1373 ( 
.A(n_1185),
.B(n_681),
.Y(n_1373)
);

INVxp67_ASAP7_75t_L g1374 ( 
.A(n_1185),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1055),
.B(n_631),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1078),
.B(n_632),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1114),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1114),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1053),
.B(n_763),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1062),
.B(n_701),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1114),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1114),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1059),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1272),
.A2(n_634),
.B1(n_647),
.B2(n_633),
.Y(n_1384)
);

NOR2x2_ASAP7_75t_L g1385 ( 
.A(n_1365),
.B(n_763),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1282),
.B(n_648),
.Y(n_1386)
);

NOR3xp33_ASAP7_75t_L g1387 ( 
.A(n_1243),
.B(n_650),
.C(n_645),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1284),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1286),
.B(n_1193),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1323),
.A2(n_704),
.B(n_724),
.C(n_723),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1187),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1187),
.Y(n_1392)
);

OA22x2_ASAP7_75t_L g1393 ( 
.A1(n_1379),
.A2(n_655),
.B1(n_661),
.B2(n_653),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1302),
.B(n_651),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1197),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1317),
.B(n_652),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1244),
.A2(n_760),
.B1(n_788),
.B2(n_703),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1317),
.B(n_656),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1304),
.B(n_659),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1222),
.B(n_662),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1348),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1188),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1320),
.B(n_660),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_1216),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1188),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1204),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1191),
.A2(n_788),
.B1(n_760),
.B2(n_664),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1219),
.Y(n_1408)
);

NOR3xp33_ASAP7_75t_L g1409 ( 
.A(n_1198),
.B(n_671),
.C(n_670),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1186),
.B(n_663),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1377),
.Y(n_1411)
);

NAND2xp33_ASAP7_75t_L g1412 ( 
.A(n_1348),
.B(n_665),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1377),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1196),
.B(n_667),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1383),
.B(n_668),
.Y(n_1415)
);

A2O1A1Ixp33_ASAP7_75t_SL g1416 ( 
.A1(n_1338),
.A2(n_732),
.B(n_739),
.C(n_727),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1260),
.B(n_673),
.Y(n_1417)
);

NAND2xp33_ASAP7_75t_SL g1418 ( 
.A(n_1360),
.B(n_669),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1378),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1230),
.B(n_674),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1236),
.B(n_1237),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1207),
.Y(n_1422)
);

NOR3xp33_ASAP7_75t_L g1423 ( 
.A(n_1257),
.B(n_700),
.C(n_685),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1363),
.A2(n_688),
.B1(n_695),
.B2(n_678),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1368),
.A2(n_708),
.B1(n_718),
.B2(n_707),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1381),
.Y(n_1426)
);

NOR2x2_ASAP7_75t_L g1427 ( 
.A(n_1373),
.B(n_775),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1381),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1225),
.B(n_702),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1248),
.B(n_719),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1330),
.B(n_720),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1382),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1238),
.B(n_722),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1348),
.B(n_728),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1292),
.B(n_731),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1251),
.B(n_736),
.Y(n_1436)
);

BUFx12f_ASAP7_75t_L g1437 ( 
.A(n_1221),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1245),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1228),
.A2(n_744),
.B1(n_747),
.B2(n_742),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1247),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1321),
.A2(n_752),
.B(n_790),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1322),
.A2(n_791),
.B(n_761),
.Y(n_1442)
);

AND2x6_ASAP7_75t_SL g1443 ( 
.A(n_1373),
.B(n_750),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1251),
.B(n_706),
.Y(n_1444)
);

O2A1O1Ixp5_ASAP7_75t_L g1445 ( 
.A1(n_1375),
.A2(n_784),
.B(n_764),
.C(n_348),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1220),
.B(n_713),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1249),
.Y(n_1447)
);

OR2x6_ASAP7_75t_L g1448 ( 
.A(n_1350),
.B(n_934),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1297),
.B(n_716),
.Y(n_1449)
);

NOR2xp67_ASAP7_75t_L g1450 ( 
.A(n_1290),
.B(n_347),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1233),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1269),
.Y(n_1452)
);

AND2x4_ASAP7_75t_SL g1453 ( 
.A(n_1345),
.B(n_775),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1250),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1262),
.B(n_721),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1190),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1293),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1192),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1241),
.A2(n_939),
.B1(n_940),
.B2(n_937),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1214),
.A2(n_937),
.B1(n_940),
.B2(n_939),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1264),
.B(n_725),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1294),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1333),
.A2(n_939),
.B1(n_940),
.B2(n_937),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1264),
.B(n_729),
.Y(n_1464)
);

AO22x1_ASAP7_75t_L g1465 ( 
.A1(n_1273),
.A2(n_734),
.B1(n_738),
.B2(n_730),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1234),
.B(n_741),
.Y(n_1466)
);

NAND2x1p5_ASAP7_75t_L g1467 ( 
.A(n_1345),
.B(n_1339),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1266),
.B(n_746),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1327),
.B(n_749),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1312),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_1214),
.B(n_753),
.Y(n_1471)
);

OAI21xp33_ASAP7_75t_L g1472 ( 
.A1(n_1261),
.A2(n_766),
.B(n_759),
.Y(n_1472)
);

NOR2x1p5_ASAP7_75t_L g1473 ( 
.A(n_1224),
.B(n_767),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1215),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1313),
.B(n_772),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1200),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1208),
.B(n_776),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1231),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1252),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1299),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1212),
.B(n_777),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1344),
.B(n_785),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1279),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1254),
.B(n_786),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1246),
.B(n_937),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1207),
.Y(n_1486)
);

CKINVDCx20_ASAP7_75t_R g1487 ( 
.A(n_1298),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1255),
.B(n_775),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1199),
.B(n_0),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1344),
.B(n_939),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1356),
.A2(n_943),
.B1(n_944),
.B2(n_940),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1256),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1346),
.B(n_943),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1306),
.B(n_1),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1267),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1356),
.A2(n_944),
.B1(n_943),
.B2(n_942),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1194),
.B(n_943),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1349),
.B(n_944),
.Y(n_1498)
);

OAI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1369),
.A2(n_944),
.B1(n_942),
.B2(n_941),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1354),
.B(n_2),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1274),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1376),
.B(n_3),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1295),
.B(n_4),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1201),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1300),
.B(n_4),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1226),
.B(n_5),
.Y(n_1506)
);

OAI21xp33_ASAP7_75t_L g1507 ( 
.A1(n_1288),
.A2(n_5),
.B(n_6),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1226),
.B(n_349),
.Y(n_1508)
);

OAI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1370),
.A2(n_942),
.B1(n_947),
.B2(n_941),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1203),
.Y(n_1510)
);

AO22x1_ASAP7_75t_L g1511 ( 
.A1(n_1372),
.A2(n_1340),
.B1(n_1374),
.B2(n_1366),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1194),
.B(n_6),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1344),
.B(n_942),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1207),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1259),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1235),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1277),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1217),
.B(n_1227),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1227),
.B(n_1239),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1329),
.B(n_7),
.Y(n_1520)
);

NOR2x2_ASAP7_75t_L g1521 ( 
.A(n_1307),
.B(n_1309),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1217),
.B(n_947),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1319),
.B(n_8),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1350),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1239),
.B(n_8),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1206),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1235),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1209),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1314),
.A2(n_947),
.B1(n_352),
.B2(n_355),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1235),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1319),
.B(n_9),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1242),
.B(n_10),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1274),
.B(n_11),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1242),
.B(n_11),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1285),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1258),
.A2(n_947),
.B1(n_14),
.B2(n_12),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1189),
.B(n_12),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1253),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1202),
.B(n_13),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1218),
.B(n_13),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1380),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1380),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1263),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1358),
.A2(n_358),
.B1(n_359),
.B2(n_351),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1218),
.B(n_14),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1314),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1546)
);

INVx8_ASAP7_75t_L g1547 ( 
.A(n_1253),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1341),
.B(n_18),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1217),
.B(n_360),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1342),
.A2(n_364),
.B1(n_365),
.B2(n_363),
.Y(n_1550)
);

INVxp33_ASAP7_75t_L g1551 ( 
.A(n_1195),
.Y(n_1551)
);

AND2x6_ASAP7_75t_L g1552 ( 
.A(n_1281),
.B(n_366),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1372),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1253),
.B(n_367),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1210),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1314),
.A2(n_1371),
.B1(n_1367),
.B2(n_1303),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1211),
.B(n_19),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1213),
.B(n_19),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1265),
.B(n_368),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1314),
.A2(n_372),
.B1(n_374),
.B2(n_371),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1205),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1229),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1275),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1563)
);

NOR2x2_ASAP7_75t_L g1564 ( 
.A(n_1291),
.B(n_20),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1268),
.B(n_21),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1265),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1278),
.B(n_23),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1270),
.B(n_23),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1276),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1278),
.B(n_24),
.Y(n_1570)
);

OR2x6_ASAP7_75t_L g1571 ( 
.A(n_1308),
.B(n_375),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1305),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1280),
.B(n_25),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1311),
.Y(n_1574)
);

OR2x6_ASAP7_75t_L g1575 ( 
.A(n_1289),
.B(n_1246),
.Y(n_1575)
);

INVx4_ASAP7_75t_L g1576 ( 
.A(n_1289),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1296),
.Y(n_1577)
);

INVx2_ASAP7_75t_SL g1578 ( 
.A(n_1223),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1223),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1296),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1283),
.B(n_376),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1352),
.B(n_1331),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1343),
.B(n_26),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1389),
.B(n_1406),
.Y(n_1584)
);

OR2x6_ASAP7_75t_L g1585 ( 
.A(n_1547),
.B(n_1283),
.Y(n_1585)
);

NAND2xp33_ASAP7_75t_SL g1586 ( 
.A(n_1408),
.B(n_1578),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1476),
.Y(n_1587)
);

AO21x2_ASAP7_75t_L g1588 ( 
.A1(n_1442),
.A2(n_1316),
.B(n_1324),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1429),
.B(n_1388),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1395),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1400),
.B(n_1288),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1428),
.Y(n_1592)
);

NOR2x1_ASAP7_75t_R g1593 ( 
.A(n_1437),
.B(n_1281),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1417),
.B(n_1275),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1579),
.B(n_1332),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1449),
.B(n_1334),
.Y(n_1596)
);

NOR3xp33_ASAP7_75t_SL g1597 ( 
.A(n_1494),
.B(n_1359),
.C(n_1351),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1519),
.B(n_1452),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1444),
.B(n_1315),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1467),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1467),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1422),
.Y(n_1602)
);

CKINVDCx8_ASAP7_75t_R g1603 ( 
.A(n_1443),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1421),
.B(n_1337),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1422),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1432),
.Y(n_1606)
);

AOI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1446),
.A2(n_1347),
.B1(n_1287),
.B2(n_1336),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1391),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1392),
.Y(n_1609)
);

NAND2xp33_ASAP7_75t_R g1610 ( 
.A(n_1561),
.B(n_1287),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1470),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1409),
.A2(n_1325),
.B1(n_1328),
.B2(n_1326),
.Y(n_1612)
);

INVx5_ASAP7_75t_L g1613 ( 
.A(n_1575),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1402),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1477),
.B(n_1353),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1542),
.B(n_1318),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1405),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1411),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1413),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1489),
.A2(n_1240),
.B1(n_1271),
.B2(n_1364),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1422),
.Y(n_1621)
);

OR2x6_ASAP7_75t_L g1622 ( 
.A(n_1547),
.B(n_1301),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1419),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1481),
.B(n_1318),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1426),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1520),
.A2(n_1240),
.B1(n_1271),
.B2(n_1355),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1457),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1456),
.Y(n_1628)
);

CKINVDCx8_ASAP7_75t_R g1629 ( 
.A(n_1443),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1462),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1466),
.B(n_1240),
.Y(n_1631)
);

BUFx12f_ASAP7_75t_L g1632 ( 
.A(n_1473),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1468),
.B(n_1240),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1480),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1438),
.Y(n_1635)
);

BUFx4f_ASAP7_75t_L g1636 ( 
.A(n_1547),
.Y(n_1636)
);

NOR3xp33_ASAP7_75t_SL g1637 ( 
.A(n_1472),
.B(n_1271),
.C(n_1232),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1455),
.B(n_1232),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1440),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1447),
.Y(n_1640)
);

INVx5_ASAP7_75t_L g1641 ( 
.A(n_1575),
.Y(n_1641)
);

INVx5_ASAP7_75t_L g1642 ( 
.A(n_1575),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1483),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1404),
.B(n_1362),
.Y(n_1644)
);

BUFx12f_ASAP7_75t_L g1645 ( 
.A(n_1501),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1454),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1451),
.B(n_1357),
.Y(n_1647)
);

NOR3xp33_ASAP7_75t_SL g1648 ( 
.A(n_1472),
.B(n_1271),
.C(n_27),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1495),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1574),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1541),
.Y(n_1651)
);

A2O1A1Ixp33_ASAP7_75t_L g1652 ( 
.A1(n_1442),
.A2(n_1357),
.B(n_1361),
.C(n_1310),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1504),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1524),
.Y(n_1654)
);

BUFx8_ASAP7_75t_SL g1655 ( 
.A(n_1487),
.Y(n_1655)
);

INVx5_ASAP7_75t_L g1656 ( 
.A(n_1527),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1510),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1553),
.B(n_1361),
.Y(n_1658)
);

BUFx8_ASAP7_75t_L g1659 ( 
.A(n_1567),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1386),
.B(n_1335),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1448),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1526),
.Y(n_1662)
);

AO221x1_ASAP7_75t_L g1663 ( 
.A1(n_1536),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.C(n_31),
.Y(n_1663)
);

NOR3xp33_ASAP7_75t_SL g1664 ( 
.A(n_1507),
.B(n_1418),
.C(n_1523),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1521),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1528),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1569),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1555),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1394),
.B(n_29),
.Y(n_1669)
);

BUFx6f_ASAP7_75t_L g1670 ( 
.A(n_1527),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1423),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1461),
.B(n_1464),
.Y(n_1672)
);

INVx3_ASAP7_75t_SL g1673 ( 
.A(n_1385),
.Y(n_1673)
);

INVx5_ASAP7_75t_L g1674 ( 
.A(n_1527),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1399),
.A2(n_1459),
.B1(n_1556),
.B2(n_1439),
.Y(n_1675)
);

CKINVDCx14_ASAP7_75t_R g1676 ( 
.A(n_1512),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1448),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1562),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1518),
.B(n_377),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1508),
.B(n_32),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1448),
.Y(n_1681)
);

INVxp67_ASAP7_75t_L g1682 ( 
.A(n_1533),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1492),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1564),
.Y(n_1684)
);

BUFx4f_ASAP7_75t_L g1685 ( 
.A(n_1552),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1511),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1515),
.Y(n_1687)
);

NAND2xp33_ASAP7_75t_R g1688 ( 
.A(n_1582),
.B(n_378),
.Y(n_1688)
);

NOR3xp33_ASAP7_75t_SL g1689 ( 
.A(n_1507),
.B(n_35),
.C(n_36),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1517),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1566),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1458),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_1506),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1475),
.B(n_36),
.Y(n_1694)
);

NOR3xp33_ASAP7_75t_SL g1695 ( 
.A(n_1531),
.B(n_37),
.C(n_38),
.Y(n_1695)
);

INVx4_ASAP7_75t_L g1696 ( 
.A(n_1566),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1508),
.B(n_38),
.Y(n_1697)
);

BUFx8_ASAP7_75t_L g1698 ( 
.A(n_1570),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1459),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1484),
.B(n_39),
.Y(n_1700)
);

BUFx4f_ASAP7_75t_L g1701 ( 
.A(n_1571),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1486),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_R g1703 ( 
.A(n_1401),
.B(n_380),
.Y(n_1703)
);

BUFx4f_ASAP7_75t_L g1704 ( 
.A(n_1571),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1474),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1441),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1486),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1500),
.B(n_42),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1478),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1479),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1441),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1711)
);

AO22x1_ASAP7_75t_L g1712 ( 
.A1(n_1552),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1436),
.B(n_46),
.Y(n_1713)
);

NAND2xp33_ASAP7_75t_SL g1714 ( 
.A(n_1551),
.B(n_47),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1401),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1514),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1535),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1497),
.B(n_382),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1580),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1577),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1514),
.Y(n_1721)
);

INVx5_ASAP7_75t_L g1722 ( 
.A(n_1552),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1557),
.Y(n_1723)
);

BUFx4f_ASAP7_75t_L g1724 ( 
.A(n_1571),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1558),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_1453),
.Y(n_1726)
);

CKINVDCx8_ASAP7_75t_R g1727 ( 
.A(n_1552),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1576),
.Y(n_1728)
);

INVxp67_ASAP7_75t_L g1729 ( 
.A(n_1488),
.Y(n_1729)
);

BUFx3_ASAP7_75t_L g1730 ( 
.A(n_1516),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_R g1731 ( 
.A(n_1516),
.B(n_383),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1403),
.B(n_48),
.Y(n_1732)
);

AND3x1_ASAP7_75t_SL g1733 ( 
.A(n_1563),
.B(n_48),
.C(n_49),
.Y(n_1733)
);

BUFx8_ASAP7_75t_L g1734 ( 
.A(n_1583),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1565),
.Y(n_1735)
);

NOR3xp33_ASAP7_75t_SL g1736 ( 
.A(n_1469),
.B(n_49),
.C(n_50),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1530),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1530),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1407),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1439),
.B(n_51),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1430),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1538),
.Y(n_1742)
);

INVx5_ASAP7_75t_L g1743 ( 
.A(n_1538),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1568),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1573),
.Y(n_1745)
);

INVx5_ASAP7_75t_L g1746 ( 
.A(n_1543),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1485),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1537),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1525),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1393),
.Y(n_1750)
);

AND2x6_ASAP7_75t_L g1751 ( 
.A(n_1560),
.B(n_384),
.Y(n_1751)
);

INVxp67_ASAP7_75t_SL g1752 ( 
.A(n_1493),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1539),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1503),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1485),
.Y(n_1755)
);

OR2x2_ASAP7_75t_SL g1756 ( 
.A(n_1532),
.B(n_52),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1471),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1410),
.B(n_53),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1498),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1534),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1396),
.A2(n_56),
.B1(n_53),
.B2(n_55),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1505),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1548),
.Y(n_1763)
);

BUFx12f_ASAP7_75t_L g1764 ( 
.A(n_1427),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1540),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1545),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1384),
.B(n_55),
.Y(n_1767)
);

INVx5_ASAP7_75t_L g1768 ( 
.A(n_1529),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1384),
.B(n_1502),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1754),
.B(n_1465),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1608),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1768),
.A2(n_1499),
.B(n_1435),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_L g1773 ( 
.A(n_1636),
.Y(n_1773)
);

INVxp67_ASAP7_75t_L g1774 ( 
.A(n_1589),
.Y(n_1774)
);

OAI21x1_ASAP7_75t_L g1775 ( 
.A1(n_1631),
.A2(n_1445),
.B(n_1463),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1748),
.B(n_1424),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1609),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1751),
.A2(n_1387),
.B1(n_1397),
.B2(n_1536),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1767),
.B(n_1414),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1768),
.A2(n_1398),
.B(n_1509),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1664),
.B(n_1546),
.C(n_1425),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1729),
.B(n_1431),
.Y(n_1782)
);

INVx3_ASAP7_75t_L g1783 ( 
.A(n_1727),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1768),
.A2(n_1581),
.B(n_1434),
.Y(n_1784)
);

OAI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1769),
.A2(n_1420),
.B(n_1415),
.Y(n_1785)
);

OAI21x1_ASAP7_75t_L g1786 ( 
.A1(n_1633),
.A2(n_1463),
.B(n_1550),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1753),
.B(n_1390),
.Y(n_1787)
);

OAI21x1_ASAP7_75t_L g1788 ( 
.A1(n_1675),
.A2(n_1559),
.B(n_1554),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1693),
.B(n_1433),
.Y(n_1789)
);

AOI21x1_ASAP7_75t_L g1790 ( 
.A1(n_1591),
.A2(n_1490),
.B(n_1549),
.Y(n_1790)
);

OAI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1596),
.A2(n_1482),
.B(n_1412),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1614),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1723),
.B(n_1572),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1685),
.A2(n_1529),
.B(n_1560),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1613),
.B(n_1522),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1725),
.B(n_1450),
.Y(n_1796)
);

BUFx6f_ASAP7_75t_L g1797 ( 
.A(n_1636),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1630),
.Y(n_1798)
);

OAI21x1_ASAP7_75t_L g1799 ( 
.A1(n_1763),
.A2(n_1544),
.B(n_1460),
.Y(n_1799)
);

NAND2x1_ASAP7_75t_L g1800 ( 
.A(n_1600),
.B(n_1491),
.Y(n_1800)
);

O2A1O1Ixp5_ASAP7_75t_L g1801 ( 
.A1(n_1740),
.A2(n_1416),
.B(n_1513),
.C(n_1496),
.Y(n_1801)
);

OAI21x1_ASAP7_75t_L g1802 ( 
.A1(n_1763),
.A2(n_386),
.B(n_385),
.Y(n_1802)
);

OAI21x1_ASAP7_75t_L g1803 ( 
.A1(n_1624),
.A2(n_390),
.B(n_387),
.Y(n_1803)
);

OAI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1735),
.A2(n_56),
.B(n_57),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1634),
.Y(n_1805)
);

OAI21x1_ASAP7_75t_L g1806 ( 
.A1(n_1600),
.A2(n_1601),
.B(n_1747),
.Y(n_1806)
);

OA21x2_ASAP7_75t_L g1807 ( 
.A1(n_1652),
.A2(n_392),
.B(n_391),
.Y(n_1807)
);

OAI21x1_ASAP7_75t_L g1808 ( 
.A1(n_1601),
.A2(n_395),
.B(n_393),
.Y(n_1808)
);

OAI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1744),
.A2(n_58),
.B(n_59),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1685),
.A2(n_548),
.B(n_399),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1682),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_1811)
);

AOI21x1_ASAP7_75t_L g1812 ( 
.A1(n_1594),
.A2(n_400),
.B(n_396),
.Y(n_1812)
);

CKINVDCx20_ASAP7_75t_R g1813 ( 
.A(n_1655),
.Y(n_1813)
);

INVxp67_ASAP7_75t_L g1814 ( 
.A(n_1665),
.Y(n_1814)
);

OAI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1745),
.A2(n_61),
.B(n_62),
.Y(n_1815)
);

AOI21xp33_ASAP7_75t_L g1816 ( 
.A1(n_1672),
.A2(n_1713),
.B(n_1615),
.Y(n_1816)
);

INVx4_ASAP7_75t_L g1817 ( 
.A(n_1613),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1691),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1755),
.A2(n_1759),
.B(n_1612),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1590),
.Y(n_1820)
);

OAI21x1_ASAP7_75t_L g1821 ( 
.A1(n_1762),
.A2(n_404),
.B(n_403),
.Y(n_1821)
);

OAI21x1_ASAP7_75t_L g1822 ( 
.A1(n_1620),
.A2(n_406),
.B(n_405),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1765),
.B(n_62),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1722),
.A2(n_547),
.B(n_408),
.Y(n_1824)
);

OAI21x1_ASAP7_75t_SL g1825 ( 
.A1(n_1660),
.A2(n_1699),
.B(n_1708),
.Y(n_1825)
);

NAND2x1p5_ASAP7_75t_L g1826 ( 
.A(n_1613),
.B(n_407),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1751),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1635),
.Y(n_1828)
);

AO31x2_ASAP7_75t_L g1829 ( 
.A1(n_1618),
.A2(n_65),
.A3(n_63),
.B(n_64),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1766),
.B(n_66),
.Y(n_1830)
);

INVx4_ASAP7_75t_L g1831 ( 
.A(n_1641),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1669),
.A2(n_66),
.B(n_67),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1651),
.Y(n_1833)
);

AOI21x1_ASAP7_75t_L g1834 ( 
.A1(n_1638),
.A2(n_1732),
.B(n_1758),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1654),
.Y(n_1835)
);

INVx2_ASAP7_75t_SL g1836 ( 
.A(n_1643),
.Y(n_1836)
);

NAND2x1p5_ASAP7_75t_L g1837 ( 
.A(n_1641),
.B(n_409),
.Y(n_1837)
);

INVx3_ASAP7_75t_SL g1838 ( 
.A(n_1611),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1752),
.A2(n_68),
.B(n_70),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1584),
.B(n_71),
.Y(n_1840)
);

BUFx2_ASAP7_75t_L g1841 ( 
.A(n_1716),
.Y(n_1841)
);

O2A1O1Ixp5_ASAP7_75t_L g1842 ( 
.A1(n_1712),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1607),
.A2(n_1597),
.B(n_1694),
.Y(n_1843)
);

INVx1_ASAP7_75t_SL g1844 ( 
.A(n_1599),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1749),
.B(n_73),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1749),
.B(n_74),
.Y(n_1846)
);

OA21x2_ASAP7_75t_L g1847 ( 
.A1(n_1623),
.A2(n_418),
.B(n_417),
.Y(n_1847)
);

INVx2_ASAP7_75t_SL g1848 ( 
.A(n_1645),
.Y(n_1848)
);

OAI21x1_ASAP7_75t_L g1849 ( 
.A1(n_1625),
.A2(n_423),
.B(n_421),
.Y(n_1849)
);

OAI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1706),
.A2(n_427),
.B(n_425),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1711),
.A2(n_430),
.B(n_428),
.Y(n_1851)
);

OAI21x1_ASAP7_75t_L g1852 ( 
.A1(n_1628),
.A2(n_435),
.B(n_431),
.Y(n_1852)
);

NAND2x1p5_ASAP7_75t_L g1853 ( 
.A(n_1641),
.B(n_438),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_SL g1854 ( 
.A1(n_1718),
.A2(n_440),
.B(n_439),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1701),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1617),
.Y(n_1856)
);

OAI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1648),
.A2(n_77),
.B(n_79),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1642),
.B(n_441),
.Y(n_1858)
);

AO31x2_ASAP7_75t_L g1859 ( 
.A1(n_1619),
.A2(n_82),
.A3(n_80),
.B(n_81),
.Y(n_1859)
);

OAI21x1_ASAP7_75t_L g1860 ( 
.A1(n_1626),
.A2(n_444),
.B(n_443),
.Y(n_1860)
);

OAI21x1_ASAP7_75t_SL g1861 ( 
.A1(n_1604),
.A2(n_80),
.B(n_82),
.Y(n_1861)
);

BUFx2_ASAP7_75t_L g1862 ( 
.A(n_1702),
.Y(n_1862)
);

AOI221x1_ASAP7_75t_L g1863 ( 
.A1(n_1714),
.A2(n_86),
.B1(n_83),
.B2(n_84),
.C(n_87),
.Y(n_1863)
);

NOR2x1_ASAP7_75t_L g1864 ( 
.A(n_1588),
.B(n_83),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1704),
.A2(n_1724),
.B1(n_1686),
.B2(n_1749),
.Y(n_1865)
);

NOR3xp33_ASAP7_75t_L g1866 ( 
.A(n_1680),
.B(n_86),
.C(n_87),
.Y(n_1866)
);

AO31x2_ASAP7_75t_L g1867 ( 
.A1(n_1653),
.A2(n_90),
.A3(n_88),
.B(n_89),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1760),
.B(n_88),
.Y(n_1868)
);

INVxp67_ASAP7_75t_L g1869 ( 
.A(n_1719),
.Y(n_1869)
);

OAI21x1_ASAP7_75t_L g1870 ( 
.A1(n_1592),
.A2(n_448),
.B(n_447),
.Y(n_1870)
);

BUFx3_ASAP7_75t_L g1871 ( 
.A(n_1707),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1721),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1739),
.A2(n_89),
.B(n_91),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1760),
.B(n_91),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1751),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_1875)
);

INVx5_ASAP7_75t_SL g1876 ( 
.A(n_1585),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1639),
.Y(n_1877)
);

BUFx6f_ASAP7_75t_L g1878 ( 
.A(n_1656),
.Y(n_1878)
);

INVx4_ASAP7_75t_L g1879 ( 
.A(n_1642),
.Y(n_1879)
);

OAI21x1_ASAP7_75t_L g1880 ( 
.A1(n_1606),
.A2(n_451),
.B(n_450),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1656),
.Y(n_1881)
);

INVx5_ASAP7_75t_L g1882 ( 
.A(n_1585),
.Y(n_1882)
);

A2O1A1Ixp33_ASAP7_75t_L g1883 ( 
.A1(n_1689),
.A2(n_95),
.B(n_92),
.C(n_94),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1760),
.B(n_454),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1695),
.B(n_96),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1627),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1691),
.Y(n_1887)
);

AOI21x1_ASAP7_75t_L g1888 ( 
.A1(n_1712),
.A2(n_461),
.B(n_459),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_SL g1889 ( 
.A1(n_1718),
.A2(n_464),
.B(n_462),
.Y(n_1889)
);

BUFx3_ASAP7_75t_L g1890 ( 
.A(n_1730),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1646),
.B(n_96),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1650),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1738),
.Y(n_1893)
);

AOI221x1_ASAP7_75t_L g1894 ( 
.A1(n_1663),
.A2(n_101),
.B1(n_98),
.B2(n_99),
.C(n_102),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1662),
.Y(n_1895)
);

A2O1A1Ixp33_ASAP7_75t_L g1896 ( 
.A1(n_1671),
.A2(n_102),
.B(n_98),
.C(n_101),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1668),
.Y(n_1897)
);

OAI22x1_ASAP7_75t_L g1898 ( 
.A1(n_1761),
.A2(n_1750),
.B1(n_1697),
.B2(n_1673),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1642),
.A2(n_1598),
.B(n_1616),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1640),
.Y(n_1900)
);

BUFx10_ASAP7_75t_L g1901 ( 
.A(n_1587),
.Y(n_1901)
);

OAI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1700),
.A2(n_103),
.B(n_104),
.Y(n_1902)
);

BUFx2_ASAP7_75t_L g1903 ( 
.A(n_1734),
.Y(n_1903)
);

AOI21x1_ASAP7_75t_L g1904 ( 
.A1(n_1657),
.A2(n_468),
.B(n_467),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1741),
.B(n_103),
.Y(n_1905)
);

INVxp67_ASAP7_75t_L g1906 ( 
.A(n_1734),
.Y(n_1906)
);

INVx1_ASAP7_75t_SL g1907 ( 
.A(n_1742),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1720),
.A2(n_473),
.B(n_472),
.Y(n_1908)
);

OAI21x1_ASAP7_75t_L g1909 ( 
.A1(n_1666),
.A2(n_478),
.B(n_475),
.Y(n_1909)
);

BUFx6f_ASAP7_75t_L g1910 ( 
.A(n_1656),
.Y(n_1910)
);

BUFx2_ASAP7_75t_L g1911 ( 
.A(n_1737),
.Y(n_1911)
);

OAI21x1_ASAP7_75t_L g1912 ( 
.A1(n_1667),
.A2(n_483),
.B(n_482),
.Y(n_1912)
);

BUFx6f_ASAP7_75t_L g1913 ( 
.A(n_1674),
.Y(n_1913)
);

CKINVDCx20_ASAP7_75t_R g1914 ( 
.A(n_1586),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1632),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1649),
.A2(n_485),
.B(n_484),
.Y(n_1916)
);

OAI22x1_ASAP7_75t_L g1917 ( 
.A1(n_1679),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_1917)
);

BUFx4f_ASAP7_75t_SL g1918 ( 
.A(n_1764),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1757),
.B(n_105),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1679),
.A2(n_493),
.B(n_492),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1644),
.A2(n_109),
.B1(n_106),
.B2(n_107),
.Y(n_1921)
);

AOI21xp33_ASAP7_75t_L g1922 ( 
.A1(n_1688),
.A2(n_109),
.B(n_110),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1681),
.A2(n_499),
.B(n_496),
.Y(n_1923)
);

OAI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1751),
.A2(n_111),
.B(n_112),
.Y(n_1924)
);

OAI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1647),
.A2(n_111),
.B(n_112),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1678),
.Y(n_1926)
);

AOI21x1_ASAP7_75t_L g1927 ( 
.A1(n_1661),
.A2(n_503),
.B(n_501),
.Y(n_1927)
);

AOI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1677),
.A2(n_507),
.B(n_504),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1794),
.A2(n_1663),
.B(n_1674),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1844),
.B(n_1756),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1844),
.B(n_1683),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1778),
.A2(n_1736),
.B1(n_1676),
.B2(n_1637),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1771),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1779),
.B(n_1692),
.Y(n_1934)
);

CKINVDCx20_ASAP7_75t_R g1935 ( 
.A(n_1813),
.Y(n_1935)
);

OR2x6_ASAP7_75t_L g1936 ( 
.A(n_1854),
.B(n_1681),
.Y(n_1936)
);

BUFx4_ASAP7_75t_SL g1937 ( 
.A(n_1914),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1789),
.B(n_1705),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1816),
.B(n_1687),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1774),
.B(n_1690),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1787),
.B(n_1710),
.Y(n_1941)
);

BUFx8_ASAP7_75t_L g1942 ( 
.A(n_1903),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1771),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1777),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1776),
.B(n_1717),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1885),
.B(n_1709),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1772),
.A2(n_1746),
.B(n_1622),
.Y(n_1947)
);

A2O1A1Ixp33_ASAP7_75t_L g1948 ( 
.A1(n_1843),
.A2(n_1595),
.B(n_1726),
.C(n_1658),
.Y(n_1948)
);

AO21x2_ASAP7_75t_L g1949 ( 
.A1(n_1780),
.A2(n_1703),
.B(n_1731),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1882),
.B(n_1746),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1798),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1845),
.B(n_1684),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1833),
.B(n_1715),
.Y(n_1953)
);

BUFx3_ASAP7_75t_L g1954 ( 
.A(n_1820),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1805),
.Y(n_1955)
);

NAND2x1p5_ASAP7_75t_L g1956 ( 
.A(n_1882),
.B(n_1743),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1828),
.Y(n_1957)
);

BUFx2_ASAP7_75t_L g1958 ( 
.A(n_1841),
.Y(n_1958)
);

BUFx2_ASAP7_75t_L g1959 ( 
.A(n_1862),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1777),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1846),
.B(n_1715),
.Y(n_1961)
);

INVx5_ASAP7_75t_L g1962 ( 
.A(n_1878),
.Y(n_1962)
);

BUFx6f_ASAP7_75t_L g1963 ( 
.A(n_1878),
.Y(n_1963)
);

AOI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1785),
.A2(n_1746),
.B(n_1622),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1878),
.Y(n_1965)
);

A2O1A1Ixp33_ASAP7_75t_SL g1966 ( 
.A1(n_1832),
.A2(n_1733),
.B(n_1610),
.C(n_1629),
.Y(n_1966)
);

BUFx2_ASAP7_75t_L g1967 ( 
.A(n_1872),
.Y(n_1967)
);

AO21x2_ASAP7_75t_L g1968 ( 
.A1(n_1825),
.A2(n_1658),
.B(n_1595),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1850),
.A2(n_1743),
.B(n_1593),
.Y(n_1969)
);

INVx2_ASAP7_75t_SL g1970 ( 
.A(n_1871),
.Y(n_1970)
);

INVx1_ASAP7_75t_SL g1971 ( 
.A(n_1835),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1924),
.A2(n_1698),
.B1(n_1659),
.B2(n_1737),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1874),
.B(n_1737),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1781),
.A2(n_1698),
.B1(n_1659),
.B2(n_1696),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1877),
.Y(n_1975)
);

INVx4_ASAP7_75t_L g1976 ( 
.A(n_1881),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1781),
.A2(n_1603),
.B1(n_1743),
.B2(n_1696),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1901),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1882),
.B(n_1691),
.Y(n_1979)
);

BUFx2_ASAP7_75t_L g1980 ( 
.A(n_1911),
.Y(n_1980)
);

AOI22xp33_ASAP7_75t_L g1981 ( 
.A1(n_1873),
.A2(n_1728),
.B1(n_1605),
.B2(n_1621),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1881),
.Y(n_1982)
);

BUFx6f_ASAP7_75t_SL g1983 ( 
.A(n_1901),
.Y(n_1983)
);

INVx8_ASAP7_75t_L g1984 ( 
.A(n_1881),
.Y(n_1984)
);

INVx2_ASAP7_75t_SL g1985 ( 
.A(n_1890),
.Y(n_1985)
);

AOI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1850),
.A2(n_1728),
.B(n_1605),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_1910),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1793),
.B(n_1892),
.Y(n_1988)
);

AOI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1898),
.A2(n_1728),
.B1(n_1605),
.B2(n_1621),
.Y(n_1989)
);

INVx3_ASAP7_75t_L g1990 ( 
.A(n_1910),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1827),
.B(n_1602),
.Y(n_1991)
);

CKINVDCx20_ASAP7_75t_R g1992 ( 
.A(n_1838),
.Y(n_1992)
);

INVxp67_ASAP7_75t_SL g1993 ( 
.A(n_1893),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1895),
.B(n_1602),
.Y(n_1994)
);

OAI22x1_ASAP7_75t_L g1995 ( 
.A1(n_1827),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_1995)
);

BUFx12f_ASAP7_75t_L g1996 ( 
.A(n_1915),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1875),
.B(n_1602),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1897),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1907),
.B(n_1621),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1907),
.B(n_1670),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1792),
.Y(n_2001)
);

INVx3_ASAP7_75t_L g2002 ( 
.A(n_1910),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1902),
.B(n_1670),
.Y(n_2003)
);

BUFx6f_ASAP7_75t_L g2004 ( 
.A(n_1913),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1869),
.B(n_1670),
.Y(n_2005)
);

A2O1A1Ixp33_ASAP7_75t_L g2006 ( 
.A1(n_1851),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_2006)
);

OAI221xp5_ASAP7_75t_L g2007 ( 
.A1(n_1875),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.C(n_119),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1770),
.B(n_508),
.Y(n_2008)
);

BUFx6f_ASAP7_75t_L g2009 ( 
.A(n_1913),
.Y(n_2009)
);

INVx4_ASAP7_75t_L g2010 ( 
.A(n_1913),
.Y(n_2010)
);

OAI21x1_ASAP7_75t_SL g2011 ( 
.A1(n_1790),
.A2(n_1834),
.B(n_1784),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1856),
.B(n_116),
.Y(n_2012)
);

INVx6_ASAP7_75t_L g2013 ( 
.A(n_1773),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1926),
.B(n_1856),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1866),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_2015)
);

BUFx2_ASAP7_75t_L g2016 ( 
.A(n_1814),
.Y(n_2016)
);

INVxp67_ASAP7_75t_L g2017 ( 
.A(n_1782),
.Y(n_2017)
);

BUFx12f_ASAP7_75t_L g2018 ( 
.A(n_1773),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1796),
.B(n_513),
.Y(n_2019)
);

BUFx3_ASAP7_75t_L g2020 ( 
.A(n_1836),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1886),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1783),
.B(n_514),
.Y(n_2022)
);

INVx5_ASAP7_75t_L g2023 ( 
.A(n_1817),
.Y(n_2023)
);

O2A1O1Ixp33_ASAP7_75t_L g2024 ( 
.A1(n_1896),
.A2(n_122),
.B(n_120),
.C(n_121),
.Y(n_2024)
);

CKINVDCx16_ASAP7_75t_R g2025 ( 
.A(n_1865),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1792),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_L g2027 ( 
.A(n_1773),
.Y(n_2027)
);

BUFx6f_ASAP7_75t_L g2028 ( 
.A(n_1797),
.Y(n_2028)
);

OAI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_1883),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_2029)
);

BUFx4f_ASAP7_75t_L g2030 ( 
.A(n_1797),
.Y(n_2030)
);

BUFx3_ASAP7_75t_L g2031 ( 
.A(n_1848),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1851),
.A2(n_518),
.B(n_517),
.Y(n_2032)
);

INVx1_ASAP7_75t_SL g2033 ( 
.A(n_1818),
.Y(n_2033)
);

BUFx6f_ASAP7_75t_L g2034 ( 
.A(n_1797),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_SL g2035 ( 
.A(n_1831),
.B(n_519),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1886),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1900),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1884),
.B(n_520),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1840),
.B(n_521),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1900),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1831),
.B(n_524),
.Y(n_2041)
);

BUFx3_ASAP7_75t_L g2042 ( 
.A(n_1887),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1879),
.B(n_525),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1879),
.B(n_527),
.Y(n_2044)
);

OAI21x1_ASAP7_75t_L g2045 ( 
.A1(n_2011),
.A2(n_1775),
.B(n_1786),
.Y(n_2045)
);

OAI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_2032),
.A2(n_1839),
.B(n_1925),
.Y(n_2046)
);

O2A1O1Ixp33_ASAP7_75t_L g2047 ( 
.A1(n_2006),
.A2(n_1855),
.B(n_1857),
.C(n_1922),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1944),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1944),
.Y(n_2049)
);

BUFx6f_ASAP7_75t_L g2050 ( 
.A(n_1954),
.Y(n_2050)
);

OAI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_2024),
.A2(n_1929),
.B(n_1809),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_2017),
.B(n_1919),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2037),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2037),
.Y(n_2054)
);

AOI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_2007),
.A2(n_1917),
.B1(n_1815),
.B2(n_1804),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_L g2056 ( 
.A(n_2025),
.B(n_1905),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_1993),
.B(n_1864),
.Y(n_2057)
);

OAI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_2015),
.A2(n_1863),
.B1(n_1894),
.B2(n_1921),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1973),
.B(n_1934),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2021),
.Y(n_2060)
);

BUFx2_ASAP7_75t_L g2061 ( 
.A(n_1959),
.Y(n_2061)
);

AO21x2_ASAP7_75t_L g2062 ( 
.A1(n_2011),
.A2(n_1888),
.B(n_1812),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1939),
.B(n_1830),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1933),
.Y(n_2064)
);

OAI21x1_ASAP7_75t_L g2065 ( 
.A1(n_1947),
.A2(n_1788),
.B(n_1864),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1943),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1960),
.Y(n_2067)
);

INVx1_ASAP7_75t_SL g2068 ( 
.A(n_1958),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2001),
.Y(n_2069)
);

OAI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_2029),
.A2(n_1811),
.B1(n_1823),
.B2(n_1891),
.Y(n_2070)
);

OAI21x1_ASAP7_75t_L g2071 ( 
.A1(n_1964),
.A2(n_1802),
.B(n_1927),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1988),
.B(n_1867),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2026),
.Y(n_2073)
);

AO21x2_ASAP7_75t_L g2074 ( 
.A1(n_1969),
.A2(n_1861),
.B(n_1928),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2036),
.B(n_1829),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1945),
.B(n_1867),
.Y(n_2076)
);

OAI21x1_ASAP7_75t_L g2077 ( 
.A1(n_1986),
.A2(n_1904),
.B(n_1803),
.Y(n_2077)
);

AO22x2_ASAP7_75t_L g2078 ( 
.A1(n_1932),
.A2(n_1997),
.B1(n_1991),
.B2(n_1977),
.Y(n_2078)
);

INVx5_ASAP7_75t_L g2079 ( 
.A(n_1936),
.Y(n_2079)
);

O2A1O1Ixp33_ASAP7_75t_SL g2080 ( 
.A1(n_1966),
.A2(n_1868),
.B(n_1906),
.C(n_1791),
.Y(n_2080)
);

CKINVDCx20_ASAP7_75t_R g2081 ( 
.A(n_1935),
.Y(n_2081)
);

OA21x2_ASAP7_75t_L g2082 ( 
.A1(n_1948),
.A2(n_1842),
.B(n_1819),
.Y(n_2082)
);

OAI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_1972),
.A2(n_1920),
.B1(n_1826),
.B2(n_1853),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2040),
.Y(n_2084)
);

OAI21x1_ASAP7_75t_L g2085 ( 
.A1(n_2014),
.A2(n_1849),
.B(n_1909),
.Y(n_2085)
);

OAI21xp5_ASAP7_75t_L g2086 ( 
.A1(n_1981),
.A2(n_1916),
.B(n_1801),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1951),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1955),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1957),
.Y(n_2089)
);

AOI21x1_ASAP7_75t_L g2090 ( 
.A1(n_2003),
.A2(n_1899),
.B(n_1847),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_L g2091 ( 
.A(n_1971),
.B(n_1783),
.Y(n_2091)
);

INVx3_ASAP7_75t_L g2092 ( 
.A(n_1950),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1975),
.Y(n_2093)
);

OAI21x1_ASAP7_75t_L g2094 ( 
.A1(n_1941),
.A2(n_1912),
.B(n_1852),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1961),
.B(n_1829),
.Y(n_2095)
);

INVx5_ASAP7_75t_L g2096 ( 
.A(n_1936),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_1967),
.B(n_1806),
.Y(n_2097)
);

OA21x2_ASAP7_75t_L g2098 ( 
.A1(n_1931),
.A2(n_1908),
.B(n_1821),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1998),
.B(n_1859),
.Y(n_2099)
);

AO21x2_ASAP7_75t_L g2100 ( 
.A1(n_1968),
.A2(n_1880),
.B(n_1870),
.Y(n_2100)
);

BUFx10_ASAP7_75t_L g2101 ( 
.A(n_1983),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1940),
.Y(n_2102)
);

CKINVDCx20_ASAP7_75t_R g2103 ( 
.A(n_1992),
.Y(n_2103)
);

INVxp67_ASAP7_75t_L g2104 ( 
.A(n_1938),
.Y(n_2104)
);

OA21x2_ASAP7_75t_L g2105 ( 
.A1(n_1989),
.A2(n_1799),
.B(n_1822),
.Y(n_2105)
);

INVxp67_ASAP7_75t_SL g2106 ( 
.A(n_1953),
.Y(n_2106)
);

OAI21x1_ASAP7_75t_L g2107 ( 
.A1(n_1956),
.A2(n_1808),
.B(n_1807),
.Y(n_2107)
);

OAI21xp33_ASAP7_75t_SL g2108 ( 
.A1(n_2019),
.A2(n_1860),
.B(n_1889),
.Y(n_2108)
);

AOI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_1995),
.A2(n_1858),
.B1(n_1810),
.B2(n_1923),
.Y(n_2109)
);

INVx3_ASAP7_75t_SL g2110 ( 
.A(n_1978),
.Y(n_2110)
);

OAI21x1_ASAP7_75t_L g2111 ( 
.A1(n_1946),
.A2(n_1807),
.B(n_1824),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1994),
.Y(n_2112)
);

CKINVDCx11_ASAP7_75t_R g2113 ( 
.A(n_1996),
.Y(n_2113)
);

OAI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_1974),
.A2(n_1800),
.B(n_1837),
.Y(n_2114)
);

INVx6_ASAP7_75t_L g2115 ( 
.A(n_1942),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2106),
.B(n_1930),
.Y(n_2116)
);

AOI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_2046),
.A2(n_1949),
.B1(n_2008),
.B2(n_1952),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2048),
.Y(n_2118)
);

NAND3xp33_ASAP7_75t_L g2119 ( 
.A(n_2051),
.B(n_2012),
.C(n_2035),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2102),
.B(n_2016),
.Y(n_2120)
);

OAI21x1_ASAP7_75t_L g2121 ( 
.A1(n_2065),
.A2(n_1847),
.B(n_1982),
.Y(n_2121)
);

AOI221xp5_ASAP7_75t_L g2122 ( 
.A1(n_2058),
.A2(n_2039),
.B1(n_2005),
.B2(n_2022),
.C(n_1980),
.Y(n_2122)
);

INVxp67_ASAP7_75t_L g2123 ( 
.A(n_2061),
.Y(n_2123)
);

AOI21xp5_ASAP7_75t_L g2124 ( 
.A1(n_2046),
.A2(n_1950),
.B(n_1858),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2060),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2095),
.B(n_1859),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2049),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2068),
.B(n_2059),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2084),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_2081),
.Y(n_2130)
);

CKINVDCx8_ASAP7_75t_R g2131 ( 
.A(n_2050),
.Y(n_2131)
);

A2O1A1Ixp33_ASAP7_75t_L g2132 ( 
.A1(n_2047),
.A2(n_2038),
.B(n_2043),
.C(n_2041),
.Y(n_2132)
);

INVx4_ASAP7_75t_L g2133 ( 
.A(n_2079),
.Y(n_2133)
);

INVx3_ASAP7_75t_L g2134 ( 
.A(n_2092),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_2097),
.B(n_1999),
.Y(n_2135)
);

HB1xp67_ASAP7_75t_L g2136 ( 
.A(n_2057),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2063),
.B(n_1999),
.Y(n_2137)
);

INVx4_ASAP7_75t_L g2138 ( 
.A(n_2079),
.Y(n_2138)
);

BUFx12f_ASAP7_75t_L g2139 ( 
.A(n_2113),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2053),
.Y(n_2140)
);

BUFx12f_ASAP7_75t_L g2141 ( 
.A(n_2101),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2112),
.B(n_2000),
.Y(n_2142)
);

CKINVDCx16_ASAP7_75t_R g2143 ( 
.A(n_2103),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2068),
.B(n_1970),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2075),
.B(n_2033),
.Y(n_2145)
);

OAI22xp33_ASAP7_75t_L g2146 ( 
.A1(n_2055),
.A2(n_2023),
.B1(n_1962),
.B2(n_2020),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_2056),
.B(n_2031),
.Y(n_2147)
);

OAI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_2055),
.A2(n_1876),
.B1(n_1985),
.B2(n_2013),
.Y(n_2148)
);

NOR3xp33_ASAP7_75t_L g2149 ( 
.A(n_2051),
.B(n_2010),
.C(n_1976),
.Y(n_2149)
);

OAI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_2109),
.A2(n_2070),
.B1(n_2096),
.B2(n_2079),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_2092),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2054),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2064),
.Y(n_2153)
);

AOI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_2070),
.A2(n_2078),
.B1(n_2052),
.B2(n_2083),
.Y(n_2154)
);

A2O1A1Ixp33_ASAP7_75t_L g2155 ( 
.A1(n_2108),
.A2(n_2043),
.B(n_2044),
.C(n_2041),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_2075),
.B(n_2000),
.Y(n_2156)
);

CKINVDCx11_ASAP7_75t_R g2157 ( 
.A(n_2110),
.Y(n_2157)
);

INVx1_ASAP7_75t_SL g2158 ( 
.A(n_2050),
.Y(n_2158)
);

INVx1_ASAP7_75t_SL g2159 ( 
.A(n_2050),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_2097),
.B(n_2042),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2066),
.Y(n_2161)
);

O2A1O1Ixp33_ASAP7_75t_L g2162 ( 
.A1(n_2080),
.A2(n_1795),
.B(n_1990),
.C(n_1982),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_2078),
.A2(n_2044),
.B1(n_1795),
.B2(n_2018),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_2057),
.B(n_2023),
.Y(n_2164)
);

BUFx12f_ASAP7_75t_L g2165 ( 
.A(n_2139),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2118),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2127),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2140),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2152),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2153),
.Y(n_2170)
);

BUFx2_ASAP7_75t_L g2171 ( 
.A(n_2133),
.Y(n_2171)
);

INVx3_ASAP7_75t_L g2172 ( 
.A(n_2134),
.Y(n_2172)
);

OAI21x1_ASAP7_75t_L g2173 ( 
.A1(n_2121),
.A2(n_2045),
.B(n_2071),
.Y(n_2173)
);

OA21x2_ASAP7_75t_L g2174 ( 
.A1(n_2154),
.A2(n_2077),
.B(n_2111),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2161),
.Y(n_2175)
);

BUFx2_ASAP7_75t_SL g2176 ( 
.A(n_2133),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2129),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2125),
.B(n_2072),
.Y(n_2178)
);

OA21x2_ASAP7_75t_L g2179 ( 
.A1(n_2154),
.A2(n_2076),
.B(n_2085),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2136),
.B(n_2067),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2145),
.Y(n_2181)
);

HB1xp67_ASAP7_75t_L g2182 ( 
.A(n_2156),
.Y(n_2182)
);

BUFx3_ASAP7_75t_L g2183 ( 
.A(n_2138),
.Y(n_2183)
);

OA21x2_ASAP7_75t_L g2184 ( 
.A1(n_2124),
.A2(n_2099),
.B(n_2094),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2126),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2116),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2120),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2134),
.Y(n_2188)
);

AO21x2_ASAP7_75t_L g2189 ( 
.A1(n_2146),
.A2(n_2099),
.B(n_2062),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2151),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2151),
.Y(n_2191)
);

INVx2_ASAP7_75t_SL g2192 ( 
.A(n_2160),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2142),
.Y(n_2193)
);

OAI21x1_ASAP7_75t_L g2194 ( 
.A1(n_2173),
.A2(n_2090),
.B(n_2163),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_2183),
.B(n_2138),
.Y(n_2195)
);

NOR2x1_ASAP7_75t_SL g2196 ( 
.A(n_2176),
.B(n_2096),
.Y(n_2196)
);

OAI22xp33_ASAP7_75t_L g2197 ( 
.A1(n_2192),
.A2(n_2119),
.B1(n_2163),
.B2(n_2150),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2166),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2192),
.B(n_2128),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2192),
.B(n_2123),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_2165),
.B(n_2141),
.Y(n_2201)
);

OAI21x1_ASAP7_75t_L g2202 ( 
.A1(n_2173),
.A2(n_2107),
.B(n_2073),
.Y(n_2202)
);

OAI221xp5_ASAP7_75t_SL g2203 ( 
.A1(n_2187),
.A2(n_2122),
.B1(n_2117),
.B2(n_2119),
.C(n_2132),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2186),
.B(n_2137),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2195),
.B(n_2185),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2198),
.Y(n_2206)
);

BUFx2_ASAP7_75t_L g2207 ( 
.A(n_2195),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2198),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2200),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2195),
.B(n_2185),
.Y(n_2210)
);

NOR2xp33_ASAP7_75t_L g2211 ( 
.A(n_2201),
.B(n_2165),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2200),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2205),
.Y(n_2213)
);

OAI221xp5_ASAP7_75t_L g2214 ( 
.A1(n_2207),
.A2(n_2203),
.B1(n_2148),
.B2(n_2187),
.C(n_2131),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2206),
.Y(n_2215)
);

HB1xp67_ASAP7_75t_L g2216 ( 
.A(n_2209),
.Y(n_2216)
);

OAI321xp33_ASAP7_75t_L g2217 ( 
.A1(n_2212),
.A2(n_2197),
.A3(n_2171),
.B1(n_2114),
.B2(n_2086),
.C(n_2204),
.Y(n_2217)
);

OAI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_2211),
.A2(n_2155),
.B1(n_2096),
.B2(n_2195),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2208),
.Y(n_2219)
);

AO21x1_ASAP7_75t_SL g2220 ( 
.A1(n_2211),
.A2(n_2196),
.B(n_2114),
.Y(n_2220)
);

NOR2x1_ASAP7_75t_L g2221 ( 
.A(n_2205),
.B(n_2171),
.Y(n_2221)
);

INVx3_ASAP7_75t_L g2222 ( 
.A(n_2210),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2222),
.B(n_2210),
.Y(n_2223)
);

NAND3xp33_ASAP7_75t_L g2224 ( 
.A(n_2214),
.B(n_2149),
.C(n_2179),
.Y(n_2224)
);

AOI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_2218),
.A2(n_2179),
.B1(n_2189),
.B2(n_2174),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2216),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2222),
.B(n_2199),
.Y(n_2227)
);

AOI221xp5_ASAP7_75t_L g2228 ( 
.A1(n_2217),
.A2(n_2186),
.B1(n_2178),
.B2(n_2193),
.C(n_2181),
.Y(n_2228)
);

NAND4xp25_ASAP7_75t_L g2229 ( 
.A(n_2221),
.B(n_2091),
.C(n_2147),
.D(n_2162),
.Y(n_2229)
);

NAND3xp33_ASAP7_75t_L g2230 ( 
.A(n_2216),
.B(n_2179),
.C(n_2174),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_L g2231 ( 
.A(n_2213),
.B(n_2165),
.Y(n_2231)
);

AOI22xp33_ASAP7_75t_L g2232 ( 
.A1(n_2220),
.A2(n_2179),
.B1(n_2174),
.B2(n_2189),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2213),
.B(n_2199),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2226),
.B(n_2215),
.Y(n_2234)
);

HB1xp67_ASAP7_75t_L g2235 ( 
.A(n_2223),
.Y(n_2235)
);

HB1xp67_ASAP7_75t_L g2236 ( 
.A(n_2227),
.Y(n_2236)
);

AOI22xp33_ASAP7_75t_L g2237 ( 
.A1(n_2224),
.A2(n_2219),
.B1(n_2179),
.B2(n_2174),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2231),
.B(n_2101),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_2228),
.B(n_2143),
.Y(n_2239)
);

OAI221xp5_ASAP7_75t_L g2240 ( 
.A1(n_2225),
.A2(n_2171),
.B1(n_2183),
.B2(n_2176),
.C(n_2115),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_2233),
.B(n_2196),
.Y(n_2241)
);

HB1xp67_ASAP7_75t_L g2242 ( 
.A(n_2230),
.Y(n_2242)
);

OAI211xp5_ASAP7_75t_SL g2243 ( 
.A1(n_2239),
.A2(n_2232),
.B(n_2157),
.C(n_2229),
.Y(n_2243)
);

NAND2x1_ASAP7_75t_L g2244 ( 
.A(n_2241),
.B(n_2115),
.Y(n_2244)
);

INVx2_ASAP7_75t_SL g2245 ( 
.A(n_2235),
.Y(n_2245)
);

INVx1_ASAP7_75t_SL g2246 ( 
.A(n_2236),
.Y(n_2246)
);

NOR2xp33_ASAP7_75t_R g2247 ( 
.A(n_2245),
.B(n_1918),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2246),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2244),
.B(n_2238),
.Y(n_2249)
);

OAI21xp5_ASAP7_75t_SL g2250 ( 
.A1(n_2243),
.A2(n_2237),
.B(n_2242),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2248),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2249),
.B(n_2234),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_2250),
.B(n_2240),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_2247),
.B(n_2130),
.Y(n_2254)
);

NAND4xp75_ASAP7_75t_L g2255 ( 
.A(n_2248),
.B(n_2242),
.C(n_1942),
.D(n_2174),
.Y(n_2255)
);

OR2x2_ASAP7_75t_L g2256 ( 
.A(n_2248),
.B(n_2182),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2252),
.B(n_2144),
.Y(n_2257)
);

OAI21xp5_ASAP7_75t_SL g2258 ( 
.A1(n_2253),
.A2(n_2251),
.B(n_2256),
.Y(n_2258)
);

NAND3xp33_ASAP7_75t_SL g2259 ( 
.A(n_2254),
.B(n_2255),
.C(n_2159),
.Y(n_2259)
);

O2A1O1Ixp33_ASAP7_75t_L g2260 ( 
.A1(n_2253),
.A2(n_2183),
.B(n_2083),
.C(n_2086),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2256),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2256),
.Y(n_2262)
);

OAI221xp5_ASAP7_75t_L g2263 ( 
.A1(n_2253),
.A2(n_2183),
.B1(n_2176),
.B2(n_2158),
.C(n_2030),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2256),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_2252),
.B(n_1962),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_L g2266 ( 
.A(n_2254),
.B(n_2193),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2257),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2261),
.B(n_2262),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2264),
.Y(n_2269)
);

AOI221x1_ASAP7_75t_L g2270 ( 
.A1(n_2259),
.A2(n_2034),
.B1(n_2028),
.B2(n_2027),
.C(n_2188),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2258),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2266),
.Y(n_2272)
);

OR2x2_ASAP7_75t_L g2273 ( 
.A(n_2265),
.B(n_2182),
.Y(n_2273)
);

INVxp67_ASAP7_75t_SL g2274 ( 
.A(n_2263),
.Y(n_2274)
);

OR2x2_ASAP7_75t_L g2275 ( 
.A(n_2260),
.B(n_2181),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2261),
.B(n_2185),
.Y(n_2276)
);

INVx2_ASAP7_75t_SL g2277 ( 
.A(n_2261),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2257),
.Y(n_2278)
);

INVxp33_ASAP7_75t_L g2279 ( 
.A(n_2258),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2268),
.Y(n_2280)
);

INVx2_ASAP7_75t_SL g2281 ( 
.A(n_2277),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2268),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2269),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2271),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2279),
.B(n_2180),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2275),
.Y(n_2286)
);

NOR2x1_ASAP7_75t_L g2287 ( 
.A(n_2272),
.B(n_2010),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2276),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2273),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2267),
.Y(n_2290)
);

INVx2_ASAP7_75t_SL g2291 ( 
.A(n_2278),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2274),
.Y(n_2292)
);

OA21x2_ASAP7_75t_L g2293 ( 
.A1(n_2270),
.A2(n_2194),
.B(n_2202),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2277),
.B(n_2170),
.Y(n_2294)
);

NOR3xp33_ASAP7_75t_L g2295 ( 
.A(n_2292),
.B(n_1937),
.C(n_1887),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2281),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2288),
.Y(n_2297)
);

NOR3x1_ASAP7_75t_L g2298 ( 
.A(n_2291),
.B(n_2194),
.C(n_2190),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_2289),
.B(n_2013),
.Y(n_2299)
);

AOI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_2284),
.A2(n_2028),
.B1(n_2034),
.B2(n_2027),
.Y(n_2300)
);

AOI211xp5_ASAP7_75t_SL g2301 ( 
.A1(n_2283),
.A2(n_1990),
.B(n_2002),
.C(n_1979),
.Y(n_2301)
);

AOI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_2285),
.A2(n_2028),
.B1(n_2034),
.B2(n_2027),
.Y(n_2302)
);

NOR2x1_ASAP7_75t_L g2303 ( 
.A(n_2280),
.B(n_2282),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2280),
.B(n_2170),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2286),
.B(n_123),
.Y(n_2305)
);

A2O1A1Ixp33_ASAP7_75t_L g2306 ( 
.A1(n_2287),
.A2(n_1984),
.B(n_2172),
.C(n_2108),
.Y(n_2306)
);

NOR2xp67_ASAP7_75t_L g2307 ( 
.A(n_2290),
.B(n_124),
.Y(n_2307)
);

INVxp67_ASAP7_75t_L g2308 ( 
.A(n_2294),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2307),
.Y(n_2309)
);

NOR3x1_ASAP7_75t_L g2310 ( 
.A(n_2296),
.B(n_2293),
.C(n_126),
.Y(n_2310)
);

OR2x2_ASAP7_75t_L g2311 ( 
.A(n_2297),
.B(n_2293),
.Y(n_2311)
);

A2O1A1Ixp33_ASAP7_75t_L g2312 ( 
.A1(n_2305),
.A2(n_1984),
.B(n_2172),
.C(n_2202),
.Y(n_2312)
);

NOR3xp33_ASAP7_75t_L g2313 ( 
.A(n_2303),
.B(n_2002),
.C(n_1979),
.Y(n_2313)
);

NAND3xp33_ASAP7_75t_L g2314 ( 
.A(n_2299),
.B(n_1962),
.C(n_1963),
.Y(n_2314)
);

NOR2x1_ASAP7_75t_L g2315 ( 
.A(n_2304),
.B(n_126),
.Y(n_2315)
);

NOR2x1p5_ASAP7_75t_L g2316 ( 
.A(n_2295),
.B(n_1963),
.Y(n_2316)
);

AOI322xp5_ASAP7_75t_L g2317 ( 
.A1(n_2308),
.A2(n_2191),
.A3(n_2190),
.B1(n_2188),
.B2(n_2180),
.C1(n_2172),
.C2(n_2164),
.Y(n_2317)
);

INVxp67_ASAP7_75t_L g2318 ( 
.A(n_2300),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2298),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2302),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_2306),
.B(n_2301),
.Y(n_2321)
);

NOR2x1_ASAP7_75t_L g2322 ( 
.A(n_2307),
.B(n_127),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2307),
.B(n_2167),
.Y(n_2323)
);

AOI22xp5_ASAP7_75t_L g2324 ( 
.A1(n_2296),
.A2(n_1876),
.B1(n_2172),
.B2(n_2191),
.Y(n_2324)
);

CKINVDCx16_ASAP7_75t_R g2325 ( 
.A(n_2296),
.Y(n_2325)
);

OR2x2_ASAP7_75t_L g2326 ( 
.A(n_2296),
.B(n_2189),
.Y(n_2326)
);

AOI21xp33_ASAP7_75t_L g2327 ( 
.A1(n_2303),
.A2(n_128),
.B(n_129),
.Y(n_2327)
);

AOI221xp5_ASAP7_75t_L g2328 ( 
.A1(n_2295),
.A2(n_2172),
.B1(n_2168),
.B2(n_2167),
.C(n_131),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2307),
.B(n_2168),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2307),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2322),
.Y(n_2331)
);

AOI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_2325),
.A2(n_2316),
.B1(n_2313),
.B2(n_2319),
.Y(n_2332)
);

AOI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_2314),
.A2(n_2189),
.B1(n_1965),
.B2(n_1987),
.Y(n_2333)
);

AO22x2_ASAP7_75t_L g2334 ( 
.A1(n_2311),
.A2(n_2169),
.B1(n_2166),
.B2(n_131),
.Y(n_2334)
);

INVxp67_ASAP7_75t_SL g2335 ( 
.A(n_2310),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2315),
.Y(n_2336)
);

NOR2x1_ASAP7_75t_L g2337 ( 
.A(n_2309),
.B(n_129),
.Y(n_2337)
);

NOR2x1p5_ASAP7_75t_L g2338 ( 
.A(n_2330),
.B(n_1963),
.Y(n_2338)
);

AOI22xp5_ASAP7_75t_L g2339 ( 
.A1(n_2321),
.A2(n_2189),
.B1(n_1987),
.B2(n_2004),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2323),
.Y(n_2340)
);

AOI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2328),
.A2(n_1987),
.B1(n_2004),
.B2(n_1965),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2329),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2327),
.B(n_130),
.Y(n_2343)
);

NOR2x1_ASAP7_75t_L g2344 ( 
.A(n_2320),
.B(n_130),
.Y(n_2344)
);

OAI22xp33_ASAP7_75t_L g2345 ( 
.A1(n_2324),
.A2(n_2004),
.B1(n_2009),
.B2(n_1965),
.Y(n_2345)
);

NOR2x1_ASAP7_75t_L g2346 ( 
.A(n_2326),
.B(n_132),
.Y(n_2346)
);

AOI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_2318),
.A2(n_2009),
.B1(n_2180),
.B2(n_2164),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2312),
.Y(n_2348)
);

AO22x1_ASAP7_75t_L g2349 ( 
.A1(n_2317),
.A2(n_2009),
.B1(n_2023),
.B2(n_135),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2322),
.Y(n_2350)
);

AOI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_2325),
.A2(n_2178),
.B1(n_2160),
.B2(n_2074),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2322),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2322),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2322),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2322),
.Y(n_2355)
);

AO22x2_ASAP7_75t_L g2356 ( 
.A1(n_2319),
.A2(n_2169),
.B1(n_2166),
.B2(n_135),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_2325),
.B(n_2169),
.Y(n_2357)
);

AOI221xp5_ASAP7_75t_L g2358 ( 
.A1(n_2327),
.A2(n_136),
.B1(n_133),
.B2(n_134),
.C(n_137),
.Y(n_2358)
);

AOI221xp5_ASAP7_75t_L g2359 ( 
.A1(n_2327),
.A2(n_138),
.B1(n_134),
.B2(n_136),
.C(n_139),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2325),
.B(n_138),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2322),
.Y(n_2361)
);

AO22x2_ASAP7_75t_L g2362 ( 
.A1(n_2319),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_2362)
);

AO22x2_ASAP7_75t_L g2363 ( 
.A1(n_2319),
.A2(n_143),
.B1(n_140),
.B2(n_142),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2322),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2322),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2325),
.B(n_143),
.Y(n_2366)
);

NOR2x1_ASAP7_75t_L g2367 ( 
.A(n_2322),
.B(n_144),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2335),
.B(n_2135),
.Y(n_2368)
);

AND2x4_ASAP7_75t_SL g2369 ( 
.A(n_2365),
.B(n_2135),
.Y(n_2369)
);

CKINVDCx6p67_ASAP7_75t_R g2370 ( 
.A(n_2360),
.Y(n_2370)
);

NOR2xp33_ASAP7_75t_L g2371 ( 
.A(n_2366),
.B(n_146),
.Y(n_2371)
);

AO22x1_ASAP7_75t_L g2372 ( 
.A1(n_2367),
.A2(n_2337),
.B1(n_2344),
.B2(n_2336),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2362),
.B(n_147),
.Y(n_2373)
);

INVxp67_ASAP7_75t_L g2374 ( 
.A(n_2363),
.Y(n_2374)
);

AOI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2332),
.A2(n_2074),
.B1(n_2104),
.B2(n_2184),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2331),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2350),
.Y(n_2377)
);

CKINVDCx20_ASAP7_75t_R g2378 ( 
.A(n_2352),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_2353),
.Y(n_2379)
);

AOI21xp33_ASAP7_75t_SL g2380 ( 
.A1(n_2354),
.A2(n_2361),
.B(n_2355),
.Y(n_2380)
);

NOR2x1_ASAP7_75t_L g2381 ( 
.A(n_2364),
.B(n_147),
.Y(n_2381)
);

AOI322xp5_ASAP7_75t_L g2382 ( 
.A1(n_2348),
.A2(n_2357),
.A3(n_2345),
.B1(n_2342),
.B2(n_2340),
.C1(n_2346),
.C2(n_2343),
.Y(n_2382)
);

AOI22xp33_ASAP7_75t_L g2383 ( 
.A1(n_2338),
.A2(n_2184),
.B1(n_2177),
.B2(n_2175),
.Y(n_2383)
);

HB1xp67_ASAP7_75t_L g2384 ( 
.A(n_2334),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_R g2385 ( 
.A(n_2358),
.B(n_148),
.Y(n_2385)
);

OAI21xp33_ASAP7_75t_L g2386 ( 
.A1(n_2347),
.A2(n_2175),
.B(n_2177),
.Y(n_2386)
);

AOI22xp5_ASAP7_75t_L g2387 ( 
.A1(n_2359),
.A2(n_2184),
.B1(n_2177),
.B2(n_2062),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2356),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_SL g2389 ( 
.A(n_2341),
.B(n_148),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2349),
.Y(n_2390)
);

OAI22xp33_ASAP7_75t_SL g2391 ( 
.A1(n_2339),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2333),
.B(n_149),
.Y(n_2392)
);

O2A1O1Ixp33_ASAP7_75t_L g2393 ( 
.A1(n_2351),
.A2(n_153),
.B(n_151),
.C(n_152),
.Y(n_2393)
);

NOR2x1_ASAP7_75t_L g2394 ( 
.A(n_2367),
.B(n_153),
.Y(n_2394)
);

NAND2xp33_ASAP7_75t_SL g2395 ( 
.A(n_2336),
.B(n_154),
.Y(n_2395)
);

OAI22xp5_ASAP7_75t_SL g2396 ( 
.A1(n_2331),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_2396)
);

AOI22xp5_ASAP7_75t_L g2397 ( 
.A1(n_2335),
.A2(n_2184),
.B1(n_2173),
.B2(n_2088),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2367),
.B(n_155),
.Y(n_2398)
);

AOI22xp33_ASAP7_75t_L g2399 ( 
.A1(n_2335),
.A2(n_2184),
.B1(n_2087),
.B2(n_2093),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_R g2400 ( 
.A(n_2331),
.B(n_157),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2362),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2367),
.B(n_157),
.Y(n_2402)
);

OR2x2_ASAP7_75t_L g2403 ( 
.A(n_2360),
.B(n_158),
.Y(n_2403)
);

AOI322xp5_ASAP7_75t_L g2404 ( 
.A1(n_2335),
.A2(n_158),
.A3(n_159),
.B1(n_160),
.B2(n_161),
.C1(n_162),
.C2(n_163),
.Y(n_2404)
);

INVxp67_ASAP7_75t_SL g2405 ( 
.A(n_2381),
.Y(n_2405)
);

NOR2x1p5_ASAP7_75t_L g2406 ( 
.A(n_2373),
.B(n_160),
.Y(n_2406)
);

INVxp33_ASAP7_75t_L g2407 ( 
.A(n_2400),
.Y(n_2407)
);

AND2x4_ASAP7_75t_L g2408 ( 
.A(n_2394),
.B(n_161),
.Y(n_2408)
);

NOR3xp33_ASAP7_75t_L g2409 ( 
.A(n_2380),
.B(n_162),
.C(n_164),
.Y(n_2409)
);

OR2x2_ASAP7_75t_L g2410 ( 
.A(n_2401),
.B(n_164),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2368),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2379),
.Y(n_2412)
);

XOR2xp5_ASAP7_75t_L g2413 ( 
.A(n_2378),
.B(n_166),
.Y(n_2413)
);

NOR2x1p5_ASAP7_75t_L g2414 ( 
.A(n_2390),
.B(n_166),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2384),
.Y(n_2415)
);

AOI22xp33_ASAP7_75t_L g2416 ( 
.A1(n_2379),
.A2(n_2089),
.B1(n_2069),
.B2(n_2105),
.Y(n_2416)
);

INVx1_ASAP7_75t_SL g2417 ( 
.A(n_2395),
.Y(n_2417)
);

NOR2x1_ASAP7_75t_L g2418 ( 
.A(n_2398),
.B(n_167),
.Y(n_2418)
);

BUFx3_ASAP7_75t_L g2419 ( 
.A(n_2379),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2403),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2369),
.Y(n_2421)
);

XNOR2x1_ASAP7_75t_L g2422 ( 
.A(n_2372),
.B(n_167),
.Y(n_2422)
);

INVxp67_ASAP7_75t_SL g2423 ( 
.A(n_2396),
.Y(n_2423)
);

NOR2xp67_ASAP7_75t_L g2424 ( 
.A(n_2374),
.B(n_168),
.Y(n_2424)
);

INVxp67_ASAP7_75t_SL g2425 ( 
.A(n_2402),
.Y(n_2425)
);

NOR2x1_ASAP7_75t_L g2426 ( 
.A(n_2388),
.B(n_169),
.Y(n_2426)
);

NOR2x1p5_ASAP7_75t_L g2427 ( 
.A(n_2370),
.B(n_169),
.Y(n_2427)
);

AOI22xp5_ASAP7_75t_L g2428 ( 
.A1(n_2376),
.A2(n_2082),
.B1(n_2105),
.B2(n_2100),
.Y(n_2428)
);

OR2x2_ASAP7_75t_L g2429 ( 
.A(n_2377),
.B(n_170),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2371),
.Y(n_2430)
);

XNOR2xp5_ASAP7_75t_L g2431 ( 
.A(n_2391),
.B(n_171),
.Y(n_2431)
);

AOI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_2389),
.A2(n_2082),
.B1(n_2100),
.B2(n_2098),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2392),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2387),
.Y(n_2434)
);

NAND4xp75_ASAP7_75t_L g2435 ( 
.A(n_2382),
.B(n_2385),
.C(n_2375),
.D(n_2404),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2397),
.Y(n_2436)
);

NAND4xp75_ASAP7_75t_L g2437 ( 
.A(n_2393),
.B(n_173),
.C(n_171),
.D(n_172),
.Y(n_2437)
);

XNOR2xp5_ASAP7_75t_L g2438 ( 
.A(n_2383),
.B(n_172),
.Y(n_2438)
);

OAI211xp5_ASAP7_75t_L g2439 ( 
.A1(n_2386),
.A2(n_175),
.B(n_173),
.C(n_174),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2399),
.Y(n_2440)
);

HB1xp67_ASAP7_75t_L g2441 ( 
.A(n_2381),
.Y(n_2441)
);

NAND2x1p5_ASAP7_75t_L g2442 ( 
.A(n_2394),
.B(n_174),
.Y(n_2442)
);

NOR4xp75_ASAP7_75t_L g2443 ( 
.A(n_2389),
.B(n_177),
.C(n_175),
.D(n_176),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2379),
.Y(n_2444)
);

NOR2x1_ASAP7_75t_L g2445 ( 
.A(n_2381),
.B(n_176),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2372),
.B(n_178),
.Y(n_2446)
);

NAND4xp75_ASAP7_75t_L g2447 ( 
.A(n_2381),
.B(n_180),
.C(n_178),
.D(n_179),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2373),
.Y(n_2448)
);

INVxp67_ASAP7_75t_SL g2449 ( 
.A(n_2381),
.Y(n_2449)
);

NOR2x1_ASAP7_75t_L g2450 ( 
.A(n_2381),
.B(n_179),
.Y(n_2450)
);

XOR2x2_ASAP7_75t_L g2451 ( 
.A(n_2394),
.B(n_181),
.Y(n_2451)
);

AND3x4_ASAP7_75t_L g2452 ( 
.A(n_2394),
.B(n_181),
.C(n_182),
.Y(n_2452)
);

INVxp67_ASAP7_75t_SL g2453 ( 
.A(n_2381),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2373),
.Y(n_2454)
);

NOR2x1_ASAP7_75t_L g2455 ( 
.A(n_2381),
.B(n_182),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2379),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2373),
.Y(n_2457)
);

AND3x1_ASAP7_75t_L g2458 ( 
.A(n_2394),
.B(n_183),
.C(n_184),
.Y(n_2458)
);

INVx3_ASAP7_75t_L g2459 ( 
.A(n_2379),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2373),
.Y(n_2460)
);

NAND4xp75_ASAP7_75t_L g2461 ( 
.A(n_2381),
.B(n_185),
.C(n_183),
.D(n_184),
.Y(n_2461)
);

NOR2x1_ASAP7_75t_L g2462 ( 
.A(n_2381),
.B(n_185),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2372),
.B(n_186),
.Y(n_2463)
);

AOI221xp5_ASAP7_75t_L g2464 ( 
.A1(n_2415),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.C(n_189),
.Y(n_2464)
);

AOI321xp33_ASAP7_75t_L g2465 ( 
.A1(n_2415),
.A2(n_187),
.A3(n_189),
.B1(n_190),
.B2(n_191),
.C(n_192),
.Y(n_2465)
);

OR2x2_ASAP7_75t_L g2466 ( 
.A(n_2442),
.B(n_190),
.Y(n_2466)
);

AOI21xp33_ASAP7_75t_SL g2467 ( 
.A1(n_2452),
.A2(n_191),
.B(n_192),
.Y(n_2467)
);

AOI211xp5_ASAP7_75t_L g2468 ( 
.A1(n_2439),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2427),
.Y(n_2469)
);

OAI322xp33_ASAP7_75t_SL g2470 ( 
.A1(n_2411),
.A2(n_2421),
.A3(n_2463),
.B1(n_2446),
.B2(n_2456),
.C1(n_2412),
.C2(n_2444),
.Y(n_2470)
);

A2O1A1Ixp33_ASAP7_75t_L g2471 ( 
.A1(n_2424),
.A2(n_196),
.B(n_194),
.C(n_195),
.Y(n_2471)
);

INVxp67_ASAP7_75t_SL g2472 ( 
.A(n_2445),
.Y(n_2472)
);

A2O1A1Ixp33_ASAP7_75t_L g2473 ( 
.A1(n_2459),
.A2(n_2419),
.B(n_2409),
.C(n_2450),
.Y(n_2473)
);

AOI322xp5_ASAP7_75t_L g2474 ( 
.A1(n_2423),
.A2(n_196),
.A3(n_197),
.B1(n_198),
.B2(n_199),
.C1(n_200),
.C2(n_203),
.Y(n_2474)
);

AOI22xp5_ASAP7_75t_L g2475 ( 
.A1(n_2417),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_2475)
);

NOR3xp33_ASAP7_75t_SL g2476 ( 
.A(n_2435),
.B(n_200),
.C(n_203),
.Y(n_2476)
);

NOR3xp33_ASAP7_75t_L g2477 ( 
.A(n_2459),
.B(n_204),
.C(n_205),
.Y(n_2477)
);

OAI211xp5_ASAP7_75t_L g2478 ( 
.A1(n_2455),
.A2(n_2462),
.B(n_2449),
.C(n_2453),
.Y(n_2478)
);

AOI21xp5_ASAP7_75t_L g2479 ( 
.A1(n_2405),
.A2(n_205),
.B(n_206),
.Y(n_2479)
);

O2A1O1Ixp5_ASAP7_75t_L g2480 ( 
.A1(n_2408),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_2480)
);

NAND3xp33_ASAP7_75t_L g2481 ( 
.A(n_2458),
.B(n_207),
.C(n_208),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2413),
.Y(n_2482)
);

OAI22xp33_ASAP7_75t_L g2483 ( 
.A1(n_2410),
.A2(n_2407),
.B1(n_2441),
.B2(n_2440),
.Y(n_2483)
);

NOR3x2_ASAP7_75t_L g2484 ( 
.A(n_2447),
.B(n_209),
.C(n_210),
.Y(n_2484)
);

OAI311xp33_ASAP7_75t_L g2485 ( 
.A1(n_2448),
.A2(n_2460),
.A3(n_2457),
.B1(n_2454),
.C1(n_2433),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_2408),
.B(n_209),
.Y(n_2486)
);

OAI22xp5_ASAP7_75t_L g2487 ( 
.A1(n_2422),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_2487)
);

AOI31xp33_ASAP7_75t_L g2488 ( 
.A1(n_2418),
.A2(n_215),
.A3(n_213),
.B(n_214),
.Y(n_2488)
);

AOI211xp5_ASAP7_75t_L g2489 ( 
.A1(n_2431),
.A2(n_215),
.B(n_213),
.C(n_214),
.Y(n_2489)
);

AND2x4_ASAP7_75t_L g2490 ( 
.A(n_2443),
.B(n_216),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2429),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_2437),
.B(n_216),
.Y(n_2492)
);

NAND3xp33_ASAP7_75t_SL g2493 ( 
.A(n_2434),
.B(n_2420),
.C(n_2430),
.Y(n_2493)
);

INVx1_ASAP7_75t_SL g2494 ( 
.A(n_2451),
.Y(n_2494)
);

AOI22x1_ASAP7_75t_L g2495 ( 
.A1(n_2414),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_2495)
);

A2O1A1Ixp33_ASAP7_75t_L g2496 ( 
.A1(n_2426),
.A2(n_219),
.B(n_217),
.C(n_218),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_2461),
.B(n_220),
.Y(n_2497)
);

NAND4xp25_ASAP7_75t_L g2498 ( 
.A(n_2436),
.B(n_220),
.C(n_221),
.D(n_222),
.Y(n_2498)
);

OAI221xp5_ASAP7_75t_SL g2499 ( 
.A1(n_2438),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.C(n_224),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2406),
.B(n_223),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2425),
.Y(n_2501)
);

A2O1A1Ixp33_ASAP7_75t_L g2502 ( 
.A1(n_2432),
.A2(n_224),
.B(n_225),
.C(n_226),
.Y(n_2502)
);

NOR3xp33_ASAP7_75t_L g2503 ( 
.A(n_2428),
.B(n_225),
.C(n_227),
.Y(n_2503)
);

OAI21xp5_ASAP7_75t_SL g2504 ( 
.A1(n_2416),
.A2(n_227),
.B(n_228),
.Y(n_2504)
);

AOI22xp5_ASAP7_75t_L g2505 ( 
.A1(n_2415),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_2505)
);

NAND4xp75_ASAP7_75t_L g2506 ( 
.A(n_2424),
.B(n_229),
.C(n_230),
.D(n_231),
.Y(n_2506)
);

NAND4xp25_ASAP7_75t_L g2507 ( 
.A(n_2411),
.B(n_231),
.C(n_232),
.D(n_233),
.Y(n_2507)
);

OAI32xp33_ASAP7_75t_L g2508 ( 
.A1(n_2415),
.A2(n_233),
.A3(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_2508)
);

AOI22xp33_ASAP7_75t_L g2509 ( 
.A1(n_2415),
.A2(n_2098),
.B1(n_235),
.B2(n_237),
.Y(n_2509)
);

OA22x2_ASAP7_75t_L g2510 ( 
.A1(n_2452),
.A2(n_234),
.B1(n_237),
.B2(n_238),
.Y(n_2510)
);

XNOR2xp5_ASAP7_75t_L g2511 ( 
.A(n_2413),
.B(n_238),
.Y(n_2511)
);

OAI21xp5_ASAP7_75t_L g2512 ( 
.A1(n_2415),
.A2(n_239),
.B(n_240),
.Y(n_2512)
);

NAND3xp33_ASAP7_75t_L g2513 ( 
.A(n_2409),
.B(n_239),
.C(n_240),
.Y(n_2513)
);

NAND5xp2_ASAP7_75t_L g2514 ( 
.A(n_2411),
.B(n_241),
.C(n_242),
.D(n_243),
.E(n_244),
.Y(n_2514)
);

NOR3xp33_ASAP7_75t_L g2515 ( 
.A(n_2415),
.B(n_242),
.C(n_244),
.Y(n_2515)
);

OAI211xp5_ASAP7_75t_SL g2516 ( 
.A1(n_2415),
.A2(n_245),
.B(n_246),
.C(n_247),
.Y(n_2516)
);

OAI21xp5_ASAP7_75t_L g2517 ( 
.A1(n_2415),
.A2(n_245),
.B(n_246),
.Y(n_2517)
);

INVx1_ASAP7_75t_SL g2518 ( 
.A(n_2408),
.Y(n_2518)
);

NOR2xp33_ASAP7_75t_L g2519 ( 
.A(n_2415),
.B(n_247),
.Y(n_2519)
);

AOI22xp5_ASAP7_75t_L g2520 ( 
.A1(n_2415),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_2520)
);

AOI221xp5_ASAP7_75t_L g2521 ( 
.A1(n_2415),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.C(n_252),
.Y(n_2521)
);

CKINVDCx20_ASAP7_75t_R g2522 ( 
.A(n_2411),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2519),
.B(n_251),
.Y(n_2523)
);

NAND3xp33_ASAP7_75t_L g2524 ( 
.A(n_2489),
.B(n_252),
.C(n_253),
.Y(n_2524)
);

OAI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2481),
.A2(n_254),
.B(n_256),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2495),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2511),
.Y(n_2527)
);

XNOR2x1_ASAP7_75t_L g2528 ( 
.A(n_2506),
.B(n_254),
.Y(n_2528)
);

OAI22xp5_ASAP7_75t_L g2529 ( 
.A1(n_2522),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_2529)
);

XNOR2xp5_ASAP7_75t_L g2530 ( 
.A(n_2484),
.B(n_257),
.Y(n_2530)
);

AND2x4_ASAP7_75t_L g2531 ( 
.A(n_2469),
.B(n_258),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2510),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2466),
.Y(n_2533)
);

XNOR2x1_ASAP7_75t_L g2534 ( 
.A(n_2494),
.B(n_259),
.Y(n_2534)
);

AND2x2_ASAP7_75t_SL g2535 ( 
.A(n_2490),
.B(n_2497),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2488),
.Y(n_2536)
);

HB1xp67_ASAP7_75t_L g2537 ( 
.A(n_2490),
.Y(n_2537)
);

BUFx2_ASAP7_75t_L g2538 ( 
.A(n_2512),
.Y(n_2538)
);

NAND4xp75_ASAP7_75t_L g2539 ( 
.A(n_2476),
.B(n_260),
.C(n_261),
.D(n_262),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2500),
.Y(n_2540)
);

NAND4xp75_ASAP7_75t_L g2541 ( 
.A(n_2492),
.B(n_261),
.C(n_263),
.D(n_264),
.Y(n_2541)
);

NAND4xp75_ASAP7_75t_L g2542 ( 
.A(n_2486),
.B(n_263),
.C(n_264),
.D(n_265),
.Y(n_2542)
);

INVx2_ASAP7_75t_SL g2543 ( 
.A(n_2518),
.Y(n_2543)
);

XNOR2x1_ASAP7_75t_L g2544 ( 
.A(n_2487),
.B(n_265),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2480),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2471),
.Y(n_2546)
);

AOI22xp5_ASAP7_75t_L g2547 ( 
.A1(n_2493),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_2547)
);

AOI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_2472),
.A2(n_267),
.B(n_270),
.Y(n_2548)
);

OAI21xp5_ASAP7_75t_L g2549 ( 
.A1(n_2473),
.A2(n_271),
.B(n_272),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2491),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2496),
.Y(n_2551)
);

XOR2x2_ASAP7_75t_L g2552 ( 
.A(n_2513),
.B(n_272),
.Y(n_2552)
);

OR2x2_ASAP7_75t_L g2553 ( 
.A(n_2498),
.B(n_273),
.Y(n_2553)
);

NOR2x1p5_ASAP7_75t_L g2554 ( 
.A(n_2507),
.B(n_273),
.Y(n_2554)
);

XNOR2x1_ASAP7_75t_L g2555 ( 
.A(n_2482),
.B(n_274),
.Y(n_2555)
);

NOR2x1_ASAP7_75t_L g2556 ( 
.A(n_2478),
.B(n_275),
.Y(n_2556)
);

OR2x2_ASAP7_75t_L g2557 ( 
.A(n_2514),
.B(n_2499),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2465),
.Y(n_2558)
);

AND2x4_ASAP7_75t_L g2559 ( 
.A(n_2501),
.B(n_275),
.Y(n_2559)
);

OA22x2_ASAP7_75t_L g2560 ( 
.A1(n_2504),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_2560)
);

NAND3xp33_ASAP7_75t_L g2561 ( 
.A(n_2468),
.B(n_278),
.C(n_279),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_L g2562 ( 
.A(n_2467),
.B(n_280),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2475),
.Y(n_2563)
);

NAND2x1_ASAP7_75t_L g2564 ( 
.A(n_2479),
.B(n_280),
.Y(n_2564)
);

AND2x4_ASAP7_75t_L g2565 ( 
.A(n_2517),
.B(n_281),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2505),
.Y(n_2566)
);

XNOR2xp5_ASAP7_75t_L g2567 ( 
.A(n_2483),
.B(n_281),
.Y(n_2567)
);

XNOR2x1_ASAP7_75t_L g2568 ( 
.A(n_2520),
.B(n_282),
.Y(n_2568)
);

AND2x2_ASAP7_75t_L g2569 ( 
.A(n_2515),
.B(n_2477),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2516),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2521),
.B(n_282),
.Y(n_2571)
);

XNOR2x1_ASAP7_75t_L g2572 ( 
.A(n_2470),
.B(n_283),
.Y(n_2572)
);

AOI211xp5_ASAP7_75t_L g2573 ( 
.A1(n_2562),
.A2(n_2485),
.B(n_2502),
.C(n_2508),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2567),
.Y(n_2574)
);

OR3x2_ASAP7_75t_L g2575 ( 
.A(n_2553),
.B(n_2558),
.C(n_2536),
.Y(n_2575)
);

NOR3xp33_ASAP7_75t_L g2576 ( 
.A(n_2543),
.B(n_2550),
.C(n_2545),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2567),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2534),
.Y(n_2578)
);

CKINVDCx16_ASAP7_75t_R g2579 ( 
.A(n_2537),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_SL g2580 ( 
.A(n_2547),
.B(n_2464),
.Y(n_2580)
);

OR2x6_ASAP7_75t_L g2581 ( 
.A(n_2564),
.B(n_2503),
.Y(n_2581)
);

HB1xp67_ASAP7_75t_L g2582 ( 
.A(n_2542),
.Y(n_2582)
);

XNOR2xp5_ASAP7_75t_L g2583 ( 
.A(n_2572),
.B(n_2509),
.Y(n_2583)
);

NAND3xp33_ASAP7_75t_SL g2584 ( 
.A(n_2523),
.B(n_2474),
.C(n_283),
.Y(n_2584)
);

OR2x2_ASAP7_75t_L g2585 ( 
.A(n_2528),
.B(n_284),
.Y(n_2585)
);

XOR2xp5_ASAP7_75t_L g2586 ( 
.A(n_2555),
.B(n_284),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2560),
.Y(n_2587)
);

INVx3_ASAP7_75t_SL g2588 ( 
.A(n_2535),
.Y(n_2588)
);

BUFx2_ASAP7_75t_L g2589 ( 
.A(n_2556),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2530),
.Y(n_2590)
);

NAND4xp25_ASAP7_75t_L g2591 ( 
.A(n_2561),
.B(n_285),
.C(n_286),
.D(n_287),
.Y(n_2591)
);

NAND4xp75_ASAP7_75t_L g2592 ( 
.A(n_2546),
.B(n_286),
.C(n_287),
.D(n_288),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2559),
.B(n_289),
.Y(n_2593)
);

OR3x1_ASAP7_75t_L g2594 ( 
.A(n_2570),
.B(n_289),
.C(n_290),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2530),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_SL g2596 ( 
.A(n_2549),
.B(n_290),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_SL g2597 ( 
.A(n_2565),
.B(n_291),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_2525),
.B(n_291),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2548),
.B(n_292),
.Y(n_2599)
);

CKINVDCx16_ASAP7_75t_R g2600 ( 
.A(n_2557),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2539),
.Y(n_2601)
);

BUFx12f_ASAP7_75t_L g2602 ( 
.A(n_2538),
.Y(n_2602)
);

INVx1_ASAP7_75t_SL g2603 ( 
.A(n_2531),
.Y(n_2603)
);

OA22x2_ASAP7_75t_L g2604 ( 
.A1(n_2526),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_2604)
);

AOI22xp33_ASAP7_75t_SL g2605 ( 
.A1(n_2524),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_2605)
);

INVx2_ASAP7_75t_SL g2606 ( 
.A(n_2554),
.Y(n_2606)
);

OA22x2_ASAP7_75t_SL g2607 ( 
.A1(n_2551),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_2607)
);

INVx1_ASAP7_75t_SL g2608 ( 
.A(n_2541),
.Y(n_2608)
);

NOR3xp33_ASAP7_75t_L g2609 ( 
.A(n_2527),
.B(n_2563),
.C(n_2532),
.Y(n_2609)
);

AOI22xp5_ASAP7_75t_SL g2610 ( 
.A1(n_2586),
.A2(n_2604),
.B1(n_2593),
.B2(n_2589),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2594),
.Y(n_2611)
);

OAI21xp5_ASAP7_75t_L g2612 ( 
.A1(n_2576),
.A2(n_2609),
.B(n_2583),
.Y(n_2612)
);

NOR3xp33_ASAP7_75t_SL g2613 ( 
.A(n_2579),
.B(n_2600),
.C(n_2584),
.Y(n_2613)
);

INVx1_ASAP7_75t_SL g2614 ( 
.A(n_2592),
.Y(n_2614)
);

HB1xp67_ASAP7_75t_L g2615 ( 
.A(n_2581),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2607),
.Y(n_2616)
);

OR3x2_ASAP7_75t_L g2617 ( 
.A(n_2585),
.B(n_2540),
.C(n_2552),
.Y(n_2617)
);

AND2x2_ASAP7_75t_SL g2618 ( 
.A(n_2587),
.B(n_2533),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2599),
.Y(n_2619)
);

OAI21x1_ASAP7_75t_SL g2620 ( 
.A1(n_2601),
.A2(n_2568),
.B(n_2544),
.Y(n_2620)
);

HB1xp67_ASAP7_75t_L g2621 ( 
.A(n_2581),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2597),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2605),
.B(n_2569),
.Y(n_2623)
);

HB1xp67_ASAP7_75t_L g2624 ( 
.A(n_2582),
.Y(n_2624)
);

AOI22xp5_ASAP7_75t_L g2625 ( 
.A1(n_2602),
.A2(n_2566),
.B1(n_2571),
.B2(n_2529),
.Y(n_2625)
);

BUFx2_ASAP7_75t_L g2626 ( 
.A(n_2588),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2603),
.B(n_297),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2608),
.B(n_298),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2596),
.Y(n_2629)
);

XOR2x1_ASAP7_75t_L g2630 ( 
.A(n_2578),
.B(n_299),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2573),
.B(n_300),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2575),
.Y(n_2632)
);

NOR3x2_ASAP7_75t_L g2633 ( 
.A(n_2630),
.B(n_2606),
.C(n_2574),
.Y(n_2633)
);

AOI22xp5_ASAP7_75t_L g2634 ( 
.A1(n_2626),
.A2(n_2577),
.B1(n_2591),
.B2(n_2595),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2627),
.B(n_2590),
.Y(n_2635)
);

OAI221xp5_ASAP7_75t_L g2636 ( 
.A1(n_2612),
.A2(n_2598),
.B1(n_2580),
.B2(n_303),
.C(n_304),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2616),
.Y(n_2637)
);

OR3x1_ASAP7_75t_L g2638 ( 
.A(n_2611),
.B(n_300),
.C(n_302),
.Y(n_2638)
);

INVx1_ASAP7_75t_SL g2639 ( 
.A(n_2628),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2631),
.Y(n_2640)
);

OAI22x1_ASAP7_75t_L g2641 ( 
.A1(n_2625),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2615),
.Y(n_2642)
);

XNOR2xp5_ASAP7_75t_L g2643 ( 
.A(n_2610),
.B(n_305),
.Y(n_2643)
);

INVxp67_ASAP7_75t_L g2644 ( 
.A(n_2621),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2624),
.Y(n_2645)
);

NAND3xp33_ASAP7_75t_SL g2646 ( 
.A(n_2614),
.B(n_305),
.C(n_306),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2618),
.B(n_306),
.Y(n_2647)
);

NOR3xp33_ASAP7_75t_SL g2648 ( 
.A(n_2623),
.B(n_307),
.C(n_308),
.Y(n_2648)
);

NOR3xp33_ASAP7_75t_L g2649 ( 
.A(n_2632),
.B(n_308),
.C(n_309),
.Y(n_2649)
);

AND2x2_ASAP7_75t_L g2650 ( 
.A(n_2613),
.B(n_310),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_SL g2651 ( 
.A(n_2642),
.B(n_2622),
.Y(n_2651)
);

OAI21xp5_ASAP7_75t_L g2652 ( 
.A1(n_2644),
.A2(n_2629),
.B(n_2619),
.Y(n_2652)
);

AOI21xp5_ASAP7_75t_L g2653 ( 
.A1(n_2645),
.A2(n_2650),
.B(n_2643),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2647),
.Y(n_2654)
);

AOI22xp5_ASAP7_75t_SL g2655 ( 
.A1(n_2641),
.A2(n_2617),
.B1(n_2620),
.B2(n_314),
.Y(n_2655)
);

OAI22xp5_ASAP7_75t_L g2656 ( 
.A1(n_2638),
.A2(n_311),
.B1(n_312),
.B2(n_315),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2637),
.Y(n_2657)
);

OAI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2634),
.A2(n_311),
.B1(n_312),
.B2(n_315),
.Y(n_2658)
);

AOI22xp5_ASAP7_75t_L g2659 ( 
.A1(n_2646),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_2659)
);

AOI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_2640),
.A2(n_316),
.B1(n_317),
.B2(n_319),
.Y(n_2660)
);

CKINVDCx20_ASAP7_75t_R g2661 ( 
.A(n_2651),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2657),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2656),
.Y(n_2663)
);

AND2x4_ASAP7_75t_L g2664 ( 
.A(n_2652),
.B(n_2648),
.Y(n_2664)
);

BUFx4f_ASAP7_75t_SL g2665 ( 
.A(n_2654),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2658),
.Y(n_2666)
);

AO221x1_ASAP7_75t_L g2667 ( 
.A1(n_2663),
.A2(n_2655),
.B1(n_2633),
.B2(n_2636),
.C(n_2659),
.Y(n_2667)
);

OAI21xp5_ASAP7_75t_L g2668 ( 
.A1(n_2661),
.A2(n_2653),
.B(n_2635),
.Y(n_2668)
);

AOI222xp33_ASAP7_75t_L g2669 ( 
.A1(n_2665),
.A2(n_2639),
.B1(n_2660),
.B2(n_2649),
.C1(n_323),
.C2(n_324),
.Y(n_2669)
);

AOI222xp33_ASAP7_75t_L g2670 ( 
.A1(n_2662),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.C1(n_323),
.C2(n_324),
.Y(n_2670)
);

OAI22xp5_ASAP7_75t_SL g2671 ( 
.A1(n_2668),
.A2(n_2664),
.B1(n_2666),
.B2(n_327),
.Y(n_2671)
);

INVxp67_ASAP7_75t_L g2672 ( 
.A(n_2669),
.Y(n_2672)
);

OR3x2_ASAP7_75t_L g2673 ( 
.A(n_2667),
.B(n_321),
.C(n_325),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_L g2674 ( 
.A(n_2671),
.B(n_2672),
.Y(n_2674)
);

OAI221xp5_ASAP7_75t_R g2675 ( 
.A1(n_2674),
.A2(n_2673),
.B1(n_2670),
.B2(n_329),
.C(n_331),
.Y(n_2675)
);

AOI22xp33_ASAP7_75t_L g2676 ( 
.A1(n_2675),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.Y(n_2676)
);

AOI21xp5_ASAP7_75t_L g2677 ( 
.A1(n_2676),
.A2(n_331),
.B(n_332),
.Y(n_2677)
);

AOI211xp5_ASAP7_75t_L g2678 ( 
.A1(n_2677),
.A2(n_333),
.B(n_334),
.C(n_335),
.Y(n_2678)
);


endmodule