module real_aes_8951_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g292 ( .A(n_0), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g108 ( .A1(n_1), .A2(n_71), .B1(n_109), .B2(n_114), .Y(n_108) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_2), .A2(n_29), .B1(n_203), .B2(n_226), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_3), .B(n_232), .Y(n_304) );
INVx1_ASAP7_75t_L g185 ( .A(n_4), .Y(n_185) );
AND2x6_ASAP7_75t_L g218 ( .A(n_4), .B(n_183), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_4), .B(n_502), .Y(n_501) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_5), .A2(n_23), .B1(n_91), .B2(n_96), .Y(n_99) );
INVx1_ASAP7_75t_L g199 ( .A(n_6), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_7), .B(n_208), .Y(n_240) );
AOI22xp5_ASAP7_75t_SL g497 ( .A1(n_7), .A2(n_80), .B1(n_81), .B2(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_7), .Y(n_498) );
INVx1_ASAP7_75t_L g284 ( .A(n_8), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_9), .B(n_233), .Y(n_271) );
AO32x2_ASAP7_75t_L g254 ( .A1(n_10), .A2(n_231), .A3(n_232), .B1(n_255), .B2(n_259), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_11), .B(n_203), .Y(n_244) );
INVx1_ASAP7_75t_L g508 ( .A(n_11), .Y(n_508) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_12), .A2(n_25), .B1(n_91), .B2(n_92), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_13), .B(n_233), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_14), .A2(n_38), .B1(n_203), .B2(n_226), .Y(n_258) );
AOI22xp33_ASAP7_75t_SL g229 ( .A1(n_15), .A2(n_59), .B1(n_203), .B2(n_208), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_16), .B(n_203), .Y(n_214) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_17), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_18), .B(n_195), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_19), .A2(n_27), .B1(n_120), .B2(n_126), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g168 ( .A1(n_20), .A2(n_45), .B1(n_169), .B2(n_170), .Y(n_168) );
INVx1_ASAP7_75t_L g170 ( .A(n_20), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_21), .B(n_195), .Y(n_219) );
INVx2_ASAP7_75t_L g205 ( .A(n_22), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_24), .B(n_203), .Y(n_308) );
OAI221xp5_ASAP7_75t_L g176 ( .A1(n_25), .A2(n_42), .B1(n_56), .B2(n_177), .C(n_178), .Y(n_176) );
INVxp67_ASAP7_75t_L g179 ( .A(n_25), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_26), .B(n_195), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_28), .A2(n_80), .B1(n_81), .B2(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_28), .Y(n_510) );
AOI222xp33_ASAP7_75t_L g152 ( .A1(n_30), .A2(n_33), .B1(n_75), .B2(n_153), .C1(n_155), .C2(n_159), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_31), .B(n_203), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_32), .A2(n_43), .B1(n_130), .B2(n_133), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_34), .A2(n_67), .B1(n_226), .B2(n_227), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_35), .B(n_203), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_36), .B(n_203), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_37), .B(n_290), .Y(n_303) );
AOI22xp33_ASAP7_75t_SL g275 ( .A1(n_39), .A2(n_46), .B1(n_203), .B2(n_208), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_40), .B(n_203), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_41), .B(n_203), .Y(n_239) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_42), .A2(n_64), .B1(n_91), .B2(n_92), .Y(n_90) );
INVxp67_ASAP7_75t_L g180 ( .A(n_42), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_44), .A2(n_63), .B1(n_139), .B2(n_142), .Y(n_138) );
INVx1_ASAP7_75t_L g169 ( .A(n_45), .Y(n_169) );
INVx1_ASAP7_75t_L g183 ( .A(n_47), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_48), .B(n_203), .Y(n_293) );
INVx1_ASAP7_75t_L g198 ( .A(n_49), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_50), .A2(n_80), .B1(n_81), .B2(n_163), .Y(n_79) );
INVx1_ASAP7_75t_SL g163 ( .A(n_50), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_51), .Y(n_177) );
AO32x2_ASAP7_75t_L g223 ( .A1(n_52), .A2(n_224), .A3(n_230), .B1(n_231), .B2(n_232), .Y(n_223) );
INVx1_ASAP7_75t_L g311 ( .A(n_53), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g84 ( .A1(n_54), .A2(n_58), .B1(n_85), .B2(n_102), .Y(n_84) );
INVx1_ASAP7_75t_L g206 ( .A(n_55), .Y(n_206) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_56), .A2(n_70), .B1(n_91), .B2(n_96), .Y(n_95) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_57), .A2(n_167), .B1(n_168), .B2(n_171), .Y(n_166) );
INVx1_ASAP7_75t_L g171 ( .A(n_57), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_57), .B(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_60), .B(n_226), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_61), .A2(n_69), .B1(n_145), .B2(n_149), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_62), .B(n_208), .Y(n_215) );
INVx2_ASAP7_75t_L g196 ( .A(n_65), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_66), .B(n_208), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_68), .A2(n_76), .B1(n_208), .B2(n_209), .Y(n_274) );
OAI22xp5_ASAP7_75t_SL g164 ( .A1(n_72), .A2(n_165), .B1(n_166), .B2(n_172), .Y(n_164) );
INVx1_ASAP7_75t_L g172 ( .A(n_72), .Y(n_172) );
INVx1_ASAP7_75t_L g91 ( .A(n_73), .Y(n_91) );
INVx1_ASAP7_75t_L g93 ( .A(n_73), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_74), .B(n_208), .Y(n_309) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_173), .B1(n_186), .B2(n_490), .C(n_496), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_164), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND4xp75_ASAP7_75t_SL g82 ( .A(n_83), .B(n_118), .C(n_137), .D(n_152), .Y(n_82) );
AND2x2_ASAP7_75t_L g83 ( .A(n_84), .B(n_108), .Y(n_83) );
BUFx3_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_97), .Y(n_87) );
AND2x4_ASAP7_75t_L g112 ( .A(n_88), .B(n_113), .Y(n_112) );
AND2x6_ASAP7_75t_L g123 ( .A(n_88), .B(n_124), .Y(n_123) );
AND2x6_ASAP7_75t_L g154 ( .A(n_88), .B(n_151), .Y(n_154) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_94), .Y(n_88) );
AND2x2_ASAP7_75t_L g128 ( .A(n_89), .B(n_95), .Y(n_128) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x2_ASAP7_75t_L g106 ( .A(n_90), .B(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_90), .B(n_95), .Y(n_117) );
AND2x2_ASAP7_75t_L g148 ( .A(n_90), .B(n_99), .Y(n_148) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g96 ( .A(n_93), .Y(n_96) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g107 ( .A(n_95), .Y(n_107) );
INVx1_ASAP7_75t_L g158 ( .A(n_95), .Y(n_158) );
AND2x2_ASAP7_75t_L g105 ( .A(n_97), .B(n_106), .Y(n_105) );
AND2x4_ASAP7_75t_L g115 ( .A(n_97), .B(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g127 ( .A(n_97), .B(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_100), .Y(n_97) );
AND2x2_ASAP7_75t_L g113 ( .A(n_98), .B(n_101), .Y(n_113) );
OR2x2_ASAP7_75t_L g125 ( .A(n_98), .B(n_101), .Y(n_125) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g151 ( .A(n_99), .B(n_101), .Y(n_151) );
AND2x2_ASAP7_75t_L g157 ( .A(n_100), .B(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g136 ( .A(n_101), .Y(n_136) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g132 ( .A(n_106), .B(n_113), .Y(n_132) );
INVx1_ASAP7_75t_L g150 ( .A(n_107), .Y(n_150) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x6_ASAP7_75t_L g143 ( .A(n_113), .B(n_128), .Y(n_143) );
BUFx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x6_ASAP7_75t_L g135 ( .A(n_117), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_129), .Y(n_118) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx11_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g141 ( .A(n_124), .B(n_128), .Y(n_141) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx8_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx6_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
AND2x2_ASAP7_75t_SL g137 ( .A(n_138), .B(n_144), .Y(n_137) );
INVx5_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx4_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x4_ASAP7_75t_L g156 ( .A(n_148), .B(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g161 ( .A(n_148), .B(n_162), .Y(n_161) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx4f_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g162 ( .A(n_158), .Y(n_162) );
BUFx4f_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
BUFx12f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_166), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_168), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
AND3x1_ASAP7_75t_SL g175 ( .A(n_176), .B(n_181), .C(n_184), .Y(n_175) );
INVxp67_ASAP7_75t_L g502 ( .A(n_176), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx1_ASAP7_75t_SL g503 ( .A(n_181), .Y(n_503) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_181), .A2(n_495), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g514 ( .A(n_181), .Y(n_514) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_182), .B(n_185), .Y(n_507) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OR2x2_ASAP7_75t_SL g513 ( .A(n_184), .B(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
OR2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_411), .Y(n_186) );
NAND3xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_360), .C(n_402), .Y(n_187) );
AOI211xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_265), .B(n_314), .C(n_336), .Y(n_188) );
OAI211xp5_ASAP7_75t_SL g189 ( .A1(n_190), .A2(n_220), .B(n_248), .C(n_260), .Y(n_189) );
INVxp67_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_191), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g423 ( .A(n_191), .B(n_340), .Y(n_423) );
BUFx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g325 ( .A(n_192), .B(n_251), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_192), .B(n_236), .Y(n_442) );
INVx1_ASAP7_75t_L g460 ( .A(n_192), .Y(n_460) );
AND2x2_ASAP7_75t_L g469 ( .A(n_192), .B(n_357), .Y(n_469) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OR2x2_ASAP7_75t_L g352 ( .A(n_193), .B(n_236), .Y(n_352) );
AND2x2_ASAP7_75t_L g410 ( .A(n_193), .B(n_357), .Y(n_410) );
INVx1_ASAP7_75t_L g454 ( .A(n_193), .Y(n_454) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OR2x2_ASAP7_75t_L g331 ( .A(n_194), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g339 ( .A(n_194), .Y(n_339) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_194), .Y(n_379) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_200), .B(n_219), .Y(n_194) );
INVx2_ASAP7_75t_L g230 ( .A(n_195), .Y(n_230) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_195), .A2(n_237), .B(n_247), .Y(n_236) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_196), .B(n_197), .Y(n_195) );
AND2x2_ASAP7_75t_L g233 ( .A(n_196), .B(n_197), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_213), .B(n_218), .Y(n_200) );
O2A1O1Ixp5_ASAP7_75t_SL g201 ( .A1(n_202), .A2(n_206), .B(n_207), .C(n_210), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g226 ( .A(n_204), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_204), .Y(n_227) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g209 ( .A(n_205), .Y(n_209) );
INVx1_ASAP7_75t_L g291 ( .A(n_205), .Y(n_291) );
INVx2_ASAP7_75t_L g285 ( .A(n_208), .Y(n_285) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g257 ( .A(n_210), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_210), .A2(n_299), .B(n_300), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_210), .A2(n_308), .B(n_309), .Y(n_307) );
INVx5_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OAI22xp5_ASAP7_75t_SL g224 ( .A1(n_211), .A2(n_225), .B1(n_228), .B2(n_229), .Y(n_224) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_212), .Y(n_217) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_212), .Y(n_228) );
INVx1_ASAP7_75t_L g242 ( .A(n_212), .Y(n_242) );
AND2x2_ASAP7_75t_L g495 ( .A(n_212), .B(n_291), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_216), .Y(n_213) );
INVx1_ASAP7_75t_L g287 ( .A(n_216), .Y(n_287) );
INVx4_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx3_ASAP7_75t_L g231 ( .A(n_218), .Y(n_231) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_218), .A2(n_238), .B(n_243), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g282 ( .A1(n_218), .A2(n_283), .B(n_288), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_218), .A2(n_298), .B(n_301), .Y(n_297) );
AND2x4_ASAP7_75t_L g494 ( .A(n_218), .B(n_495), .Y(n_494) );
INVxp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_234), .Y(n_221) );
AND2x2_ASAP7_75t_L g318 ( .A(n_222), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g351 ( .A(n_222), .Y(n_351) );
OR2x2_ASAP7_75t_L g477 ( .A(n_222), .B(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_222), .B(n_236), .Y(n_481) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g251 ( .A(n_223), .Y(n_251) );
INVx1_ASAP7_75t_L g263 ( .A(n_223), .Y(n_263) );
AND2x2_ASAP7_75t_L g340 ( .A(n_223), .B(n_253), .Y(n_340) );
AND2x2_ASAP7_75t_L g380 ( .A(n_223), .B(n_254), .Y(n_380) );
INVx2_ASAP7_75t_L g246 ( .A(n_228), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_228), .A2(n_256), .B1(n_257), .B2(n_258), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_228), .A2(n_257), .B1(n_274), .B2(n_275), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g272 ( .A(n_231), .B(n_273), .C(n_276), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_231), .A2(n_307), .B(n_310), .Y(n_306) );
INVx4_ASAP7_75t_L g276 ( .A(n_232), .Y(n_276) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_232), .A2(n_297), .B(n_304), .Y(n_296) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g259 ( .A(n_233), .Y(n_259) );
INVxp67_ASAP7_75t_L g422 ( .A(n_234), .Y(n_422) );
AND2x4_ASAP7_75t_L g447 ( .A(n_234), .B(n_340), .Y(n_447) );
BUFx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_SL g338 ( .A(n_235), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g252 ( .A(n_236), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g326 ( .A(n_236), .B(n_254), .Y(n_326) );
INVx1_ASAP7_75t_L g332 ( .A(n_236), .Y(n_332) );
INVx2_ASAP7_75t_L g358 ( .A(n_236), .Y(n_358) );
AND2x2_ASAP7_75t_L g374 ( .A(n_236), .B(n_375), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_241), .Y(n_238) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_246), .Y(n_243) );
O2A1O1Ixp5_ASAP7_75t_L g310 ( .A1(n_246), .A2(n_289), .B(n_311), .C(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_249), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_252), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
BUFx2_ASAP7_75t_L g329 ( .A(n_251), .Y(n_329) );
AND2x2_ASAP7_75t_L g437 ( .A(n_251), .B(n_253), .Y(n_437) );
AND2x2_ASAP7_75t_L g354 ( .A(n_252), .B(n_339), .Y(n_354) );
AND2x2_ASAP7_75t_L g453 ( .A(n_252), .B(n_454), .Y(n_453) );
NOR2xp67_ASAP7_75t_L g375 ( .A(n_253), .B(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g478 ( .A(n_253), .B(n_339), .Y(n_478) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
BUFx2_ASAP7_75t_L g264 ( .A(n_254), .Y(n_264) );
AND2x2_ASAP7_75t_L g357 ( .A(n_254), .B(n_358), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g288 ( .A1(n_257), .A2(n_289), .B(n_292), .C(n_293), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_257), .A2(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g281 ( .A(n_259), .Y(n_281) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
AND2x2_ASAP7_75t_L g403 ( .A(n_262), .B(n_338), .Y(n_403) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_263), .B(n_339), .Y(n_388) );
INVx2_ASAP7_75t_L g387 ( .A(n_264), .Y(n_387) );
OAI222xp33_ASAP7_75t_L g391 ( .A1(n_264), .A2(n_331), .B1(n_392), .B2(n_394), .C1(n_395), .C2(n_398), .Y(n_391) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_277), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g316 ( .A(n_269), .Y(n_316) );
OR2x2_ASAP7_75t_L g427 ( .A(n_269), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g349 ( .A(n_270), .Y(n_349) );
NOR2x1_ASAP7_75t_L g400 ( .A(n_270), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g406 ( .A(n_270), .B(n_320), .Y(n_406) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g367 ( .A(n_271), .Y(n_367) );
AO21x1_ASAP7_75t_L g366 ( .A1(n_273), .A2(n_276), .B(n_367), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_277), .A2(n_370), .B1(n_409), .B2(n_410), .Y(n_408) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_295), .Y(n_277) );
INVx3_ASAP7_75t_L g342 ( .A(n_278), .Y(n_342) );
OR2x2_ASAP7_75t_L g475 ( .A(n_278), .B(n_351), .Y(n_475) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g348 ( .A(n_279), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g364 ( .A(n_279), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g372 ( .A(n_279), .B(n_320), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_279), .B(n_296), .Y(n_428) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g319 ( .A(n_280), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g323 ( .A(n_280), .B(n_296), .Y(n_323) );
AND2x2_ASAP7_75t_L g399 ( .A(n_280), .B(n_346), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_280), .B(n_305), .Y(n_439) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_294), .Y(n_280) );
OA21x2_ASAP7_75t_L g305 ( .A1(n_281), .A2(n_306), .B(n_313), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B(n_286), .C(n_287), .Y(n_283) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_295), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g355 ( .A(n_295), .B(n_316), .Y(n_355) );
AND2x2_ASAP7_75t_L g359 ( .A(n_295), .B(n_349), .Y(n_359) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_305), .Y(n_295) );
INVx3_ASAP7_75t_L g320 ( .A(n_296), .Y(n_320) );
AND2x2_ASAP7_75t_L g345 ( .A(n_296), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g480 ( .A(n_296), .B(n_463), .Y(n_480) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_305), .Y(n_334) );
INVx2_ASAP7_75t_L g346 ( .A(n_305), .Y(n_346) );
AND2x2_ASAP7_75t_L g390 ( .A(n_305), .B(n_366), .Y(n_390) );
INVx1_ASAP7_75t_L g433 ( .A(n_305), .Y(n_433) );
OR2x2_ASAP7_75t_L g464 ( .A(n_305), .B(n_366), .Y(n_464) );
AND2x2_ASAP7_75t_L g484 ( .A(n_305), .B(n_320), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B(n_321), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g322 ( .A(n_316), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_316), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g441 ( .A(n_318), .Y(n_441) );
INVx2_ASAP7_75t_SL g335 ( .A(n_319), .Y(n_335) );
AND2x2_ASAP7_75t_L g455 ( .A(n_319), .B(n_349), .Y(n_455) );
INVx2_ASAP7_75t_L g401 ( .A(n_320), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_320), .B(n_433), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_324), .B1(n_327), .B2(n_333), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_323), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_SL g489 ( .A(n_323), .Y(n_489) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g414 ( .A(n_325), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_325), .B(n_357), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_326), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g430 ( .A(n_326), .B(n_379), .Y(n_430) );
INVx2_ASAP7_75t_L g486 ( .A(n_326), .Y(n_486) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x2_ASAP7_75t_L g356 ( .A(n_329), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_329), .B(n_374), .Y(n_407) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_331), .B(n_351), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g468 ( .A(n_334), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_SL g418 ( .A1(n_335), .A2(n_419), .B(n_421), .C(n_424), .Y(n_418) );
OR2x2_ASAP7_75t_L g445 ( .A(n_335), .B(n_349), .Y(n_445) );
OAI221xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_341), .B1(n_343), .B2(n_350), .C(n_353), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_338), .B(n_340), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_338), .B(n_387), .Y(n_394) );
AND2x2_ASAP7_75t_L g436 ( .A(n_338), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g472 ( .A(n_338), .Y(n_472) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_339), .Y(n_363) );
INVx1_ASAP7_75t_L g376 ( .A(n_339), .Y(n_376) );
NOR2xp67_ASAP7_75t_L g396 ( .A(n_342), .B(n_397), .Y(n_396) );
INVxp67_ASAP7_75t_L g450 ( .A(n_342), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_342), .B(n_390), .Y(n_466) );
INVx2_ASAP7_75t_L g452 ( .A(n_343), .Y(n_452) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_347), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g393 ( .A(n_345), .B(n_364), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_L g402 ( .A1(n_345), .A2(n_361), .B(n_403), .C(n_404), .Y(n_402) );
AND2x2_ASAP7_75t_L g371 ( .A(n_346), .B(n_366), .Y(n_371) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_350), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
OR2x2_ASAP7_75t_L g419 ( .A(n_351), .B(n_420), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_356), .B2(n_359), .Y(n_353) );
INVx1_ASAP7_75t_L g473 ( .A(n_355), .Y(n_473) );
INVx1_ASAP7_75t_L g420 ( .A(n_357), .Y(n_420) );
INVx1_ASAP7_75t_L g471 ( .A(n_359), .Y(n_471) );
AOI211xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_364), .B(n_368), .C(n_391), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g383 ( .A(n_363), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g434 ( .A(n_364), .Y(n_434) );
AND2x2_ASAP7_75t_L g483 ( .A(n_364), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI21xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_373), .B(n_381), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVx2_ASAP7_75t_L g397 ( .A(n_371), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_371), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g389 ( .A(n_372), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g465 ( .A(n_372), .Y(n_465) );
OAI32xp33_ASAP7_75t_L g476 ( .A1(n_372), .A2(n_424), .A3(n_431), .B1(n_472), .B2(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_SL g373 ( .A(n_374), .B(n_377), .Y(n_373) );
INVx1_ASAP7_75t_SL g444 ( .A(n_374), .Y(n_444) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g384 ( .A(n_380), .Y(n_384) );
OAI21xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_385), .B(n_389), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g456 ( .A1(n_383), .A2(n_431), .B1(n_457), .B2(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_387), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g424 ( .A(n_390), .Y(n_424) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g417 ( .A(n_401), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B(n_408), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_410), .A2(n_452), .B1(n_453), .B2(n_455), .C(n_456), .Y(n_451) );
NAND5xp2_ASAP7_75t_L g411 ( .A(n_412), .B(n_435), .C(n_451), .D(n_461), .E(n_479), .Y(n_411) );
AOI211xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_415), .B(n_418), .C(n_425), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g482 ( .A(n_419), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_429), .B2(n_431), .Y(n_425) );
INVx1_ASAP7_75t_SL g458 ( .A(n_428), .Y(n_458) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI322xp33_ASAP7_75t_L g440 ( .A1(n_431), .A2(n_441), .A3(n_442), .B1(n_443), .B2(n_444), .C1(n_445), .C2(n_446), .Y(n_440) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g443 ( .A(n_433), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_433), .B(n_458), .Y(n_457) );
AOI211xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_438), .B(n_440), .C(n_448), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp33_ASAP7_75t_L g470 ( .A1(n_444), .A2(n_471), .B1(n_472), .B2(n_473), .Y(n_470) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g487 ( .A(n_454), .Y(n_487) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_469), .B1(n_470), .B2(n_474), .C(n_476), .Y(n_461) );
OAI211xp5_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_465), .B(n_466), .C(n_467), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g488 ( .A(n_464), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_482), .B2(n_483), .C(n_485), .Y(n_479) );
AOI21xp33_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_487), .B(n_488), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OAI322xp33_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_499), .A3(n_503), .B1(n_504), .B2(n_508), .C1(n_509), .C2(n_511), .Y(n_496) );
INVx1_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
endmodule