module real_jpeg_32192_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_553;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_572;
wire n_405;
wire n_412;
wire n_548;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_0),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_0),
.Y(n_374)
);

BUFx12f_ASAP7_75t_L g509 ( 
.A(n_0),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_1),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_1),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_1),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_1),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_1),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g327 ( 
.A(n_1),
.B(n_213),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_1),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_1),
.B(n_372),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_2),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_3),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_3),
.B(n_302),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_3),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_3),
.B(n_334),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_3),
.B(n_322),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_3),
.B(n_460),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_3),
.B(n_372),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_4),
.A2(n_13),
.B1(n_21),
.B2(n_24),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_5),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_5),
.B(n_184),
.Y(n_183)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_5),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_5),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_SL g382 ( 
.A(n_5),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_5),
.B(n_38),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_5),
.B(n_463),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_6),
.B(n_81),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g137 ( 
.A(n_6),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_6),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_6),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_6),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_6),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_6),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_6),
.B(n_314),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_7),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_8),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_9),
.Y(n_96)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_9),
.Y(n_512)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_10),
.Y(n_214)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_10),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_L g200 ( 
.A(n_11),
.B(n_201),
.Y(n_200)
);

NAND2x1_ASAP7_75t_L g306 ( 
.A(n_11),
.B(n_41),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_11),
.B(n_334),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_11),
.B(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_11),
.B(n_475),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_SL g510 ( 
.A(n_11),
.B(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_11),
.B(n_518),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_12),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_12),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_12),
.B(n_48),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_12),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_12),
.B(n_66),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_12),
.B(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_12),
.B(n_532),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_14),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_14),
.B(n_94),
.Y(n_93)
);

NAND2x1_ASAP7_75t_SL g132 ( 
.A(n_14),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_14),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_14),
.B(n_44),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_14),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_14),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_14),
.B(n_569),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_15),
.Y(n_135)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_15),
.Y(n_324)
);

NAND2x1_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_16),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_16),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_16),
.B(n_59),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_16),
.B(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_16),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_17),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_17),
.Y(n_239)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_17),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_18),
.B(n_99),
.Y(n_98)
);

NAND2x1_ASAP7_75t_L g186 ( 
.A(n_18),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_18),
.B(n_216),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_18),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_18),
.B(n_437),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_18),
.B(n_480),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_18),
.B(n_487),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_18),
.B(n_507),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_19),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_19),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_19),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_19),
.B(n_245),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_19),
.B(n_94),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_19),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_19),
.B(n_372),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_561),
.B2(n_578),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_285),
.B(n_556),
.Y(n_26)
);

NOR2x1_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_254),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_223),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_167),
.Y(n_29)
);

NOR2xp67_ASAP7_75t_SL g558 ( 
.A(n_30),
.B(n_167),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_105),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_31),
.B(n_106),
.C(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_56),
.C(n_76),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_34),
.B(n_56),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_46),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_36),
.B(n_47),
.C(n_51),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.C(n_43),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_37),
.A2(n_43),
.B1(n_97),
.B2(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_37),
.A2(n_103),
.B1(n_111),
.B2(n_116),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_39),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_39),
.Y(n_460)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_39),
.Y(n_488)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_41),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_42),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_42),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_42),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_42),
.Y(n_281)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_42),
.Y(n_418)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_43),
.A2(n_93),
.B1(n_97),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_57),
.C(n_69),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_47),
.B(n_70),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_50),
.Y(n_218)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_53),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_53),
.Y(n_570)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_54),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_57),
.B(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.C(n_65),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_58),
.B(n_62),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_61),
.Y(n_303)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_65),
.B(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_68),
.Y(n_193)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_77),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_92),
.C(n_101),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_78),
.B(n_92),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_86),
.Y(n_78)
);

XNOR2x1_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_80),
.B(n_83),
.C(n_86),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_82),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_85),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_88),
.B(n_309),
.Y(n_456)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g518 ( 
.A(n_90),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_91),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_98),
.Y(n_92)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_93),
.Y(n_180)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_96),
.Y(n_369)
);

XNOR2x1_ASAP7_75t_L g178 ( 
.A(n_98),
.B(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_101),
.B(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_116),
.C(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_140),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_123),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_107),
.B(n_124),
.C(n_127),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_117),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_109),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_109),
.A2(n_115),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_109),
.B(n_116),
.C(n_117),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_109),
.B(n_267),
.C(n_268),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_111),
.Y(n_116)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp67_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.C(n_136),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_162),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_136),
.B1(n_137),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_140),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_160),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_141)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

XNOR2x1_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_154),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_148),
.B1(n_149),
.B2(n_153),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_147),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_148),
.B(n_153),
.C(n_154),
.Y(n_240)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_151),
.Y(n_441)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_152),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_156),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_158),
.B(n_159),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_158),
.B(n_159),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_160),
.A2(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_165),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_R g167 ( 
.A(n_168),
.B(n_171),
.C(n_174),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_171),
.Y(n_346)
);

XNOR2x2_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_175),
.B(n_345),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_198),
.C(n_220),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_196),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_177),
.B(n_181),
.C(n_196),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_181),
.Y(n_357)
);

OAI21x1_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_189),
.B(n_194),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_186),
.B(n_195),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_189),
.Y(n_387)
);

INVx3_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_196),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_198),
.B(n_221),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_209),
.B(n_219),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.C(n_207),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_200),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_SL g339 ( 
.A(n_200),
.B(n_204),
.C(n_207),
.Y(n_339)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_204),
.A2(n_207),
.B1(n_208),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_204),
.Y(n_297)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

NAND2xp33_ASAP7_75t_SL g219 ( 
.A(n_210),
.B(n_215),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_210),
.B(n_215),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_210),
.B(n_215),
.Y(n_340)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_214),
.Y(n_385)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_214),
.Y(n_481)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_223),
.A2(n_558),
.B(n_559),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_224),
.B(n_226),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_251),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_229),
.C(n_251),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_241),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_230),
.B(n_250),
.C(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_240),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_236),
.C(n_240),
.Y(n_258)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_249),
.B2(n_250),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_267),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_254),
.A2(n_557),
.B(n_560),
.Y(n_556)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_255),
.B(n_256),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_283),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g563 ( 
.A(n_258),
.B(n_259),
.C(n_283),
.Y(n_563)
);

XNOR2x1_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_269),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_266),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_261),
.B(n_266),
.C(n_269),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_267),
.B(n_272),
.C(n_278),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_278),
.B1(n_279),
.B2(n_282),
.Y(n_269)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_271),
.A2(n_272),
.B1(n_572),
.B2(n_573),
.Y(n_571)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI21x1_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_395),
.B(n_553),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_347),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_287),
.A2(n_554),
.B(n_555),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_344),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g555 ( 
.A(n_288),
.B(n_344),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.C(n_342),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_290),
.B(n_342),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_293),
.B(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_317),
.C(n_335),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_294),
.B(n_351),
.Y(n_350)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_299),
.C(n_311),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_296),
.B(n_298),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_299),
.A2(n_300),
.B1(n_311),
.B2(n_312),
.Y(n_422)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_304),
.B(n_307),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_362),
.Y(n_361)
);

AOI21xp33_ASAP7_75t_SL g307 ( 
.A1(n_302),
.A2(n_308),
.B(n_310),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_304),
.A2(n_305),
.B1(n_310),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_309),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

OA21x2_ASAP7_75t_SL g406 ( 
.A1(n_312),
.A2(n_313),
.B(n_316),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_318),
.A2(n_336),
.B1(n_337),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_318),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_328),
.C(n_332),
.Y(n_318)
);

XOR2x1_ASAP7_75t_L g391 ( 
.A(n_319),
.B(n_392),
.Y(n_391)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_325),
.C(n_327),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_320),
.A2(n_321),
.B1(n_327),
.B2(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_323),
.Y(n_477)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_325),
.B(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_328),
.A2(n_329),
.B1(n_332),
.B2(n_333),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_337)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_339),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_393),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_348),
.B(n_393),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_353),
.C(n_358),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_350),
.B(n_354),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_358),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_386),
.C(n_389),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_359),
.A2(n_360),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.C(n_375),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_361),
.B(n_445),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_364),
.A2(n_375),
.B1(n_376),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_364),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_370),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_365),
.A2(n_366),
.B1(n_370),
.B2(n_371),
.Y(n_442)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_374),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_374),
.Y(n_534)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

MAJx2_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_381),
.C(n_382),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_377),
.A2(n_378),
.B1(n_382),
.B2(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_381),
.B(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_382),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_385),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_386),
.A2(n_390),
.B1(n_391),
.B2(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_386),
.Y(n_401)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_449),
.B(n_551),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_423),
.B(n_426),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_397),
.B(n_423),
.C(n_552),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_402),
.C(n_419),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_398),
.B(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_402),
.B(n_420),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_406),
.C(n_407),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_406),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_407),
.B(n_429),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_413),
.C(n_415),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_408),
.B(n_465),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_409),
.A2(n_410),
.B1(n_411),
.B2(n_412),
.Y(n_455)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_413),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_465)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_418),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_447),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_427),
.B(n_447),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_430),
.C(n_443),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_428),
.B(n_467),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_430),
.B(n_444),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_434),
.C(n_442),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_453),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_442),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.C(n_439),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_435),
.B(n_439),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_436),
.B(n_500),
.Y(n_499)
);

INVx3_ASAP7_75t_SL g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_441),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_468),
.B(n_550),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_466),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_SL g550 ( 
.A(n_451),
.B(n_466),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_454),
.C(n_464),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_452),
.B(n_548),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_454),
.B(n_464),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.C(n_457),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_455),
.B(n_456),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_457),
.B(n_494),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_461),
.Y(n_457)
);

AO22x1_ASAP7_75t_L g490 ( 
.A1(n_458),
.A2(n_459),
.B1(n_461),
.B2(n_462),
.Y(n_490)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_469),
.A2(n_545),
.B(n_549),
.Y(n_468)
);

OAI21x1_ASAP7_75t_SL g469 ( 
.A1(n_470),
.A2(n_502),
.B(n_544),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_491),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_471),
.B(n_491),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_484),
.C(n_490),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_472),
.A2(n_473),
.B1(n_540),
.B2(n_542),
.Y(n_539)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_474),
.B(n_478),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_497),
.C(n_498),
.Y(n_496)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_482),
.Y(n_478)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_479),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_482),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_484),
.A2(n_485),
.B1(n_490),
.B2(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_489),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_486),
.B(n_489),
.Y(n_520)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_490),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_492),
.A2(n_493),
.B1(n_495),
.B2(n_501),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_492),
.B(n_496),
.C(n_499),
.Y(n_546)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_495),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_499),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_537),
.B(n_543),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_504),
.A2(n_521),
.B(n_536),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_513),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_505),
.B(n_513),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_506),
.B(n_510),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_506),
.B(n_510),
.Y(n_529)
);

INVx4_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx8_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_510),
.B(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_520),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_515),
.A2(n_516),
.B1(n_517),
.B2(n_519),
.Y(n_514)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_515),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_516),
.B(n_519),
.C(n_520),
.Y(n_538)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_522),
.A2(n_530),
.B(n_535),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_529),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_529),
.Y(n_535)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx3_ASAP7_75t_SL g532 ( 
.A(n_533),
.Y(n_532)
);

INVx8_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_539),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_538),
.B(n_539),
.Y(n_543)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_540),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_SL g545 ( 
.A(n_546),
.B(n_547),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_546),
.B(n_547),
.Y(n_549)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_561),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_562),
.B(n_577),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_564),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_563),
.B(n_564),
.Y(n_577)
);

BUFx24_ASAP7_75t_SL g580 ( 
.A(n_564),
.Y(n_580)
);

FAx1_ASAP7_75t_SL g564 ( 
.A(n_565),
.B(n_566),
.CI(n_567),
.CON(n_564),
.SN(n_564)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_571),
.Y(n_567)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_574),
.B(n_576),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);


endmodule