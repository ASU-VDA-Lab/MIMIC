module fake_jpeg_7477_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_14),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_16),
.B(n_19),
.Y(n_24)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_21),
.Y(n_23)
);

CKINVDCx9p33_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_0),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_14),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_36),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_22),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_10),
.B1(n_17),
.B2(n_21),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_16),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_15),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_17),
.C(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_42),
.B1(n_43),
.B2(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_35),
.B1(n_21),
.B2(n_17),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_44),
.C(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_39),
.B(n_45),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_51),
.C(n_50),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_54),
.A2(n_55),
.B(n_28),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_46),
.C(n_32),
.Y(n_55)
);

BUFx24_ASAP7_75t_SL g57 ( 
.A(n_56),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_8),
.Y(n_59)
);


endmodule