module fake_jpeg_2548_n_154 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_55),
.Y(n_65)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_70),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_51),
.B1(n_55),
.B2(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_44),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_54),
.C(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_79),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_42),
.B(n_47),
.C(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_82),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_62),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_86),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_48),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_87),
.B(n_0),
.Y(n_103)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_41),
.B(n_43),
.C(n_49),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_66),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_89),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_41),
.C(n_50),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_88),
.B1(n_81),
.B2(n_79),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_71),
.B1(n_48),
.B2(n_50),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_71),
.B1(n_46),
.B2(n_60),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_46),
.B1(n_1),
.B2(n_2),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_18),
.C(n_39),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_105),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_96),
.B(n_97),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_40),
.B1(n_23),
.B2(n_24),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_5),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_107),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_31),
.B(n_36),
.C(n_34),
.D(n_33),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_119),
.B(n_9),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_6),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_7),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_7),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_8),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_8),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_37),
.B(n_30),
.C(n_29),
.Y(n_122)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_28),
.B(n_26),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_129),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_9),
.C(n_11),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_117),
.C(n_113),
.Y(n_140)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_11),
.B(n_12),
.C(n_13),
.D(n_14),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_134),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_128),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_121),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_121),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_113),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_143),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_140),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_131),
.B(n_122),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_139),
.B(n_108),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_138),
.B(n_126),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_145),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_145),
.B1(n_124),
.B2(n_133),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_141),
.B(n_132),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_141),
.B(n_125),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_119),
.Y(n_154)
);


endmodule