module fake_jpeg_15060_n_149 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_149);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_31),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_13),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_46),
.B(n_48),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_13),
.C(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_49),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_21),
.B1(n_22),
.B2(n_13),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_26),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_21),
.B1(n_24),
.B2(n_17),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_19),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_36),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_32),
.B1(n_25),
.B2(n_34),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_45),
.B1(n_31),
.B2(n_39),
.Y(n_70)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_14),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_14),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_63),
.B1(n_29),
.B2(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_25),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_57),
.B1(n_54),
.B2(n_60),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_80),
.B1(n_69),
.B2(n_71),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_54),
.B1(n_60),
.B2(n_29),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_42),
.B(n_30),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_64),
.B(n_75),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_47),
.B(n_58),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_30),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_44),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_66),
.B1(n_77),
.B2(n_71),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_30),
.C(n_27),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_27),
.C(n_30),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_96),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_104),
.B1(n_83),
.B2(n_84),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_66),
.B1(n_44),
.B2(n_17),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_50),
.B1(n_80),
.B2(n_20),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_8),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_105),
.Y(n_116)
);

AO21x2_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_92),
.B(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_7),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_89),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_112),
.B(n_42),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_104),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_79),
.B(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

OAI322xp33_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_104),
.A3(n_98),
.B1(n_93),
.B2(n_96),
.C1(n_97),
.C2(n_95),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_119),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_94),
.B1(n_50),
.B2(n_2),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_124),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_115),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_129),
.C(n_130),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_107),
.C(n_109),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_108),
.C(n_42),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_20),
.C(n_23),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_137),
.Y(n_140)
);

AOI31xp67_ASAP7_75t_SL g134 ( 
.A1(n_131),
.A2(n_125),
.A3(n_128),
.B(n_121),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_5),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_4),
.B(n_12),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_135),
.A2(n_4),
.B(n_12),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_138),
.A2(n_11),
.B(n_1),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_0),
.C(n_2),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_144),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_0),
.B(n_1),
.Y(n_143)
);

NOR2x1_ASAP7_75t_SL g145 ( 
.A(n_143),
.B(n_3),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_145),
.A2(n_23),
.B(n_140),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_146),
.B(n_23),
.Y(n_148)
);

XNOR2x2_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_23),
.Y(n_149)
);


endmodule