module fake_jpeg_13001_n_567 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_567);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_567;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_55),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_23),
.B(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_59),
.Y(n_108)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_25),
.B(n_9),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_66),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_70),
.Y(n_170)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_78),
.Y(n_156)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_23),
.B(n_10),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_85),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_51),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_35),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_89),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_99),
.Y(n_126)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_26),
.B(n_10),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_96),
.B(n_103),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_26),
.B(n_18),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_12),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_31),
.B(n_8),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_20),
.B1(n_46),
.B2(n_32),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_111),
.A2(n_140),
.B1(n_141),
.B2(n_144),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_114),
.B(n_115),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_51),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_51),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_119),
.B(n_152),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_60),
.A2(n_19),
.B1(n_46),
.B2(n_20),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_123),
.A2(n_142),
.B1(n_33),
.B2(n_42),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_50),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_149),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_73),
.A2(n_19),
.B1(n_46),
.B2(n_32),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_79),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_64),
.A2(n_32),
.B1(n_22),
.B2(n_24),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_91),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_89),
.B(n_50),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_50),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_67),
.A2(n_49),
.B1(n_48),
.B2(n_43),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_158),
.A2(n_48),
.B1(n_31),
.B2(n_43),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_69),
.B(n_49),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_42),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_93),
.Y(n_168)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_171),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_66),
.B(n_21),
.C(n_29),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_172),
.B(n_179),
.Y(n_273)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

BUFx2_ASAP7_75t_SL g244 ( 
.A(n_173),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_42),
.B(n_33),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_205),
.C(n_31),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_175),
.A2(n_207),
.B1(n_30),
.B2(n_27),
.Y(n_245)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_176),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_177),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_126),
.Y(n_179)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_182),
.Y(n_270)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_187),
.B(n_188),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_108),
.B(n_86),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_113),
.B(n_37),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_189),
.B(n_195),
.Y(n_239)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_190),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

INVx4_ASAP7_75t_SL g192 ( 
.A(n_151),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_192),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_126),
.A2(n_29),
.B(n_30),
.C(n_27),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g284 ( 
.A1(n_193),
.A2(n_228),
.B(n_229),
.Y(n_284)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_138),
.B(n_43),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

INVx3_ASAP7_75t_SL g260 ( 
.A(n_196),
.Y(n_260)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_197),
.Y(n_250)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_199),
.Y(n_280)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_201),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_118),
.B(n_37),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_202),
.B(n_219),
.Y(n_265)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_203),
.Y(n_281)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_204),
.B(n_206),
.Y(n_251)
);

NAND2x1_ASAP7_75t_L g205 ( 
.A(n_139),
.B(n_153),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_120),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_123),
.A2(n_70),
.B1(n_72),
.B2(n_80),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_142),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_208),
.B(n_209),
.Y(n_255)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_210),
.B(n_212),
.Y(n_264)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_137),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_211),
.Y(n_254)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_125),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_213),
.Y(n_288)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_147),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_122),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_215),
.B(n_218),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_110),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_217),
.Y(n_277)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_129),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_128),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_139),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_220),
.Y(n_241)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_133),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_221),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_156),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_222),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_132),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_223),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_110),
.A2(n_55),
.B1(n_87),
.B2(n_92),
.Y(n_224)
);

OAI22x1_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_141),
.B1(n_140),
.B2(n_144),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_117),
.B(n_37),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_225),
.B(n_232),
.Y(n_267)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_132),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_226),
.B(n_227),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_161),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_155),
.Y(n_228)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_156),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_230),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_278)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_146),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_233),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_111),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_134),
.B1(n_135),
.B2(n_159),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_234),
.A2(n_245),
.B1(n_259),
.B2(n_222),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_236),
.A2(n_7),
.B1(n_15),
.B2(n_4),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_246),
.A2(n_8),
.B(n_17),
.C(n_15),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_185),
.B(n_178),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_257),
.B(n_271),
.C(n_275),
.Y(n_304)
);

AOI32xp33_ASAP7_75t_L g258 ( 
.A1(n_179),
.A2(n_148),
.A3(n_98),
.B1(n_49),
.B2(n_48),
.Y(n_258)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_258),
.B(n_14),
.CI(n_15),
.CON(n_331),
.SN(n_331)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_174),
.A2(n_160),
.B1(n_127),
.B2(n_154),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_193),
.B(n_230),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_272),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_216),
.A2(n_84),
.B1(n_127),
.B2(n_154),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_278),
.B1(n_287),
.B2(n_172),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_205),
.B(n_148),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_180),
.B(n_216),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_97),
.C(n_90),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_226),
.B(n_135),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_283),
.B(n_184),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_181),
.B(n_30),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_192),
.C(n_191),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_224),
.A2(n_160),
.B1(n_166),
.B2(n_170),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_289),
.A2(n_291),
.B1(n_293),
.B2(n_295),
.Y(n_341)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_290),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_211),
.B1(n_213),
.B2(n_134),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_182),
.B(n_227),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_292),
.A2(n_280),
.B(n_237),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_262),
.A2(n_166),
.B1(n_170),
.B2(n_173),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_294),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_267),
.A2(n_287),
.B1(n_273),
.B2(n_236),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_267),
.A2(n_171),
.B1(n_196),
.B2(n_176),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_296),
.A2(n_298),
.B1(n_299),
.B2(n_301),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_273),
.A2(n_220),
.B(n_217),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_297),
.A2(n_280),
.B(n_237),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_245),
.A2(n_190),
.B1(n_214),
.B2(n_101),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_305),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_259),
.A2(n_255),
.B1(n_235),
.B2(n_265),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_252),
.Y(n_302)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_252),
.Y(n_303)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_303),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_273),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_194),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_306),
.B(n_327),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_307),
.B(n_264),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_308),
.B(n_309),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_239),
.A2(n_102),
.B1(n_199),
.B2(n_229),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_246),
.A2(n_199),
.B1(n_1),
.B2(n_2),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_310),
.B(n_313),
.Y(n_359)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_268),
.Y(n_312)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_312),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_258),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g314 ( 
.A(n_257),
.B(n_271),
.C(n_284),
.Y(n_314)
);

XNOR2x1_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_325),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_238),
.A2(n_8),
.B1(n_17),
.B2(n_16),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_315),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_316),
.A2(n_321),
.B(n_324),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_275),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_317),
.B(n_323),
.Y(n_362)
);

O2A1O1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_251),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_318)
);

O2A1O1Ixp33_ASAP7_75t_L g357 ( 
.A1(n_318),
.A2(n_247),
.B(n_281),
.C(n_249),
.Y(n_357)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_283),
.A2(n_11),
.B(n_15),
.Y(n_319)
);

OAI21xp33_ASAP7_75t_L g349 ( 
.A1(n_319),
.A2(n_331),
.B(n_256),
.Y(n_349)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_320),
.Y(n_380)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_270),
.Y(n_322)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_322),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_276),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_323)
);

AO22x1_ASAP7_75t_L g324 ( 
.A1(n_278),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_250),
.B(n_243),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_238),
.A2(n_5),
.B1(n_12),
.B2(n_13),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_326),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_250),
.B(n_5),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_269),
.B(n_12),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_328),
.B(n_281),
.Y(n_363)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_268),
.Y(n_329)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_329),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_243),
.B(n_13),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_330),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_242),
.A2(n_14),
.B1(n_18),
.B2(n_286),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_242),
.A2(n_14),
.B1(n_286),
.B2(n_266),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_266),
.A2(n_240),
.B1(n_241),
.B2(n_248),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_248),
.Y(n_335)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_276),
.A2(n_260),
.B1(n_240),
.B2(n_241),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_336),
.A2(n_260),
.B1(n_253),
.B2(n_279),
.Y(n_368)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_274),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_337),
.B(n_274),
.Y(n_360)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_279),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_338),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_339),
.A2(n_351),
.B(n_371),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_342),
.B(n_309),
.C(n_317),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_334),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_345),
.B(n_350),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_349),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_311),
.Y(n_350)
);

OA21x2_ASAP7_75t_L g351 ( 
.A1(n_311),
.A2(n_282),
.B(n_288),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_295),
.A2(n_260),
.B1(n_254),
.B2(n_288),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_352),
.A2(n_368),
.B1(n_369),
.B2(n_299),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_354),
.A2(n_318),
.B(n_323),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_357),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_360),
.B(n_364),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_290),
.B(n_294),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_361),
.B(n_363),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_333),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_289),
.A2(n_274),
.B1(n_253),
.B2(n_247),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_292),
.A2(n_300),
.B(n_297),
.Y(n_371)
);

OAI32xp33_ASAP7_75t_L g372 ( 
.A1(n_325),
.A2(n_249),
.A3(n_244),
.B1(n_256),
.B2(n_277),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_374),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_301),
.B(n_277),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_336),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_377),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_332),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_307),
.B(n_321),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_378),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_361),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_382),
.B(n_390),
.Y(n_431)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_380),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_383),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_375),
.A2(n_304),
.B1(n_291),
.B2(n_331),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_385),
.A2(n_394),
.B1(n_397),
.B2(n_378),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_347),
.B(n_304),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_386),
.B(n_388),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_347),
.B(n_314),
.Y(n_388)
);

NAND2xp33_ASAP7_75t_SL g421 ( 
.A(n_389),
.B(n_354),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_368),
.Y(n_390)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_391),
.Y(n_426)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_344),
.Y(n_392)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_392),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_341),
.A2(n_369),
.B1(n_350),
.B2(n_345),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_393),
.A2(n_398),
.B1(n_399),
.B2(n_409),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_365),
.A2(n_331),
.B1(n_293),
.B2(n_310),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_360),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_396),
.B(n_402),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_365),
.A2(n_316),
.B1(n_313),
.B2(n_302),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_341),
.A2(n_351),
.B1(n_352),
.B2(n_340),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_351),
.A2(n_340),
.B1(n_343),
.B2(n_377),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_376),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_343),
.B(n_303),
.Y(n_404)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_404),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_351),
.B(n_338),
.Y(n_405)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_405),
.Y(n_447)
);

OAI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_357),
.A2(n_316),
.B1(n_296),
.B2(n_324),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_406),
.A2(n_367),
.B1(n_370),
.B2(n_324),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_376),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_353),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_371),
.A2(n_316),
.B(n_335),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_408),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_359),
.A2(n_364),
.B1(n_346),
.B2(n_358),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_376),
.B(n_330),
.Y(n_411)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_411),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_418),
.Y(n_428)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_380),
.Y(n_414)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_414),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_347),
.B(n_298),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_355),
.Y(n_444)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_417),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_342),
.B(n_379),
.C(n_348),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_404),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_419),
.B(n_421),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_393),
.A2(n_359),
.B1(n_374),
.B2(n_358),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_425),
.A2(n_443),
.B1(n_437),
.B2(n_422),
.Y(n_469)
);

CKINVDCx14_ASAP7_75t_R g427 ( 
.A(n_403),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_433),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_386),
.B(n_348),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_429),
.B(n_430),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_339),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_412),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_434),
.A2(n_442),
.B1(n_445),
.B2(n_450),
.Y(n_455)
);

OAI21xp33_ASAP7_75t_L g435 ( 
.A1(n_382),
.A2(n_357),
.B(n_356),
.Y(n_435)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_435),
.Y(n_463)
);

OA21x2_ASAP7_75t_L g437 ( 
.A1(n_405),
.A2(n_372),
.B(n_362),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_437),
.B(n_441),
.Y(n_471)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_439),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_403),
.B(n_363),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_390),
.A2(n_346),
.B1(n_362),
.B2(n_373),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_398),
.A2(n_373),
.B1(n_355),
.B2(n_376),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_389),
.Y(n_473)
);

FAx1_ASAP7_75t_SL g445 ( 
.A(n_388),
.B(n_356),
.CI(n_316),
.CON(n_445),
.SN(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_413),
.B(n_320),
.Y(n_446)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_394),
.A2(n_353),
.B1(n_367),
.B2(n_366),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_451),
.A2(n_391),
.B1(n_412),
.B2(n_384),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_410),
.C(n_411),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_453),
.C(n_454),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_410),
.C(n_415),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_385),
.C(n_400),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_387),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_461),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_426),
.A2(n_395),
.B1(n_397),
.B2(n_416),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_457),
.A2(n_458),
.B1(n_464),
.B2(n_469),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_426),
.A2(n_395),
.B1(n_416),
.B2(n_408),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_420),
.B(n_400),
.C(n_401),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_459),
.B(n_462),
.C(n_468),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_424),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_420),
.B(n_387),
.C(n_399),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_422),
.A2(n_384),
.B1(n_396),
.B2(n_409),
.Y(n_464)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_467),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_407),
.C(n_402),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_473),
.B(n_479),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_432),
.B(n_417),
.C(n_392),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_452),
.C(n_453),
.Y(n_502)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_436),
.Y(n_475)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_475),
.Y(n_491)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_436),
.Y(n_476)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_476),
.Y(n_497)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_432),
.Y(n_477)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_477),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_431),
.B(n_366),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_423),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_431),
.B(n_381),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_466),
.B(n_447),
.Y(n_480)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_480),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_471),
.A2(n_450),
.B1(n_442),
.B2(n_447),
.Y(n_481)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_481),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_457),
.A2(n_451),
.B1(n_449),
.B2(n_448),
.Y(n_484)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_484),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_478),
.B(n_474),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_485),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_463),
.A2(n_449),
.B(n_437),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_486),
.A2(n_456),
.B(n_459),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_460),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_489),
.B(n_492),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_464),
.A2(n_425),
.B1(n_443),
.B2(n_445),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_493),
.B(n_470),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_455),
.A2(n_445),
.B(n_440),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_494),
.A2(n_473),
.B(n_454),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_465),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_495),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_458),
.A2(n_440),
.B1(n_438),
.B2(n_414),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_501),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_462),
.A2(n_383),
.B1(n_381),
.B2(n_370),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_502),
.Y(n_505)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_468),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_506),
.A2(n_492),
.B(n_511),
.Y(n_533)
);

INVx4_ASAP7_75t_L g507 ( 
.A(n_495),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_507),
.B(n_511),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_518),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_470),
.C(n_461),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_512),
.B(n_487),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_472),
.C(n_322),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_515),
.B(n_516),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_329),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_312),
.C(n_337),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_517),
.B(n_501),
.C(n_485),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_487),
.B(n_483),
.Y(n_518)
);

BUFx24_ASAP7_75t_SL g520 ( 
.A(n_486),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_521),
.Y(n_525)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_480),
.B(n_498),
.C(n_491),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_522),
.B(n_523),
.Y(n_547)
);

AOI21x1_ASAP7_75t_L g524 ( 
.A1(n_503),
.A2(n_494),
.B(n_488),
.Y(n_524)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_524),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_505),
.B(n_482),
.C(n_488),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_526),
.B(n_527),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_505),
.B(n_483),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_491),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_528),
.B(n_529),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_519),
.A2(n_497),
.B1(n_498),
.B2(n_490),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_515),
.A2(n_482),
.B(n_497),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_530),
.B(n_533),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_517),
.B(n_490),
.C(n_493),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_531),
.B(n_509),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_504),
.B(n_514),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_534),
.B(n_525),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_537),
.B(n_538),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_513),
.Y(n_538)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_528),
.Y(n_540)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_540),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_532),
.B(n_509),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_544),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_523),
.B(n_527),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_545),
.B(n_531),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_540),
.A2(n_533),
.B(n_508),
.Y(n_548)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_548),
.Y(n_558)
);

INVx11_ASAP7_75t_L g551 ( 
.A(n_541),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_551),
.B(n_552),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_543),
.A2(n_535),
.B(n_507),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_554),
.B(n_547),
.C(n_549),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_555),
.B(n_556),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_553),
.B(n_539),
.C(n_547),
.Y(n_556)
);

BUFx24_ASAP7_75t_SL g559 ( 
.A(n_558),
.Y(n_559)
);

AO21x1_ASAP7_75t_L g563 ( 
.A1(n_559),
.A2(n_546),
.B(n_536),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_557),
.A2(n_548),
.B(n_551),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_560),
.A2(n_550),
.B(n_552),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_562),
.A2(n_563),
.B(n_561),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_564),
.A2(n_546),
.B(n_535),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_565),
.B(n_522),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_566),
.A2(n_518),
.B(n_512),
.Y(n_567)
);


endmodule