module fake_jpeg_21647_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_18),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_26)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_10),
.B(n_15),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_0),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_13),
.C(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_30),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_7),
.B1(n_14),
.B2(n_2),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_23),
.B1(n_14),
.B2(n_18),
.Y(n_33)
);

AND2x6_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_15),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_27),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_29),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_21),
.B1(n_17),
.B2(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_39),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_26),
.B(n_28),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_31),
.B1(n_35),
.B2(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_25),
.Y(n_45)
);

AO21x1_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_40),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_42),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_47),
.A2(n_48),
.B(n_40),
.Y(n_49)
);

AOI322xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.A3(n_0),
.B1(n_1),
.B2(n_2),
.C1(n_3),
.C2(n_5),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);


endmodule