module fake_jpeg_28570_n_469 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_469);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_469;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx8_ASAP7_75t_SL g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_50),
.B(n_73),
.Y(n_110)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_56),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_31),
.A2(n_16),
.B(n_15),
.C(n_14),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_66),
.A2(n_39),
.B(n_36),
.C(n_25),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

CKINVDCx6p67_ASAP7_75t_R g151 ( 
.A(n_71),
.Y(n_151)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_37),
.B(n_39),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_101),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_19),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_116),
.B(n_136),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_50),
.B(n_21),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_142),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_20),
.B1(n_30),
.B2(n_34),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_160),
.B1(n_75),
.B2(n_86),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_69),
.B(n_32),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_55),
.B(n_21),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_56),
.B(n_32),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_153),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_71),
.B(n_44),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_57),
.B(n_44),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_158),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_71),
.B(n_22),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_64),
.A2(n_30),
.B1(n_34),
.B2(n_20),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_126),
.A2(n_23),
.B1(n_45),
.B2(n_40),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_161),
.A2(n_210),
.B1(n_211),
.B2(n_122),
.Y(n_234)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g249 ( 
.A(n_163),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_164),
.B(n_168),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_110),
.B(n_46),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_165),
.B(n_167),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g223 ( 
.A(n_166),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_110),
.B(n_74),
.C(n_98),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_158),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_132),
.B(n_36),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_169),
.B(n_203),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_172),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_151),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_171),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_151),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_173),
.B(n_175),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_115),
.B(n_101),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_180),
.A2(n_194),
.B1(n_198),
.B2(n_114),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_181),
.B(n_183),
.Y(n_247)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_118),
.B(n_101),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_81),
.B1(n_76),
.B2(n_84),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_185),
.A2(n_204),
.B1(n_135),
.B2(n_155),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_143),
.A2(n_23),
.B1(n_25),
.B2(n_42),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_199),
.Y(n_229)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_105),
.B(n_17),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_193),
.Y(n_213)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_107),
.B(n_17),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_108),
.A2(n_94),
.B1(n_92),
.B2(n_91),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_120),
.B(n_26),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_42),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_128),
.A2(n_95),
.B1(n_85),
.B2(n_34),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_121),
.A2(n_23),
.B1(n_26),
.B2(n_22),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_145),
.Y(n_201)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_104),
.B(n_87),
.Y(n_203)
);

AO22x1_ASAP7_75t_SL g204 ( 
.A1(n_124),
.A2(n_30),
.B1(n_34),
.B2(n_45),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_111),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_208),
.B(n_209),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_154),
.Y(n_209)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

INVx3_ASAP7_75t_SL g211 ( 
.A(n_137),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_220),
.A2(n_241),
.B1(n_242),
.B2(n_170),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_227),
.B(n_232),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_165),
.B(n_46),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_176),
.C(n_186),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_191),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_234),
.A2(n_208),
.B(n_206),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_177),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_235),
.B(n_181),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_238),
.A2(n_250),
.B1(n_251),
.B2(n_197),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_166),
.A2(n_133),
.B1(n_147),
.B2(n_159),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_189),
.A2(n_150),
.B1(n_129),
.B2(n_131),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_207),
.A2(n_148),
.B1(n_134),
.B2(n_127),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_211),
.A2(n_139),
.B1(n_130),
.B2(n_141),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_238),
.A2(n_184),
.B1(n_167),
.B2(n_178),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_253),
.A2(n_257),
.B1(n_269),
.B2(n_273),
.Y(n_312)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_248),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_267),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_256),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_213),
.A2(n_178),
.B1(n_193),
.B2(n_196),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_258),
.A2(n_265),
.B1(n_270),
.B2(n_283),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_259),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_87),
.Y(n_304)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_261),
.Y(n_298)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_263),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_212),
.B(n_231),
.C(n_232),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_244),
.C(n_214),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_223),
.A2(n_114),
.B1(n_201),
.B2(n_199),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_266),
.A2(n_280),
.B1(n_282),
.B2(n_236),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_229),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_213),
.A2(n_176),
.B1(n_204),
.B2(n_192),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_223),
.A2(n_204),
.B1(n_179),
.B2(n_163),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_173),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_272),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_229),
.A2(n_200),
.B1(n_187),
.B2(n_202),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_216),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_275),
.Y(n_297)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_276),
.Y(n_307)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_243),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_279),
.A2(n_281),
.B1(n_218),
.B2(n_244),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_227),
.A2(n_149),
.B1(n_205),
.B2(n_174),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_219),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_220),
.A2(n_210),
.B1(n_182),
.B2(n_190),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_229),
.A2(n_195),
.B1(n_40),
.B2(n_13),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_218),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_221),
.B(n_239),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_260),
.A2(n_215),
.B(n_212),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_286),
.A2(n_303),
.B(n_306),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_242),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_289),
.B(n_290),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_217),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_292),
.A2(n_283),
.B1(n_261),
.B2(n_254),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_293),
.Y(n_326)
);

OA21x2_ASAP7_75t_L g294 ( 
.A1(n_258),
.A2(n_247),
.B(n_224),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_294),
.B(n_281),
.Y(n_335)
);

OAI32xp33_ASAP7_75t_L g299 ( 
.A1(n_269),
.A2(n_230),
.A3(n_219),
.B1(n_228),
.B2(n_221),
.Y(n_299)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_299),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_285),
.A2(n_249),
.B(n_226),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_304),
.B(n_276),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_255),
.A2(n_228),
.B(n_226),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_309),
.A2(n_293),
.B(n_294),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_257),
.Y(n_323)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_316),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_295),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_317),
.B(n_332),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_315),
.A2(n_275),
.B1(n_282),
.B2(n_259),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_320),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_322),
.B(n_335),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_323),
.B(n_289),
.C(n_304),
.Y(n_366)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_300),
.A2(n_280),
.B1(n_285),
.B2(n_277),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_325),
.A2(n_330),
.B1(n_339),
.B2(n_298),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_327),
.A2(n_328),
.B1(n_344),
.B2(n_302),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_287),
.A2(n_268),
.B1(n_274),
.B2(n_262),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_309),
.Y(n_329)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_329),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_300),
.A2(n_284),
.B1(n_252),
.B2(n_263),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_288),
.Y(n_331)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_331),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_295),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_297),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_341),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_338),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_315),
.A2(n_279),
.B(n_278),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_288),
.Y(n_364)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_337),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_214),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_294),
.A2(n_249),
.B1(n_268),
.B2(n_271),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_340),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_312),
.B(n_237),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_292),
.A2(n_271),
.B1(n_237),
.B2(n_12),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_342),
.A2(n_298),
.B1(n_302),
.B2(n_305),
.Y(n_365)
);

BUFx12f_ASAP7_75t_L g343 ( 
.A(n_298),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_343),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_312),
.A2(n_33),
.B1(n_47),
.B2(n_43),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_349),
.A2(n_318),
.B1(n_326),
.B2(n_339),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_343),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_351),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_331),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_343),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_355),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_335),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_338),
.B(n_321),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_358),
.B(n_359),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_313),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_322),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_361),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_337),
.Y(n_362)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_362),
.Y(n_373)
);

OAI21xp33_ASAP7_75t_L g388 ( 
.A1(n_364),
.A2(n_296),
.B(n_311),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_365),
.A2(n_368),
.B1(n_330),
.B2(n_318),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_370),
.C(n_319),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_323),
.B(n_290),
.C(n_303),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_334),
.B(n_314),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_371),
.B(n_319),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_374),
.A2(n_378),
.B1(n_381),
.B2(n_391),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_375),
.A2(n_345),
.B1(n_363),
.B2(n_4),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_379),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_349),
.A2(n_344),
.B1(n_326),
.B2(n_299),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_357),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_393),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_348),
.A2(n_325),
.B1(n_305),
.B2(n_307),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_336),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_383),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_320),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_301),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_385),
.B(n_386),
.C(n_389),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_307),
.C(n_296),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_367),
.Y(n_387)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_387),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_390),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_311),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_291),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_348),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_361),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_SL g393 ( 
.A(n_371),
.B(n_0),
.C(n_3),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_347),
.Y(n_407)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_395),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_384),
.A2(n_368),
.B1(n_352),
.B2(n_364),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_402),
.A2(n_406),
.B1(n_377),
.B2(n_3),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_352),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_403),
.B(n_47),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_386),
.B(n_357),
.C(n_356),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_405),
.C(n_47),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_382),
.C(n_372),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_376),
.A2(n_365),
.B1(n_346),
.B2(n_354),
.Y(n_406)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_407),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_373),
.B(n_347),
.Y(n_408)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_408),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_363),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_409),
.B(n_410),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g410 ( 
.A(n_383),
.B(n_345),
.CI(n_356),
.CON(n_410),
.SN(n_410)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_0),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_390),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_416),
.Y(n_436)
);

BUFx24_ASAP7_75t_SL g415 ( 
.A(n_400),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_415),
.B(n_397),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_395),
.A2(n_379),
.B(n_388),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_417),
.B(n_421),
.Y(n_428)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_420),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_422),
.B(n_403),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_47),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_423),
.B(n_424),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_401),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_47),
.C(n_43),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_412),
.C(n_399),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_427),
.B(n_431),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_426),
.B(n_396),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_430),
.B(n_47),
.C(n_43),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_413),
.A2(n_411),
.B1(n_402),
.B2(n_410),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_432),
.A2(n_0),
.B1(n_5),
.B2(n_8),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_419),
.A2(n_405),
.B(n_396),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_434),
.A2(n_422),
.B(n_412),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_435),
.B(n_437),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_425),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_438),
.Y(n_447)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_420),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_439),
.Y(n_441)
);

AOI21x1_ASAP7_75t_L g442 ( 
.A1(n_436),
.A2(n_410),
.B(n_399),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_444),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_448),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_432),
.A2(n_421),
.B(n_4),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_435),
.C(n_437),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_43),
.C(n_5),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_446),
.B(n_433),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_449),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_451),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_447),
.B(n_440),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_454),
.B(n_455),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_427),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_456),
.B(n_446),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_451),
.B(n_453),
.C(n_452),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_457),
.B(n_458),
.C(n_428),
.Y(n_463)
);

NOR3xp33_ASAP7_75t_L g461 ( 
.A(n_459),
.B(n_445),
.C(n_444),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_461),
.B(n_462),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_460),
.A2(n_429),
.B(n_428),
.Y(n_462)
);

A2O1A1O1Ixp25_ASAP7_75t_L g465 ( 
.A1(n_463),
.A2(n_5),
.B(n_9),
.C(n_10),
.D(n_11),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_465),
.A2(n_9),
.B(n_11),
.Y(n_466)
);

MAJx2_ASAP7_75t_L g467 ( 
.A(n_466),
.B(n_464),
.C(n_11),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_11),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_43),
.Y(n_469)
);


endmodule