module fake_jpeg_27984_n_236 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_5),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_32),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_18),
.B1(n_21),
.B2(n_20),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_46),
.B1(n_39),
.B2(n_35),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_22),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_15),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_37),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_43),
.B1(n_18),
.B2(n_40),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_69),
.B1(n_70),
.B2(n_46),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_34),
.B(n_37),
.C(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

AOI32xp33_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_34),
.A3(n_21),
.B1(n_27),
.B2(n_30),
.Y(n_62)
);

MAJx2_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_50),
.C(n_47),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_39),
.B1(n_42),
.B2(n_31),
.Y(n_70)
);

NOR2x1_ASAP7_75t_R g71 ( 
.A(n_55),
.B(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_27),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_74),
.B1(n_68),
.B2(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_48),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_87),
.B1(n_72),
.B2(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_45),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_58),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_75),
.B1(n_89),
.B2(n_86),
.Y(n_93)
);

BUFx4f_ASAP7_75t_SL g83 ( 
.A(n_59),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_88),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_95),
.B1(n_105),
.B2(n_108),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_88),
.B1(n_86),
.B2(n_85),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_94),
.A2(n_31),
.B1(n_47),
.B2(n_49),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_61),
.B1(n_73),
.B2(n_71),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_63),
.C(n_71),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_100),
.C(n_109),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_63),
.A3(n_70),
.B1(n_62),
.B2(n_66),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_63),
.C(n_66),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_59),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_80),
.B1(n_87),
.B2(n_76),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_54),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_78),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_72),
.B1(n_57),
.B2(n_53),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_57),
.B1(n_56),
.B2(n_67),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_33),
.C(n_24),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_107),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_112),
.Y(n_151)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_29),
.B1(n_13),
.B2(n_14),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_64),
.B1(n_46),
.B2(n_83),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_120),
.A2(n_121),
.B1(n_126),
.B2(n_130),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_64),
.B1(n_83),
.B2(n_26),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_83),
.B(n_1),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_19),
.B(n_1),
.Y(n_147)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_29),
.B1(n_24),
.B2(n_12),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_15),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_121),
.B(n_120),
.C(n_116),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_104),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_17),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_47),
.B1(n_49),
.B2(n_22),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_99),
.B1(n_19),
.B2(n_49),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_25),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_135),
.Y(n_163)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_128),
.B(n_118),
.CI(n_97),
.CON(n_135),
.SN(n_135)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_98),
.B1(n_106),
.B2(n_104),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_136),
.A2(n_143),
.B1(n_147),
.B2(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_117),
.B(n_5),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_113),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_119),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_49),
.B1(n_11),
.B2(n_14),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_49),
.B1(n_11),
.B2(n_14),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_112),
.B1(n_119),
.B2(n_16),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_155),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_137),
.B(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_126),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_128),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_170),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_131),
.C(n_133),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_171),
.C(n_146),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_135),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_125),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_169),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_9),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_17),
.C(n_13),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_14),
.B1(n_11),
.B2(n_16),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_150),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_175),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_136),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_162),
.B1(n_145),
.B2(n_138),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_177),
.A2(n_182),
.B1(n_147),
.B2(n_136),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_153),
.C(n_146),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_13),
.C(n_17),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_184),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_138),
.B1(n_148),
.B2(n_146),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_157),
.B1(n_16),
.B2(n_11),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_149),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_167),
.Y(n_186)
);

BUFx24_ASAP7_75t_SL g196 ( 
.A(n_186),
.Y(n_196)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

XOR2x2_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_168),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_190),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_143),
.B1(n_157),
.B2(n_171),
.Y(n_190)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_184),
.B1(n_173),
.B2(n_180),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_195),
.C(n_198),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_174),
.B(n_16),
.CI(n_23),
.CON(n_194),
.SN(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_176),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_13),
.C(n_23),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_201),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_179),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_205),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_189),
.A2(n_7),
.B(n_1),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_12),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_199),
.C(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_193),
.C(n_196),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_213),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_193),
.C(n_194),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_7),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_216),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_202),
.B(n_7),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_2),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_207),
.C(n_23),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_3),
.B(n_4),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_222),
.B(n_224),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_217),
.B(n_5),
.Y(n_222)
);

AO21x1_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_227),
.B(n_223),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_3),
.C(n_4),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_228),
.B(n_219),
.Y(n_230)
);

AOI321xp33_ASAP7_75t_SL g227 ( 
.A1(n_221),
.A2(n_3),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C(n_0),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_SL g232 ( 
.A1(n_229),
.A2(n_230),
.B(n_8),
.C(n_10),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_8),
.C(n_9),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_232),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_233),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_234),
.A2(n_10),
.B(n_0),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_10),
.Y(n_236)
);


endmodule