module fake_jpeg_3450_n_689 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_689);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_689;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx11_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_58),
.Y(n_208)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_28),
.Y(n_59)
);

INVx5_ASAP7_75t_SL g176 ( 
.A(n_59),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_27),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_60),
.B(n_68),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_61),
.Y(n_157)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_62),
.Y(n_134)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_67),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_70),
.Y(n_168)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_71),
.Y(n_181)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_72),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_73),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_75),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_76),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_77),
.Y(n_173)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_79),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_80),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_82),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_84),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_24),
.B(n_35),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_88),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_87),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_11),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_91),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_92),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_93),
.Y(n_207)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

BUFx8_ASAP7_75t_L g197 ( 
.A(n_99),
.Y(n_197)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_100),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_101),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_105),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_38),
.B(n_11),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_124),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_52),
.Y(n_107)
);

INVx5_ASAP7_75t_SL g217 ( 
.A(n_107),
.Y(n_217)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_108),
.Y(n_230)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_114),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_116),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_118),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_120),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_47),
.B(n_10),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_33),
.B(n_45),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_21),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_43),
.Y(n_128)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_128),
.Y(n_226)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_129),
.Y(n_234)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_130),
.Y(n_235)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_131),
.Y(n_233)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_41),
.Y(n_132)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_59),
.A2(n_41),
.B1(n_34),
.B2(n_22),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_139),
.A2(n_169),
.B1(n_170),
.B2(n_211),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_75),
.A2(n_54),
.B1(n_37),
.B2(n_39),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_143),
.B(n_195),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_68),
.A2(n_54),
.B1(n_33),
.B2(n_45),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_147),
.A2(n_156),
.B1(n_159),
.B2(n_210),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_150),
.B(n_158),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_60),
.A2(n_41),
.B1(n_21),
.B2(n_20),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_153),
.A2(n_172),
.B1(n_182),
.B2(n_0),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_86),
.A2(n_41),
.B1(n_22),
.B2(n_20),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_25),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_41),
.B1(n_25),
.B2(n_39),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_88),
.B(n_40),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_162),
.B(n_171),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_107),
.A2(n_34),
.B1(n_40),
.B2(n_37),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_87),
.A2(n_106),
.B1(n_98),
.B2(n_82),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_125),
.B(n_34),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_128),
.A2(n_55),
.B1(n_50),
.B2(n_3),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_66),
.A2(n_55),
.B1(n_50),
.B2(n_13),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_108),
.B(n_13),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_186),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_69),
.B(n_12),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_187),
.B(n_192),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_73),
.B(n_12),
.Y(n_188)
);

INVxp67_ASAP7_75t_R g262 ( 
.A(n_188),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_74),
.B(n_14),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_76),
.B(n_14),
.Y(n_195)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_79),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_202),
.Y(n_317)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_80),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_81),
.B(n_19),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_224),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_83),
.A2(n_55),
.B1(n_50),
.B2(n_3),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_85),
.A2(n_50),
.B1(n_55),
.B2(n_115),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_90),
.A2(n_55),
.B1(n_50),
.B2(n_3),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_213),
.A2(n_215),
.B1(n_210),
.B2(n_211),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_96),
.B(n_9),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_2),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_123),
.A2(n_119),
.B1(n_112),
.B2(n_101),
.Y(n_215)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_99),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_220),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_59),
.A2(n_55),
.B1(n_9),
.B2(n_14),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_221),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_60),
.B(n_7),
.Y(n_224)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_63),
.Y(n_231)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_136),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_236),
.Y(n_346)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_237),
.Y(n_336)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_238),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_136),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_240),
.Y(n_326)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_241),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_140),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_243),
.A2(n_246),
.B1(n_248),
.B2(n_272),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_251),
.A2(n_254),
.B1(n_313),
.B2(n_314),
.Y(n_374)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_252),
.Y(n_340)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_164),
.Y(n_253)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_253),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_183),
.A2(n_15),
.B1(n_18),
.B2(n_17),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_152),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_198),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_256),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_257),
.B(n_295),
.Y(n_361)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_259),
.Y(n_337)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_151),
.Y(n_260)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_260),
.Y(n_327)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_261),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_176),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_263),
.B(n_264),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_176),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_137),
.B(n_15),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_265),
.B(n_288),
.Y(n_333)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_154),
.Y(n_266)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_178),
.Y(n_268)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_268),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_137),
.A2(n_15),
.B1(n_18),
.B2(n_17),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_269),
.B(n_287),
.Y(n_347)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_196),
.Y(n_270)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_270),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_140),
.B(n_9),
.C(n_16),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_271),
.B(n_285),
.C(n_201),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_224),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_134),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_273),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_170),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_274),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_145),
.A2(n_18),
.B1(n_19),
.B2(n_6),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_275),
.A2(n_315),
.B1(n_320),
.B2(n_321),
.Y(n_380)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_141),
.Y(n_276)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_276),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_155),
.A2(n_145),
.B1(n_192),
.B2(n_187),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_277),
.A2(n_292),
.B1(n_299),
.B2(n_319),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_161),
.Y(n_278)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_278),
.Y(n_366)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_134),
.Y(n_279)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_279),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_149),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_280),
.Y(n_385)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_218),
.Y(n_281)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_281),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_175),
.Y(n_282)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_282),
.Y(n_388)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_175),
.Y(n_283)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_283),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_146),
.B(n_19),
.C(n_5),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_149),
.Y(n_286)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_286),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_SL g287 ( 
.A(n_186),
.B(n_228),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_229),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_216),
.Y(n_289)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_289),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_150),
.B(n_4),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_296),
.Y(n_350)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_157),
.Y(n_291)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_291),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_172),
.A2(n_188),
.B1(n_214),
.B2(n_162),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_199),
.Y(n_293)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_293),
.Y(n_373)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_226),
.Y(n_294)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_294),
.Y(n_378)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_173),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_197),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_194),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_297),
.B(n_301),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_213),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_299)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_180),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_233),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_303),
.Y(n_362)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_184),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_190),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_304),
.B(n_305),
.Y(n_377)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_205),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_135),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_306),
.B(n_312),
.Y(n_363)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_207),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_307),
.Y(n_332)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_168),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_308),
.Y(n_376)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_142),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_309),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_230),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_310),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_158),
.Y(n_312)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_177),
.Y(n_313)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_208),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_181),
.B(n_5),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_163),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_318),
.Y(n_328)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_144),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_139),
.A2(n_5),
.B1(n_221),
.B2(n_169),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_204),
.B(n_212),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_143),
.A2(n_232),
.B1(n_200),
.B2(n_185),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_160),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_322),
.B(n_324),
.Y(n_370)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_225),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_323),
.A2(n_296),
.B1(n_314),
.B2(n_291),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_143),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_219),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_325),
.B(n_166),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_284),
.A2(n_292),
.B1(n_239),
.B2(n_246),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_330),
.A2(n_353),
.B1(n_368),
.B2(n_372),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_274),
.A2(n_232),
.B1(n_200),
.B2(n_185),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_335),
.A2(n_358),
.B1(n_372),
.B2(n_353),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_338),
.B(n_348),
.Y(n_415)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_298),
.B(n_165),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_341),
.Y(n_403)
);

AND2x2_ASAP7_75t_SL g343 ( 
.A(n_300),
.B(n_257),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_343),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_249),
.B(n_167),
.C(n_197),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_284),
.A2(n_133),
.B1(n_138),
.B2(n_148),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_247),
.A2(n_177),
.B1(n_179),
.B2(n_217),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_239),
.A2(n_191),
.B1(n_223),
.B2(n_225),
.Y(n_368)
);

AND2x2_ASAP7_75t_SL g371 ( 
.A(n_262),
.B(n_217),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_262),
.A2(n_166),
.B1(n_179),
.B2(n_189),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_375),
.B(n_386),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_243),
.B(n_271),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_268),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_285),
.B(n_242),
.C(n_322),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_342),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_389),
.B(n_390),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_329),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_370),
.A2(n_323),
.B1(n_266),
.B2(n_261),
.Y(n_391)
);

OAI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_391),
.A2(n_396),
.B1(n_409),
.B2(n_357),
.Y(n_473)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_328),
.Y(n_392)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_392),
.Y(n_440)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_333),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_393),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_354),
.A2(n_251),
.B(n_287),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_394),
.A2(n_359),
.B(n_378),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_352),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_395),
.B(n_397),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_328),
.Y(n_397)
);

XOR2x2_ASAP7_75t_SL g398 ( 
.A(n_330),
.B(n_269),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_398),
.B(n_408),
.Y(n_479)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_375),
.Y(n_399)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_399),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_354),
.A2(n_244),
.B(n_254),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_400),
.A2(n_384),
.B(n_332),
.Y(n_439)
);

AO22x1_ASAP7_75t_SL g401 ( 
.A1(n_345),
.A2(n_318),
.B1(n_305),
.B2(n_304),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_401),
.B(n_418),
.Y(n_454)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_388),
.Y(n_402)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_402),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_350),
.B(n_267),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_405),
.B(n_407),
.Y(n_442)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_388),
.Y(n_406)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_406),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_387),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_368),
.A2(n_295),
.B1(n_297),
.B2(n_307),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_377),
.Y(n_410)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_410),
.Y(n_451)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_387),
.Y(n_411)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_411),
.Y(n_459)
);

NAND2xp67_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_270),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_412),
.B(n_423),
.Y(n_478)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_387),
.Y(n_416)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_416),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_355),
.A2(n_236),
.B1(n_301),
.B2(n_294),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_417),
.A2(n_420),
.B1(n_426),
.B2(n_430),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_281),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_355),
.A2(n_245),
.B1(n_317),
.B2(n_282),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_419),
.A2(n_428),
.B1(n_432),
.B2(n_433),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_380),
.A2(n_240),
.B1(n_286),
.B2(n_280),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_356),
.Y(n_421)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_421),
.Y(n_474)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_356),
.Y(n_422)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_422),
.Y(n_482)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_334),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_255),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_436),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_380),
.A2(n_313),
.B1(n_317),
.B2(n_238),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_334),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_427),
.B(n_429),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_345),
.A2(n_260),
.B1(n_311),
.B2(n_278),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_337),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_343),
.A2(n_250),
.B1(n_347),
.B2(n_341),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_336),
.B(n_250),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_431),
.B(n_434),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_386),
.A2(n_347),
.B1(n_338),
.B2(n_361),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_361),
.A2(n_363),
.B1(n_348),
.B2(n_371),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_336),
.B(n_363),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_343),
.A2(n_341),
.B1(n_374),
.B2(n_361),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_435),
.A2(n_385),
.B1(n_326),
.B2(n_369),
.Y(n_467)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

OA21x2_ASAP7_75t_L g438 ( 
.A1(n_364),
.A2(n_362),
.B(n_360),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_339),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_439),
.A2(n_450),
.B(n_480),
.Y(n_523)
);

AOI22x1_ASAP7_75t_SL g445 ( 
.A1(n_435),
.A2(n_369),
.B1(n_357),
.B2(n_326),
.Y(n_445)
);

OA22x2_ASAP7_75t_L g503 ( 
.A1(n_445),
.A2(n_462),
.B1(n_409),
.B2(n_391),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_438),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_452),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_415),
.B(n_351),
.C(n_373),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_448),
.B(n_465),
.C(n_477),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_413),
.A2(n_351),
.B1(n_365),
.B2(n_346),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_449),
.A2(n_464),
.B1(n_407),
.B2(n_428),
.Y(n_484)
);

A2O1A1Ixp33_ASAP7_75t_L g452 ( 
.A1(n_425),
.A2(n_379),
.B(n_376),
.C(n_349),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_438),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_461),
.B(n_466),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_397),
.A2(n_365),
.B1(n_326),
.B2(n_385),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_413),
.A2(n_432),
.B1(n_428),
.B2(n_399),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_415),
.B(n_373),
.C(n_360),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_438),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_467),
.A2(n_470),
.B1(n_471),
.B2(n_396),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_392),
.B(n_379),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_468),
.B(n_469),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_418),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_417),
.A2(n_376),
.B1(n_346),
.B2(n_344),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_408),
.A2(n_346),
.B1(n_344),
.B2(n_331),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_473),
.A2(n_426),
.B1(n_420),
.B2(n_414),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_437),
.A2(n_367),
.B(n_349),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_475),
.A2(n_412),
.B(n_422),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_404),
.B(n_339),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_481),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_415),
.B(n_367),
.C(n_359),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_404),
.B(n_378),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_483),
.A2(n_484),
.B1(n_445),
.B2(n_460),
.Y(n_537)
);

FAx1_ASAP7_75t_SL g485 ( 
.A(n_448),
.B(n_430),
.CI(n_403),
.CON(n_485),
.SN(n_485)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_485),
.B(n_491),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_464),
.A2(n_424),
.B1(n_394),
.B2(n_432),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_486),
.A2(n_522),
.B1(n_459),
.B2(n_472),
.Y(n_533)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_487),
.Y(n_526)
);

AO22x1_ASAP7_75t_L g488 ( 
.A1(n_447),
.A2(n_434),
.B1(n_414),
.B2(n_398),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_488),
.Y(n_546)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_458),
.Y(n_489)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_489),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_455),
.B(n_442),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_442),
.B(n_405),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_492),
.B(n_493),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_451),
.B(n_389),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_465),
.B(n_433),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_494),
.B(n_514),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_477),
.B(n_403),
.C(n_398),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_495),
.B(n_498),
.C(n_501),
.Y(n_528)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_458),
.Y(n_496)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_496),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_410),
.C(n_411),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_456),
.Y(n_499)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_499),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_481),
.B(n_479),
.C(n_463),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_451),
.B(n_390),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_502),
.B(n_505),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_503),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_416),
.C(n_406),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_504),
.B(n_509),
.C(n_517),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_453),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_478),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_507),
.B(n_471),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_453),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_508),
.B(n_519),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_463),
.B(n_402),
.C(n_394),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_461),
.A2(n_400),
.B(n_431),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_510),
.A2(n_439),
.B(n_480),
.Y(n_524)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_456),
.Y(n_511)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_511),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_466),
.A2(n_419),
.B1(n_414),
.B2(n_401),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_513),
.A2(n_516),
.B1(n_521),
.B2(n_452),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_440),
.B(n_401),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_515),
.A2(n_480),
.B(n_478),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_450),
.A2(n_401),
.B1(n_412),
.B2(n_427),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_440),
.B(n_421),
.C(n_423),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_443),
.Y(n_518)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_518),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_468),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_444),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_520),
.B(n_482),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_450),
.A2(n_469),
.B1(n_454),
.B2(n_460),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_449),
.A2(n_429),
.B1(n_395),
.B2(n_436),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_524),
.A2(n_547),
.B(n_559),
.Y(n_588)
);

MAJx2_ASAP7_75t_L g532 ( 
.A(n_494),
.B(n_444),
.C(n_441),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_SL g562 ( 
.A(n_532),
.B(n_557),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_533),
.A2(n_545),
.B1(n_554),
.B2(n_558),
.Y(n_563)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_535),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_SL g573 ( 
.A1(n_537),
.A2(n_526),
.B1(n_529),
.B2(n_558),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_490),
.B(n_441),
.C(n_459),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_540),
.B(n_507),
.C(n_511),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_488),
.A2(n_478),
.B1(n_472),
.B2(n_445),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_543),
.Y(n_568)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_500),
.Y(n_544)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_544),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_521),
.A2(n_454),
.B1(n_452),
.B2(n_457),
.Y(n_545)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_548),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_517),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_549),
.B(n_506),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_498),
.B(n_331),
.Y(n_550)
);

CKINVDCx14_ASAP7_75t_R g564 ( 
.A(n_550),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_500),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_551),
.B(n_555),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_490),
.B(n_457),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_504),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_523),
.A2(n_467),
.B1(n_475),
.B2(n_470),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_489),
.B(n_446),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_556),
.B(n_561),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_SL g557 ( 
.A(n_495),
.B(n_501),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_486),
.A2(n_462),
.B1(n_446),
.B2(n_443),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_523),
.A2(n_482),
.B(n_474),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_499),
.A2(n_474),
.B1(n_327),
.B2(n_366),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_560),
.A2(n_487),
.B1(n_513),
.B2(n_516),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_496),
.B(n_383),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_565),
.B(n_567),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_534),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_566),
.B(n_577),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_570),
.A2(n_573),
.B1(n_587),
.B2(n_545),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_557),
.B(n_509),
.C(n_512),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_572),
.B(n_576),
.C(n_590),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_553),
.B(n_512),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_575),
.B(n_585),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_528),
.B(n_510),
.C(n_515),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_552),
.B(n_327),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_578),
.B(n_581),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_556),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_SL g582 ( 
.A(n_530),
.B(n_488),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_582),
.B(n_583),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_SL g583 ( 
.A(n_530),
.B(n_485),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_506),
.Y(n_584)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_584),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_528),
.B(n_485),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_552),
.B(n_497),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_586),
.B(n_589),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_526),
.A2(n_497),
.B1(n_484),
.B2(n_514),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_540),
.B(n_340),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_538),
.B(n_532),
.C(n_531),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_538),
.B(n_522),
.C(n_503),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_591),
.B(n_537),
.C(n_529),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_541),
.B(n_483),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_592),
.B(n_554),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g628 ( 
.A(n_595),
.B(n_607),
.Y(n_628)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_579),
.Y(n_598)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_598),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_580),
.A2(n_544),
.B1(n_533),
.B2(n_535),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_601),
.A2(n_613),
.B1(n_587),
.B2(n_592),
.Y(n_629)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_574),
.Y(n_604)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_604),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_588),
.A2(n_524),
.B(n_547),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_605),
.A2(n_611),
.B(n_569),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_584),
.B(n_539),
.Y(n_606)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_606),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_565),
.B(n_559),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_567),
.B(n_543),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_608),
.B(n_609),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_590),
.B(n_541),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_610),
.B(n_612),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_571),
.A2(n_546),
.B(n_539),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_575),
.B(n_576),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_572),
.B(n_536),
.C(n_527),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_614),
.B(n_564),
.C(n_582),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_588),
.A2(n_546),
.B(n_525),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_615),
.A2(n_555),
.B(n_561),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_585),
.B(n_562),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_616),
.B(n_617),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_571),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_SL g618 ( 
.A1(n_563),
.A2(n_536),
.B1(n_527),
.B2(n_531),
.Y(n_618)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_618),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_620),
.B(n_634),
.Y(n_641)
);

BUFx24_ASAP7_75t_SL g621 ( 
.A(n_609),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g646 ( 
.A(n_621),
.B(n_638),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_606),
.B(n_574),
.Y(n_622)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_622),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_624),
.A2(n_637),
.B(n_639),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_601),
.A2(n_563),
.B1(n_570),
.B2(n_580),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_625),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_597),
.B(n_591),
.C(n_562),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_626),
.B(n_627),
.C(n_594),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_597),
.B(n_583),
.C(n_568),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_629),
.B(n_607),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_599),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_631),
.B(n_602),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_SL g634 ( 
.A1(n_596),
.A2(n_605),
.B1(n_595),
.B2(n_611),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_614),
.B(n_560),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_615),
.A2(n_542),
.B(n_503),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g640 ( 
.A1(n_618),
.A2(n_542),
.B1(n_503),
.B2(n_366),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_L g650 ( 
.A(n_640),
.B(n_603),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_643),
.B(n_648),
.Y(n_666)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_644),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_623),
.A2(n_593),
.B1(n_610),
.B2(n_608),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_SL g669 ( 
.A1(n_645),
.A2(n_625),
.B1(n_639),
.B2(n_637),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_619),
.A2(n_612),
.B(n_603),
.Y(n_649)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_649),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_650),
.B(n_651),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g651 ( 
.A(n_631),
.B(n_594),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_624),
.A2(n_616),
.B(n_600),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_652),
.A2(n_627),
.B(n_626),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_634),
.B(n_600),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_653),
.B(n_654),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_620),
.B(n_340),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_633),
.B(n_383),
.C(n_381),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_655),
.B(n_628),
.C(n_623),
.Y(n_664)
);

XNOR2xp5_ASAP7_75t_L g656 ( 
.A(n_633),
.B(n_381),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_656),
.B(n_628),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_658),
.B(n_669),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_642),
.B(n_622),
.Y(n_661)
);

OAI21x1_ASAP7_75t_SL g670 ( 
.A1(n_661),
.A2(n_657),
.B(n_641),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_646),
.B(n_632),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_662),
.B(n_645),
.Y(n_674)
);

XNOR2xp5_ASAP7_75t_L g672 ( 
.A(n_664),
.B(n_665),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_SL g665 ( 
.A1(n_642),
.A2(n_640),
.B1(n_636),
.B2(n_635),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_SL g671 ( 
.A(n_668),
.B(n_641),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_670),
.B(n_671),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_659),
.A2(n_643),
.B(n_652),
.Y(n_673)
);

OAI321xp33_ASAP7_75t_L g682 ( 
.A1(n_673),
.A2(n_661),
.A3(n_658),
.B1(n_669),
.B2(n_630),
.C(n_647),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_674),
.B(n_676),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_SL g676 ( 
.A1(n_660),
.A2(n_657),
.B(n_647),
.Y(n_676)
);

XNOR2xp5_ASAP7_75t_L g677 ( 
.A(n_668),
.B(n_648),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g678 ( 
.A(n_677),
.B(n_666),
.C(n_664),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_678),
.B(n_681),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g681 ( 
.A(n_672),
.B(n_663),
.C(n_667),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_682),
.A2(n_671),
.B(n_675),
.Y(n_684)
);

INVxp33_ASAP7_75t_L g685 ( 
.A(n_684),
.Y(n_685)
);

MAJIxp5_ASAP7_75t_L g686 ( 
.A(n_685),
.B(n_683),
.C(n_680),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_686),
.A2(n_679),
.B(n_675),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_687),
.A2(n_630),
.B(n_650),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_688),
.B(n_655),
.Y(n_689)
);


endmodule