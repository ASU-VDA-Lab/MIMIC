module fake_jpeg_16665_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_18),
.Y(n_23)
);

OR2x2_ASAP7_75t_SL g16 ( 
.A(n_10),
.B(n_1),
.Y(n_16)
);

OA22x2_ASAP7_75t_L g27 ( 
.A1(n_16),
.A2(n_20),
.B1(n_21),
.B2(n_12),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_11),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_26),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_6),
.B1(n_12),
.B2(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_17),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_32),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_33),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_27),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_31),
.B1(n_29),
.B2(n_26),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_27),
.Y(n_41)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_38),
.A3(n_27),
.B1(n_24),
.B2(n_37),
.C1(n_21),
.C2(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_22),
.Y(n_43)
);


endmodule