module fake_jpeg_8829_n_229 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_118;
wire n_128;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_SL g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_37),
.B(n_45),
.Y(n_73)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_47),
.Y(n_51)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_20),
.Y(n_54)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_35),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_28),
.B1(n_25),
.B2(n_18),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_61),
.B1(n_43),
.B2(n_48),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_28),
.B1(n_25),
.B2(n_29),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_67),
.B1(n_21),
.B2(n_22),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_19),
.B(n_29),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_30),
.C(n_17),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_28),
.B1(n_19),
.B2(n_27),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_27),
.B1(n_35),
.B2(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_31),
.Y(n_71)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_26),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_46),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_41),
.Y(n_76)
);

CKINVDCx9p33_ASAP7_75t_R g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_78),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_79),
.B(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_83),
.B(n_102),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_47),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_89),
.Y(n_116)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_86),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

AND2x4_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_23),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_95),
.B1(n_107),
.B2(n_66),
.Y(n_124)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_103),
.Y(n_110)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_0),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_100),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_0),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_21),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_24),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_1),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_22),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_42),
.B1(n_43),
.B2(n_24),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_51),
.Y(n_114)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_87),
.B(n_53),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_60),
.C(n_76),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_92),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_90),
.B1(n_89),
.B2(n_60),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_107),
.B1(n_68),
.B2(n_66),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_33),
.A3(n_32),
.B1(n_52),
.B2(n_72),
.Y(n_126)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_81),
.A2(n_56),
.B1(n_66),
.B2(n_52),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_111),
.B1(n_127),
.B2(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_81),
.B(n_72),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_88),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_144),
.C(n_123),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_136),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_150),
.B(n_154),
.Y(n_161)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_110),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_151),
.C(n_2),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_143),
.B1(n_111),
.B2(n_131),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_1),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_82),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_108),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_148),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_105),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_149),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_122),
.A2(n_68),
.B(n_78),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_109),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_101),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

OR2x2_ASAP7_75t_SL g155 ( 
.A(n_125),
.B(n_32),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_113),
.B(n_116),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_159),
.A2(n_162),
.B(n_163),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_116),
.B1(n_121),
.B2(n_126),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_133),
.C(n_144),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_155),
.B(n_154),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_150),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_141),
.A2(n_138),
.B(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_169),
.B(n_172),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_132),
.B1(n_130),
.B2(n_123),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_123),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_163),
.C(n_167),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_112),
.A3(n_32),
.B1(n_46),
.B2(n_23),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_143),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_173),
.B(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_15),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_187),
.B1(n_188),
.B2(n_157),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_182),
.B(n_184),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_162),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_185),
.C(n_186),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_140),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_137),
.C(n_135),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_135),
.C(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_152),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_166),
.B(n_146),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_160),
.C(n_170),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_190),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_199),
.Y(n_204)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_184),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_172),
.C(n_156),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_197),
.C(n_180),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_156),
.C(n_136),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_132),
.B1(n_130),
.B2(n_106),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_198),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_206)
);

FAx1_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_2),
.CI(n_3),
.CON(n_199),
.SN(n_199)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_177),
.A2(n_99),
.B1(n_10),
.B2(n_11),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_14),
.B(n_5),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_200),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_206),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_14),
.B1(n_15),
.B2(n_6),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_208),
.A2(n_209),
.B(n_210),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_199),
.B1(n_195),
.B2(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_203),
.B(n_191),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_216),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_207),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_7),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_208),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_209),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_217),
.A2(n_218),
.B(n_211),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_204),
.Y(n_218)
);

INVx11_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_205),
.B(n_212),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_220),
.B(n_204),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_226),
.B(n_224),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_221),
.Y(n_229)
);


endmodule