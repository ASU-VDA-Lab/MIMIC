module real_aes_7305_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_505;
wire n_434;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_SL g132 ( .A1(n_0), .A2(n_29), .B1(n_133), .B2(n_137), .Y(n_132) );
INVx1_ASAP7_75t_L g213 ( .A(n_1), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_2), .A2(n_167), .B1(n_168), .B2(n_169), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_2), .Y(n_167) );
AOI21xp33_ASAP7_75t_L g245 ( .A1(n_2), .A2(n_229), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g185 ( .A(n_3), .Y(n_185) );
AND2x6_ASAP7_75t_L g207 ( .A(n_3), .B(n_183), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_3), .B(n_508), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_4), .A2(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g251 ( .A(n_5), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_6), .B(n_308), .Y(n_307) );
AO22x2_ASAP7_75t_L g86 ( .A1(n_7), .A2(n_24), .B1(n_87), .B2(n_88), .Y(n_86) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_8), .A2(n_12), .B1(n_142), .B2(n_145), .Y(n_141) );
INVx1_ASAP7_75t_L g199 ( .A(n_9), .Y(n_199) );
INVx1_ASAP7_75t_L g322 ( .A(n_10), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g98 ( .A1(n_11), .A2(n_47), .B1(n_99), .B2(n_104), .Y(n_98) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_13), .A2(n_25), .B1(n_87), .B2(n_91), .Y(n_90) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_14), .B(n_234), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_15), .B(n_229), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_16), .B(n_241), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g319 ( .A1(n_17), .A2(n_320), .B(n_321), .C(n_323), .Y(n_319) );
OAI22xp5_ASAP7_75t_SL g164 ( .A1(n_18), .A2(n_165), .B1(n_166), .B2(n_172), .Y(n_164) );
INVx1_ASAP7_75t_L g172 ( .A(n_18), .Y(n_172) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_19), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_20), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g266 ( .A(n_21), .Y(n_266) );
AOI22xp33_ASAP7_75t_SL g149 ( .A1(n_22), .A2(n_36), .B1(n_150), .B2(n_153), .Y(n_149) );
INVx2_ASAP7_75t_L g205 ( .A(n_23), .Y(n_205) );
OAI221xp5_ASAP7_75t_L g176 ( .A1(n_25), .A2(n_41), .B1(n_50), .B2(n_177), .C(n_178), .Y(n_176) );
INVxp67_ASAP7_75t_L g179 ( .A(n_25), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_26), .A2(n_80), .B1(n_162), .B2(n_163), .Y(n_79) );
INVx1_ASAP7_75t_L g162 ( .A(n_26), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_27), .A2(n_207), .B(n_209), .C(n_281), .Y(n_280) );
AOI22xp33_ASAP7_75t_SL g121 ( .A1(n_28), .A2(n_61), .B1(n_122), .B2(n_126), .Y(n_121) );
INVx1_ASAP7_75t_L g264 ( .A(n_30), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_31), .B(n_217), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_32), .B(n_118), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_33), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_34), .B(n_229), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_35), .A2(n_37), .B1(n_157), .B2(n_159), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_38), .A2(n_209), .B1(n_219), .B2(n_262), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g289 ( .A(n_39), .Y(n_289) );
CKINVDCx16_ASAP7_75t_R g201 ( .A(n_40), .Y(n_201) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_41), .A2(n_60), .B1(n_87), .B2(n_91), .Y(n_94) );
INVxp67_ASAP7_75t_L g180 ( .A(n_41), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_42), .A2(n_237), .B(n_249), .C(n_250), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_43), .Y(n_299) );
INVx1_ASAP7_75t_L g247 ( .A(n_44), .Y(n_247) );
INVx1_ASAP7_75t_L g183 ( .A(n_45), .Y(n_183) );
INVx1_ASAP7_75t_L g198 ( .A(n_46), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_48), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_49), .Y(n_97) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_50), .A2(n_66), .B1(n_87), .B2(n_88), .Y(n_96) );
OAI22xp5_ASAP7_75t_SL g169 ( .A1(n_51), .A2(n_58), .B1(n_170), .B2(n_171), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g170 ( .A(n_51), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_SL g233 ( .A1(n_52), .A2(n_234), .B(n_235), .C(n_237), .Y(n_233) );
INVxp67_ASAP7_75t_L g236 ( .A(n_53), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_54), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_55), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g292 ( .A(n_56), .Y(n_292) );
A2O1A1Ixp33_ASAP7_75t_L g293 ( .A1(n_57), .A2(n_207), .B(n_209), .C(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g171 ( .A(n_58), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_59), .A2(n_80), .B1(n_163), .B2(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_59), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_62), .B(n_214), .Y(n_282) );
INVx2_ASAP7_75t_L g196 ( .A(n_63), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_64), .B(n_234), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_65), .A2(n_207), .B(n_209), .C(n_212), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_67), .B(n_224), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_68), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g304 ( .A1(n_69), .A2(n_207), .B(n_209), .C(n_305), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_70), .Y(n_312) );
INVx1_ASAP7_75t_L g232 ( .A(n_71), .Y(n_232) );
CKINVDCx16_ASAP7_75t_R g318 ( .A(n_72), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_73), .B(n_214), .Y(n_306) );
INVx1_ASAP7_75t_L g87 ( .A(n_74), .Y(n_87) );
INVx1_ASAP7_75t_L g89 ( .A(n_74), .Y(n_89) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_75), .B(n_227), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_76), .A2(n_229), .B(n_230), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_76), .A2(n_80), .B1(n_163), .B2(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_76), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_173), .B1(n_186), .B2(n_498), .C(n_502), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_164), .Y(n_78) );
INVx1_ASAP7_75t_L g163 ( .A(n_80), .Y(n_163) );
AND2x4_ASAP7_75t_L g80 ( .A(n_81), .B(n_130), .Y(n_80) );
NOR2xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_108), .Y(n_81) );
OAI21xp5_ASAP7_75t_SL g82 ( .A1(n_83), .A2(n_97), .B(n_98), .Y(n_82) );
INVx4_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
AND2x6_ASAP7_75t_L g84 ( .A(n_85), .B(n_92), .Y(n_84) );
AND2x4_ASAP7_75t_L g105 ( .A(n_85), .B(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_90), .Y(n_85) );
AND2x2_ASAP7_75t_L g103 ( .A(n_86), .B(n_94), .Y(n_103) );
INVx2_ASAP7_75t_L g116 ( .A(n_86), .Y(n_116) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g91 ( .A(n_89), .Y(n_91) );
OR2x2_ASAP7_75t_L g115 ( .A(n_90), .B(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g120 ( .A(n_90), .B(n_116), .Y(n_120) );
INVx2_ASAP7_75t_L g125 ( .A(n_90), .Y(n_125) );
INVx1_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
AND2x2_ASAP7_75t_L g144 ( .A(n_92), .B(n_136), .Y(n_144) );
AND2x6_ASAP7_75t_L g147 ( .A(n_92), .B(n_114), .Y(n_147) );
AND2x4_ASAP7_75t_L g152 ( .A(n_92), .B(n_120), .Y(n_152) );
AND2x2_ASAP7_75t_L g92 ( .A(n_93), .B(n_95), .Y(n_92) );
AND2x2_ASAP7_75t_L g113 ( .A(n_93), .B(n_96), .Y(n_113) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
AND2x2_ASAP7_75t_L g135 ( .A(n_94), .B(n_107), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_94), .B(n_96), .Y(n_140) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g102 ( .A(n_96), .Y(n_102) );
INVx1_ASAP7_75t_L g107 ( .A(n_96), .Y(n_107) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x4_ASAP7_75t_L g100 ( .A(n_101), .B(n_103), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g124 ( .A(n_102), .B(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g123 ( .A(n_103), .B(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g127 ( .A(n_103), .B(n_128), .Y(n_127) );
BUFx2_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND3xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_117), .C(n_121), .Y(n_108) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx4_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x6_ASAP7_75t_L g119 ( .A(n_113), .B(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g158 ( .A(n_113), .B(n_136), .Y(n_158) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g136 ( .A(n_116), .B(n_125), .Y(n_136) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g155 ( .A(n_120), .B(n_135), .Y(n_155) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OR2x6_ASAP7_75t_L g161 ( .A(n_129), .B(n_140), .Y(n_161) );
NOR2x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_148), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_141), .Y(n_131) );
BUFx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x4_ASAP7_75t_L g138 ( .A(n_136), .B(n_139), .Y(n_138) );
BUFx2_ASAP7_75t_SL g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx4_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx11_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_156), .Y(n_148) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx6_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx8_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx6_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_166), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
AND3x1_ASAP7_75t_SL g175 ( .A(n_176), .B(n_181), .C(n_184), .Y(n_175) );
INVxp67_ASAP7_75t_L g508 ( .A(n_176), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_181), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_181), .A2(n_209), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g518 ( .A(n_181), .Y(n_518) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_182), .B(n_185), .Y(n_512) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OR2x2_ASAP7_75t_SL g517 ( .A(n_184), .B(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
BUFx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2x1_ASAP7_75t_L g187 ( .A(n_188), .B(n_414), .Y(n_187) );
NOR5xp2_ASAP7_75t_L g188 ( .A(n_189), .B(n_337), .C(n_369), .D(n_384), .E(n_401), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_253), .B(n_274), .C(n_325), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_225), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_191), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_191), .B(n_389), .Y(n_452) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_192), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_192), .B(n_271), .Y(n_338) );
AND2x2_ASAP7_75t_L g379 ( .A(n_192), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_192), .B(n_348), .Y(n_383) );
OR2x2_ASAP7_75t_L g420 ( .A(n_192), .B(n_259), .Y(n_420) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g258 ( .A(n_193), .B(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g328 ( .A(n_193), .Y(n_328) );
OR2x2_ASAP7_75t_L g491 ( .A(n_193), .B(n_331), .Y(n_491) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_200), .B(n_221), .Y(n_193) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_194), .A2(n_260), .B(n_268), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_194), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g287 ( .A(n_194), .Y(n_287) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_195), .Y(n_227) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
AND2x2_ASAP7_75t_SL g224 ( .A(n_196), .B(n_197), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_208), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g260 ( .A1(n_202), .A2(n_239), .B1(n_261), .B2(n_267), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g291 ( .A1(n_202), .A2(n_292), .B(n_293), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g202 ( .A(n_203), .B(n_207), .Y(n_202) );
AND2x4_ASAP7_75t_L g229 ( .A(n_203), .B(n_207), .Y(n_229) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_206), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g210 ( .A(n_205), .Y(n_210) );
INVx1_ASAP7_75t_L g220 ( .A(n_205), .Y(n_220) );
INVx1_ASAP7_75t_L g211 ( .A(n_206), .Y(n_211) );
INVx3_ASAP7_75t_L g215 ( .A(n_206), .Y(n_215) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_206), .Y(n_217) );
INVx1_ASAP7_75t_L g234 ( .A(n_206), .Y(n_234) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_206), .Y(n_263) );
INVx4_ASAP7_75t_SL g239 ( .A(n_207), .Y(n_239) );
BUFx3_ASAP7_75t_L g501 ( .A(n_207), .Y(n_501) );
INVx5_ASAP7_75t_L g231 ( .A(n_209), .Y(n_231) );
AND2x2_ASAP7_75t_L g500 ( .A(n_209), .B(n_501), .Y(n_500) );
AND2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_210), .Y(n_238) );
BUFx3_ASAP7_75t_L g286 ( .A(n_210), .Y(n_286) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_216), .C(n_218), .Y(n_212) );
INVx5_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_215), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_215), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g249 ( .A(n_217), .Y(n_249) );
INVx4_ASAP7_75t_L g308 ( .A(n_217), .Y(n_308) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_223), .B(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_223), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g302 ( .A(n_224), .Y(n_302) );
OA21x2_ASAP7_75t_L g314 ( .A1(n_224), .A2(n_315), .B(n_324), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_225), .A2(n_394), .B1(n_395), .B2(n_398), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_225), .B(n_328), .Y(n_477) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_243), .Y(n_225) );
AND2x2_ASAP7_75t_L g273 ( .A(n_226), .B(n_259), .Y(n_273) );
AND2x2_ASAP7_75t_L g330 ( .A(n_226), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g335 ( .A(n_226), .Y(n_335) );
INVx3_ASAP7_75t_L g348 ( .A(n_226), .Y(n_348) );
OR2x2_ASAP7_75t_L g368 ( .A(n_226), .B(n_331), .Y(n_368) );
AND2x2_ASAP7_75t_L g387 ( .A(n_226), .B(n_244), .Y(n_387) );
BUFx2_ASAP7_75t_L g419 ( .A(n_226), .Y(n_419) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_240), .Y(n_226) );
INVx4_ASAP7_75t_L g242 ( .A(n_227), .Y(n_242) );
BUFx2_ASAP7_75t_L g316 ( .A(n_229), .Y(n_316) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .C(n_239), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_231), .A2(n_239), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_231), .A2(n_239), .B(n_318), .C(n_319), .Y(n_317) );
OAI322xp33_ASAP7_75t_L g502 ( .A1(n_232), .A2(n_503), .A3(n_505), .B1(n_509), .B2(n_510), .C1(n_513), .C2(n_515), .Y(n_502) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_238), .Y(n_309) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_241), .A2(n_245), .B(n_252), .Y(n_244) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_SL g288 ( .A(n_242), .B(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g334 ( .A(n_243), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
BUFx2_ASAP7_75t_L g257 ( .A(n_244), .Y(n_257) );
INVx2_ASAP7_75t_L g272 ( .A(n_244), .Y(n_272) );
OR2x2_ASAP7_75t_L g350 ( .A(n_244), .B(n_331), .Y(n_350) );
AND2x2_ASAP7_75t_L g380 ( .A(n_244), .B(n_259), .Y(n_380) );
AND2x2_ASAP7_75t_L g397 ( .A(n_244), .B(n_328), .Y(n_397) );
AND2x2_ASAP7_75t_L g437 ( .A(n_244), .B(n_348), .Y(n_437) );
AND2x2_ASAP7_75t_SL g473 ( .A(n_244), .B(n_273), .Y(n_473) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp33_ASAP7_75t_SL g254 ( .A(n_255), .B(n_270), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_256), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
OAI21xp33_ASAP7_75t_L g411 ( .A1(n_257), .A2(n_273), .B(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_257), .B(n_259), .Y(n_467) );
AND2x2_ASAP7_75t_L g403 ( .A(n_258), .B(n_404), .Y(n_403) );
INVx3_ASAP7_75t_L g331 ( .A(n_259), .Y(n_331) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_259), .Y(n_429) );
OAI22xp5_ASAP7_75t_SL g262 ( .A1(n_263), .A2(n_264), .B1(n_265), .B2(n_266), .Y(n_262) );
INVx2_ASAP7_75t_L g265 ( .A(n_263), .Y(n_265) );
INVx4_ASAP7_75t_L g320 ( .A(n_263), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_270), .B(n_328), .Y(n_496) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_271), .A2(n_439), .B1(n_440), .B2(n_445), .Y(n_438) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
AND2x2_ASAP7_75t_L g329 ( .A(n_272), .B(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g367 ( .A(n_272), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g404 ( .A(n_272), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_273), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g458 ( .A(n_273), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_300), .Y(n_275) );
INVx4_ASAP7_75t_L g344 ( .A(n_276), .Y(n_344) );
AND2x2_ASAP7_75t_L g422 ( .A(n_276), .B(n_389), .Y(n_422) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_290), .Y(n_276) );
INVx3_ASAP7_75t_L g341 ( .A(n_277), .Y(n_341) );
AND2x2_ASAP7_75t_L g355 ( .A(n_277), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_277), .Y(n_359) );
INVx2_ASAP7_75t_L g373 ( .A(n_277), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_277), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g430 ( .A(n_277), .B(n_425), .Y(n_430) );
AND2x2_ASAP7_75t_L g495 ( .A(n_277), .B(n_465), .Y(n_495) );
OR2x6_ASAP7_75t_L g277 ( .A(n_278), .B(n_288), .Y(n_277) );
AOI21xp5_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_280), .B(n_287), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_284), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_284), .A2(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g323 ( .A(n_286), .Y(n_323) );
INVx1_ASAP7_75t_L g297 ( .A(n_287), .Y(n_297) );
AND2x2_ASAP7_75t_L g336 ( .A(n_290), .B(n_314), .Y(n_336) );
INVx2_ASAP7_75t_L g356 ( .A(n_290), .Y(n_356) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_297), .B(n_298), .Y(n_290) );
INVx1_ASAP7_75t_L g361 ( .A(n_300), .Y(n_361) );
AND2x2_ASAP7_75t_L g407 ( .A(n_300), .B(n_355), .Y(n_407) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_313), .Y(n_300) );
INVx2_ASAP7_75t_L g346 ( .A(n_301), .Y(n_346) );
INVx1_ASAP7_75t_L g354 ( .A(n_301), .Y(n_354) );
AND2x2_ASAP7_75t_L g372 ( .A(n_301), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_301), .B(n_356), .Y(n_410) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B(n_311), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_310), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B(n_309), .Y(n_305) );
AND2x2_ASAP7_75t_L g389 ( .A(n_313), .B(n_346), .Y(n_389) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g342 ( .A(n_314), .Y(n_342) );
AND2x2_ASAP7_75t_L g425 ( .A(n_314), .B(n_356), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_320), .B(n_322), .Y(n_321) );
OAI21xp5_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_332), .B(n_336), .Y(n_325) );
INVx1_ASAP7_75t_SL g370 ( .A(n_326), .Y(n_370) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_327), .B(n_334), .Y(n_427) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g376 ( .A(n_328), .B(n_331), .Y(n_376) );
AND2x2_ASAP7_75t_L g405 ( .A(n_328), .B(n_349), .Y(n_405) );
OR2x2_ASAP7_75t_L g408 ( .A(n_328), .B(n_368), .Y(n_408) );
AOI222xp33_ASAP7_75t_L g472 ( .A1(n_329), .A2(n_421), .B1(n_473), .B2(n_474), .C1(n_476), .C2(n_478), .Y(n_472) );
BUFx2_ASAP7_75t_L g386 ( .A(n_331), .Y(n_386) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g375 ( .A(n_334), .B(n_376), .Y(n_375) );
INVx3_ASAP7_75t_SL g392 ( .A(n_334), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_334), .B(n_386), .Y(n_446) );
AND2x2_ASAP7_75t_L g381 ( .A(n_336), .B(n_341), .Y(n_381) );
INVx1_ASAP7_75t_L g400 ( .A(n_336), .Y(n_400) );
OAI221xp5_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_339), .B1(n_343), .B2(n_347), .C(n_351), .Y(n_337) );
OR2x2_ASAP7_75t_L g409 ( .A(n_339), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g394 ( .A(n_341), .B(n_364), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_341), .B(n_354), .Y(n_434) );
AND2x2_ASAP7_75t_L g439 ( .A(n_341), .B(n_389), .Y(n_439) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_341), .Y(n_449) );
NAND2x1_ASAP7_75t_SL g460 ( .A(n_341), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g345 ( .A(n_342), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g365 ( .A(n_342), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_342), .B(n_360), .Y(n_391) );
INVx1_ASAP7_75t_L g457 ( .A(n_342), .Y(n_457) );
INVx1_ASAP7_75t_L g432 ( .A(n_343), .Y(n_432) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g444 ( .A(n_344), .Y(n_444) );
NOR2xp67_ASAP7_75t_L g456 ( .A(n_344), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g461 ( .A(n_345), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_345), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g364 ( .A(n_346), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_346), .B(n_356), .Y(n_377) );
INVx1_ASAP7_75t_L g443 ( .A(n_346), .Y(n_443) );
INVx1_ASAP7_75t_L g464 ( .A(n_347), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OAI21xp5_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_357), .B(n_366), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
AND2x2_ASAP7_75t_L g497 ( .A(n_353), .B(n_430), .Y(n_497) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g465 ( .A(n_354), .B(n_425), .Y(n_465) );
AOI32xp33_ASAP7_75t_L g378 ( .A1(n_355), .A2(n_361), .A3(n_379), .B1(n_381), .B2(n_382), .Y(n_378) );
AOI322xp5_ASAP7_75t_L g480 ( .A1(n_355), .A2(n_387), .A3(n_470), .B1(n_481), .B2(n_482), .C1(n_483), .C2(n_485), .Y(n_480) );
INVx2_ASAP7_75t_L g360 ( .A(n_356), .Y(n_360) );
INVx1_ASAP7_75t_L g470 ( .A(n_356), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_361), .B1(n_362), .B2(n_363), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_358), .B(n_364), .Y(n_413) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_359), .B(n_425), .Y(n_475) );
INVx1_ASAP7_75t_L g362 ( .A(n_360), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_360), .B(n_389), .Y(n_479) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_368), .B(n_463), .Y(n_462) );
OAI221xp5_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_371), .B1(n_374), .B2(n_377), .C(n_378), .Y(n_369) );
OR2x2_ASAP7_75t_L g390 ( .A(n_371), .B(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g399 ( .A(n_371), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g424 ( .A(n_372), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g428 ( .A(n_382), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_388), .B1(n_390), .B2(n_392), .C(n_393), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_386), .A2(n_417), .B1(n_421), .B2(n_422), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_387), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g492 ( .A(n_387), .Y(n_492) );
INVx1_ASAP7_75t_L g486 ( .A(n_389), .Y(n_486) );
INVx1_ASAP7_75t_SL g421 ( .A(n_390), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_392), .B(n_420), .Y(n_482) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_397), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g463 ( .A(n_397), .Y(n_463) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
OAI221xp5_ASAP7_75t_SL g401 ( .A1(n_402), .A2(n_406), .B1(n_408), .B2(n_409), .C(n_411), .Y(n_401) );
NOR2xp33_ASAP7_75t_SL g402 ( .A(n_403), .B(n_405), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_403), .A2(n_421), .B1(n_467), .B2(n_468), .Y(n_466) );
CKINVDCx14_ASAP7_75t_R g406 ( .A(n_407), .Y(n_406) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_408), .A2(n_486), .B(n_487), .Y(n_485) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR3xp33_ASAP7_75t_SL g414 ( .A(n_415), .B(n_447), .C(n_471), .Y(n_414) );
NAND4xp25_ASAP7_75t_L g415 ( .A(n_416), .B(n_423), .C(n_431), .D(n_438), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g494 ( .A(n_419), .Y(n_494) );
INVx3_ASAP7_75t_SL g488 ( .A(n_420), .Y(n_488) );
OR2x2_ASAP7_75t_L g493 ( .A(n_420), .B(n_494), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_428), .B2(n_430), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_425), .B(n_443), .Y(n_484) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI21xp5_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_433), .B(n_435), .Y(n_431) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_444), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI211xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_450), .B(n_453), .C(n_466), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g481 ( .A(n_452), .Y(n_481) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_458), .B1(n_459), .B2(n_462), .C1(n_464), .C2(n_465), .Y(n_453) );
INVxp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND4xp25_ASAP7_75t_SL g490 ( .A(n_463), .B(n_491), .C(n_492), .D(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND3xp33_ASAP7_75t_SL g471 ( .A(n_472), .B(n_480), .C(n_489), .Y(n_471) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_517), .Y(n_516) );
endmodule