module real_aes_162_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g532 ( .A(n_0), .B(n_229), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_1), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g163 ( .A(n_2), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_3), .B(n_535), .Y(n_554) );
NAND2xp33_ASAP7_75t_SL g525 ( .A(n_4), .B(n_184), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_5), .B(n_197), .Y(n_220) );
INVx1_ASAP7_75t_L g517 ( .A(n_6), .Y(n_517) );
INVx1_ASAP7_75t_L g254 ( .A(n_7), .Y(n_254) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_8), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_9), .Y(n_271) );
AND2x2_ASAP7_75t_L g552 ( .A(n_10), .B(n_153), .Y(n_552) );
INVx2_ASAP7_75t_L g154 ( .A(n_11), .Y(n_154) );
NOR3xp33_ASAP7_75t_L g114 ( .A(n_12), .B(n_115), .C(n_117), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_12), .Y(n_128) );
INVx1_ASAP7_75t_L g230 ( .A(n_13), .Y(n_230) );
AOI221x1_ASAP7_75t_L g520 ( .A1(n_14), .A2(n_186), .B1(n_521), .B2(n_523), .C(n_524), .Y(n_520) );
OAI22xp5_ASAP7_75t_SL g806 ( .A1(n_14), .A2(n_58), .B1(n_807), .B2(n_808), .Y(n_806) );
INVxp67_ASAP7_75t_L g808 ( .A(n_14), .Y(n_808) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_15), .B(n_535), .Y(n_588) );
INVx1_ASAP7_75t_L g112 ( .A(n_16), .Y(n_112) );
INVx1_ASAP7_75t_L g227 ( .A(n_17), .Y(n_227) );
INVx1_ASAP7_75t_SL g175 ( .A(n_18), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_19), .B(n_178), .Y(n_200) );
AOI33xp33_ASAP7_75t_L g245 ( .A1(n_20), .A2(n_48), .A3(n_160), .B1(n_171), .B2(n_246), .B3(n_247), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_21), .A2(n_523), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_22), .B(n_229), .Y(n_557) );
AOI221xp5_ASAP7_75t_SL g597 ( .A1(n_23), .A2(n_39), .B1(n_523), .B2(n_535), .C(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g264 ( .A(n_24), .Y(n_264) );
OR2x2_ASAP7_75t_L g155 ( .A(n_25), .B(n_93), .Y(n_155) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_25), .A2(n_93), .B(n_154), .Y(n_188) );
INVxp67_ASAP7_75t_L g519 ( .A(n_26), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_27), .B(n_232), .Y(n_592) );
AND2x2_ASAP7_75t_L g546 ( .A(n_28), .B(n_152), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_29), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_30), .B(n_126), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_31), .A2(n_523), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_32), .B(n_232), .Y(n_599) );
AND2x2_ASAP7_75t_L g165 ( .A(n_33), .B(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g170 ( .A(n_33), .Y(n_170) );
AND2x2_ASAP7_75t_L g184 ( .A(n_33), .B(n_163), .Y(n_184) );
INVxp67_ASAP7_75t_L g117 ( .A(n_34), .Y(n_117) );
OR2x6_ASAP7_75t_L g129 ( .A(n_34), .B(n_111), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_35), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_36), .B(n_158), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_37), .A2(n_187), .B1(n_193), .B2(n_197), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_38), .B(n_202), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_40), .A2(n_84), .B1(n_168), .B2(n_523), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_41), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_42), .B(n_229), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_43), .B(n_204), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_44), .B(n_178), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_45), .Y(n_196) );
AND2x2_ASAP7_75t_L g536 ( .A(n_46), .B(n_152), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_47), .B(n_152), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_49), .B(n_178), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_50), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_50), .A2(n_63), .B1(n_443), .B2(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_51), .B(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g161 ( .A(n_52), .Y(n_161) );
INVx1_ASAP7_75t_L g180 ( .A(n_52), .Y(n_180) );
AOI22x1_ASAP7_75t_L g133 ( .A1(n_53), .A2(n_134), .B1(n_135), .B2(n_136), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_53), .Y(n_134) );
AND2x2_ASAP7_75t_L g296 ( .A(n_54), .B(n_152), .Y(n_296) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_55), .A2(n_77), .B1(n_158), .B2(n_168), .C(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_56), .B(n_158), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_57), .B(n_535), .Y(n_545) );
INVx1_ASAP7_75t_L g807 ( .A(n_58), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_59), .B(n_187), .Y(n_273) );
AOI21xp5_ASAP7_75t_SL g209 ( .A1(n_60), .A2(n_168), .B(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g573 ( .A(n_61), .B(n_152), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_62), .B(n_232), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_63), .Y(n_819) );
INVx1_ASAP7_75t_L g223 ( .A(n_64), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_65), .B(n_229), .Y(n_571) );
AND2x2_ASAP7_75t_SL g593 ( .A(n_66), .B(n_153), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_67), .A2(n_523), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g294 ( .A(n_68), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_69), .B(n_232), .Y(n_558) );
AND2x2_ASAP7_75t_SL g565 ( .A(n_70), .B(n_204), .Y(n_565) );
XOR2xp5_ASAP7_75t_L g132 ( .A(n_71), .B(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_72), .A2(n_104), .B1(n_137), .B2(n_138), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_72), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_73), .A2(n_168), .B(n_293), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_74), .A2(n_817), .B1(n_818), .B2(n_820), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_74), .Y(n_817) );
INVx1_ASAP7_75t_L g166 ( .A(n_75), .Y(n_166) );
INVx1_ASAP7_75t_L g182 ( .A(n_75), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_76), .B(n_158), .Y(n_248) );
AND2x2_ASAP7_75t_L g185 ( .A(n_78), .B(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g224 ( .A(n_79), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_80), .A2(n_168), .B(n_174), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_81), .A2(n_168), .B(n_199), .C(n_203), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_82), .A2(n_87), .B1(n_158), .B2(n_535), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_83), .B(n_535), .Y(n_572) );
INVx1_ASAP7_75t_L g113 ( .A(n_85), .Y(n_113) );
AND2x2_ASAP7_75t_SL g207 ( .A(n_86), .B(n_186), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_88), .A2(n_168), .B1(n_243), .B2(n_244), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_89), .B(n_229), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_90), .B(n_229), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_91), .A2(n_106), .B1(n_118), .B2(n_829), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_92), .A2(n_523), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g211 ( .A(n_94), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_95), .B(n_232), .Y(n_570) );
AND2x2_ASAP7_75t_L g249 ( .A(n_96), .B(n_186), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_97), .A2(n_262), .B(n_263), .C(n_265), .Y(n_261) );
INVxp67_ASAP7_75t_L g522 ( .A(n_98), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_99), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_100), .B(n_232), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_101), .A2(n_523), .B(n_590), .Y(n_589) );
BUFx2_ASAP7_75t_L g123 ( .A(n_102), .Y(n_123) );
INVx1_ASAP7_75t_SL g804 ( .A(n_102), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_103), .B(n_178), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_104), .Y(n_138) );
BUFx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_SL g829 ( .A(n_109), .Y(n_829) );
AND2x2_ASAP7_75t_SL g109 ( .A(n_110), .B(n_114), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_802), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_130), .Y(n_124) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x6_ASAP7_75t_SL g507 ( .A(n_128), .B(n_129), .Y(n_507) );
OR2x6_ASAP7_75t_SL g798 ( .A(n_128), .B(n_799), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_128), .B(n_799), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_129), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B1(n_139), .B2(n_800), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OAI22x1_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_506), .B1(n_508), .B2(n_796), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_141), .A2(n_506), .B1(n_509), .B2(n_801), .Y(n_800) );
AND3x1_ASAP7_75t_L g141 ( .A(n_142), .B(n_500), .C(n_503), .Y(n_141) );
NAND5xp2_ASAP7_75t_L g142 ( .A(n_143), .B(n_400), .C(n_430), .D(n_444), .E(n_470), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OAI21xp33_ASAP7_75t_L g500 ( .A1(n_144), .A2(n_443), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g813 ( .A(n_144), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_349), .Y(n_144) );
NOR3xp33_ASAP7_75t_SL g145 ( .A(n_146), .B(n_297), .C(n_331), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_214), .B(n_236), .C(n_275), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_189), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_149), .B(n_287), .Y(n_352) );
AND2x2_ASAP7_75t_L g439 ( .A(n_149), .B(n_217), .Y(n_439) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OR2x2_ASAP7_75t_L g235 ( .A(n_150), .B(n_206), .Y(n_235) );
INVx1_ASAP7_75t_L g277 ( .A(n_150), .Y(n_277) );
INVx2_ASAP7_75t_L g282 ( .A(n_150), .Y(n_282) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_150), .Y(n_310) );
INVx1_ASAP7_75t_L g324 ( .A(n_150), .Y(n_324) );
AND2x2_ASAP7_75t_L g328 ( .A(n_150), .B(n_219), .Y(n_328) );
AND2x2_ASAP7_75t_L g409 ( .A(n_150), .B(n_218), .Y(n_409) );
AO21x2_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_156), .B(n_185), .Y(n_150) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_151), .A2(n_540), .B(n_546), .Y(n_539) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_151), .A2(n_567), .B(n_573), .Y(n_566) );
AO21x2_ASAP7_75t_L g604 ( .A1(n_151), .A2(n_540), .B(n_546), .Y(n_604) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_152), .Y(n_151) );
OA21x2_ASAP7_75t_L g596 ( .A1(n_152), .A2(n_597), .B(n_601), .Y(n_596) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_154), .B(n_155), .Y(n_153) );
AND2x4_ASAP7_75t_L g197 ( .A(n_154), .B(n_155), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_167), .Y(n_156) );
INVx1_ASAP7_75t_L g274 ( .A(n_158), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_158), .A2(n_168), .B1(n_516), .B2(n_518), .Y(n_515) );
AND2x4_ASAP7_75t_L g158 ( .A(n_159), .B(n_164), .Y(n_158) );
INVx1_ASAP7_75t_L g194 ( .A(n_159), .Y(n_194) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_162), .Y(n_159) );
OR2x6_ASAP7_75t_L g176 ( .A(n_160), .B(n_172), .Y(n_176) );
INVxp33_ASAP7_75t_L g246 ( .A(n_160), .Y(n_246) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g173 ( .A(n_161), .B(n_163), .Y(n_173) );
AND2x4_ASAP7_75t_L g232 ( .A(n_161), .B(n_181), .Y(n_232) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g195 ( .A(n_164), .Y(n_195) );
BUFx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x6_ASAP7_75t_L g523 ( .A(n_165), .B(n_173), .Y(n_523) );
INVx2_ASAP7_75t_L g172 ( .A(n_166), .Y(n_172) );
AND2x6_ASAP7_75t_L g229 ( .A(n_166), .B(n_179), .Y(n_229) );
INVxp67_ASAP7_75t_L g272 ( .A(n_168), .Y(n_272) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_173), .Y(n_168) );
NOR2x1p5_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
INVx1_ASAP7_75t_L g247 ( .A(n_171), .Y(n_247) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_183), .Y(n_174) );
INVx2_ASAP7_75t_L g202 ( .A(n_176), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_176), .A2(n_183), .B(n_211), .C(n_212), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_176), .A2(n_223), .B1(n_224), .B2(n_225), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_SL g253 ( .A1(n_176), .A2(n_183), .B(n_254), .C(n_255), .Y(n_253) );
INVxp67_ASAP7_75t_L g262 ( .A(n_176), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g293 ( .A1(n_176), .A2(n_183), .B(n_294), .C(n_295), .Y(n_293) );
INVx1_ASAP7_75t_L g225 ( .A(n_178), .Y(n_225) );
AND2x4_ASAP7_75t_L g535 ( .A(n_178), .B(n_184), .Y(n_535) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_181), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_183), .A2(n_200), .B(n_201), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_183), .B(n_197), .Y(n_233) );
INVx1_ASAP7_75t_L g243 ( .A(n_183), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_183), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_183), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_183), .A2(n_557), .B(n_558), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_183), .A2(n_570), .B(n_571), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_183), .A2(n_591), .B(n_592), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_183), .A2(n_599), .B(n_600), .Y(n_598) );
INVx5_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_184), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_186), .A2(n_261), .B1(n_266), .B2(n_267), .Y(n_260) );
INVx3_ASAP7_75t_L g267 ( .A(n_186), .Y(n_267) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_187), .B(n_270), .Y(n_269) );
AOI21x1_ASAP7_75t_L g528 ( .A1(n_187), .A2(n_529), .B(n_536), .Y(n_528) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
BUFx4f_ASAP7_75t_L g204 ( .A(n_188), .Y(n_204) );
AND2x4_ASAP7_75t_SL g189 ( .A(n_190), .B(n_205), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g234 ( .A(n_191), .Y(n_234) );
AND2x2_ASAP7_75t_L g278 ( .A(n_191), .B(n_219), .Y(n_278) );
AND2x2_ASAP7_75t_L g299 ( .A(n_191), .B(n_206), .Y(n_299) );
INVx1_ASAP7_75t_L g322 ( .A(n_191), .Y(n_322) );
AND2x4_ASAP7_75t_L g389 ( .A(n_191), .B(n_218), .Y(n_389) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_198), .Y(n_191) );
NOR3xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .C(n_196), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_197), .A2(n_209), .B(n_213), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_197), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_197), .B(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_197), .B(n_522), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_197), .B(n_225), .C(n_525), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_197), .A2(n_554), .B(n_555), .Y(n_553) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_203), .A2(n_241), .B(n_249), .Y(n_240) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_203), .A2(n_241), .B(n_249), .Y(n_304) );
AOI21x1_ASAP7_75t_L g561 ( .A1(n_203), .A2(n_562), .B(n_565), .Y(n_561) );
INVx2_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_204), .A2(n_252), .B(n_256), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_204), .A2(n_588), .B(n_589), .Y(n_587) );
AND2x4_ASAP7_75t_L g405 ( .A(n_205), .B(n_322), .Y(n_405) );
OR2x2_ASAP7_75t_L g446 ( .A(n_205), .B(n_447), .Y(n_446) );
NOR2xp67_ASAP7_75t_SL g465 ( .A(n_205), .B(n_338), .Y(n_465) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_205), .B(n_397), .Y(n_483) );
INVx4_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2x1_ASAP7_75t_SL g283 ( .A(n_206), .B(n_219), .Y(n_283) );
AND2x4_ASAP7_75t_L g321 ( .A(n_206), .B(n_322), .Y(n_321) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_206), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_206), .B(n_281), .Y(n_359) );
INVx2_ASAP7_75t_L g373 ( .A(n_206), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_206), .B(n_325), .Y(n_395) );
AND2x2_ASAP7_75t_L g487 ( .A(n_206), .B(n_345), .Y(n_487) );
OR2x6_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NOR2x1_ASAP7_75t_L g215 ( .A(n_216), .B(n_235), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_217), .B(n_324), .Y(n_338) );
AND2x2_ASAP7_75t_SL g347 ( .A(n_217), .B(n_327), .Y(n_347) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_234), .Y(n_217) );
INVx1_ASAP7_75t_L g325 ( .A(n_218), .Y(n_325) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g345 ( .A(n_219), .Y(n_345) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_226), .B(n_233), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_225), .B(n_264), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B1(n_230), .B2(n_231), .Y(n_226) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVxp67_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g378 ( .A(n_234), .Y(n_378) );
INVx2_ASAP7_75t_SL g423 ( .A(n_235), .Y(n_423) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_257), .Y(n_237) );
NAND2x1p5_ASAP7_75t_L g332 ( .A(n_238), .B(n_333), .Y(n_332) );
BUFx2_ASAP7_75t_L g369 ( .A(n_238), .Y(n_369) );
AND2x2_ASAP7_75t_L g493 ( .A(n_238), .B(n_318), .Y(n_493) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_250), .Y(n_238) );
AND2x4_ASAP7_75t_L g306 ( .A(n_239), .B(n_288), .Y(n_306) );
INVx1_ASAP7_75t_L g317 ( .A(n_239), .Y(n_317) );
AND2x2_ASAP7_75t_L g348 ( .A(n_239), .B(n_303), .Y(n_348) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_240), .B(n_251), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_240), .B(n_289), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_242), .B(n_248), .Y(n_241) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVxp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g286 ( .A(n_251), .Y(n_286) );
AND2x4_ASAP7_75t_L g354 ( .A(n_251), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g366 ( .A(n_251), .Y(n_366) );
INVx1_ASAP7_75t_L g408 ( .A(n_251), .Y(n_408) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_251), .Y(n_420) );
AND2x2_ASAP7_75t_L g436 ( .A(n_251), .B(n_259), .Y(n_436) );
BUFx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g383 ( .A(n_258), .B(n_341), .Y(n_383) );
INVx1_ASAP7_75t_SL g385 ( .A(n_258), .Y(n_385) );
AND2x2_ASAP7_75t_L g406 ( .A(n_258), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g285 ( .A(n_259), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g313 ( .A(n_259), .Y(n_313) );
INVx2_ASAP7_75t_L g319 ( .A(n_259), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_259), .B(n_289), .Y(n_334) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_268), .Y(n_259) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_267), .A2(n_290), .B(n_296), .Y(n_289) );
AO21x2_ASAP7_75t_L g303 ( .A1(n_267), .A2(n_290), .B(n_296), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .B1(n_273), .B2(n_274), .Y(n_268) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_279), .B(n_284), .Y(n_275) );
INVx1_ASAP7_75t_L g415 ( .A(n_276), .Y(n_415) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx2_ASAP7_75t_L g335 ( .A(n_278), .Y(n_335) );
AND2x2_ASAP7_75t_L g391 ( .A(n_278), .B(n_327), .Y(n_391) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g305 ( .A(n_280), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_280), .B(n_321), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_280), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g412 ( .A(n_280), .B(n_405), .Y(n_412) );
AND2x2_ASAP7_75t_L g486 ( .A(n_280), .B(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_281), .Y(n_474) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_282), .Y(n_394) );
AND2x2_ASAP7_75t_L g307 ( .A(n_283), .B(n_308), .Y(n_307) );
OAI21xp33_ASAP7_75t_L g495 ( .A1(n_283), .A2(n_496), .B(n_498), .Y(n_495) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx3_ASAP7_75t_L g381 ( .A(n_285), .Y(n_381) );
NAND2x1_ASAP7_75t_SL g425 ( .A(n_285), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g428 ( .A(n_285), .B(n_306), .Y(n_428) );
AND2x2_ASAP7_75t_L g340 ( .A(n_287), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g477 ( .A(n_287), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g488 ( .A(n_287), .B(n_436), .Y(n_488) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2x1p5_ASAP7_75t_L g364 ( .A(n_288), .B(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g419 ( .A(n_289), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
OAI21xp5_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_311), .B(n_314), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B1(n_306), .B2(n_307), .Y(n_298) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_299), .Y(n_356) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_305), .Y(n_300) );
AND2x2_ASAP7_75t_L g329 ( .A(n_301), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g435 ( .A(n_301), .B(n_436), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_301), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_301), .B(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g318 ( .A(n_303), .B(n_319), .Y(n_318) );
NOR2xp67_ASAP7_75t_L g399 ( .A(n_303), .B(n_319), .Y(n_399) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_303), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g355 ( .A(n_304), .Y(n_355) );
AND2x2_ASAP7_75t_L g363 ( .A(n_304), .B(n_319), .Y(n_363) );
INVx1_ASAP7_75t_L g426 ( .A(n_304), .Y(n_426) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2x1_ASAP7_75t_L g344 ( .A(n_309), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g456 ( .A(n_312), .B(n_341), .Y(n_456) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g330 ( .A(n_313), .Y(n_330) );
AND2x2_ASAP7_75t_L g353 ( .A(n_313), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g441 ( .A(n_313), .B(n_348), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_320), .B1(n_326), .B2(n_329), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g449 ( .A(n_316), .B(n_450), .Y(n_449) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g479 ( .A(n_319), .B(n_366), .Y(n_479) );
AND2x2_ASAP7_75t_SL g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx2_ASAP7_75t_L g346 ( .A(n_321), .Y(n_346) );
OAI21xp33_ASAP7_75t_SL g492 ( .A1(n_321), .A2(n_493), .B(n_494), .Y(n_492) );
AND2x4_ASAP7_75t_SL g323 ( .A(n_324), .B(n_325), .Y(n_323) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_324), .Y(n_482) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_SL g424 ( .A1(n_327), .A2(n_425), .B(n_427), .C(n_429), .Y(n_424) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_328), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g429 ( .A(n_328), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_328), .B(n_405), .Y(n_469) );
INVx1_ASAP7_75t_SL g336 ( .A(n_329), .Y(n_336) );
AND2x2_ASAP7_75t_L g417 ( .A(n_330), .B(n_354), .Y(n_417) );
INVx1_ASAP7_75t_L g462 ( .A(n_330), .Y(n_462) );
OAI221xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .B1(n_336), .B2(n_337), .C(n_339), .Y(n_331) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_332), .Y(n_451) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g499 ( .A(n_334), .B(n_342), .Y(n_499) );
OR2x2_ASAP7_75t_L g358 ( .A(n_335), .B(n_359), .Y(n_358) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_335), .B(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_335), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g497 ( .A(n_335), .B(n_394), .Y(n_497) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI32xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_343), .A3(n_346), .B1(n_347), .B2(n_348), .Y(n_339) );
INVx1_ASAP7_75t_L g360 ( .A(n_341), .Y(n_360) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_343), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g455 ( .A(n_344), .Y(n_455) );
OAI22xp33_ASAP7_75t_SL g437 ( .A1(n_346), .A2(n_438), .B1(n_440), .B2(n_442), .Y(n_437) );
INVx1_ASAP7_75t_L g468 ( .A(n_347), .Y(n_468) );
AOI211x1_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_356), .B(n_357), .C(n_374), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_351), .B(n_436), .Y(n_442) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g398 ( .A(n_354), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g464 ( .A(n_354), .Y(n_464) );
OAI222xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B1(n_361), .B2(n_367), .C1(n_368), .C2(n_370), .Y(n_357) );
INVxp67_ASAP7_75t_L g454 ( .A(n_358), .Y(n_454) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_362), .B(n_447), .Y(n_494) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g410 ( .A(n_363), .B(n_407), .Y(n_410) );
INVx3_ASAP7_75t_L g450 ( .A(n_365), .Y(n_450) );
BUFx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g388 ( .A(n_373), .B(n_389), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_379), .B1(n_382), .B2(n_387), .C(n_390), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_376), .A2(n_433), .B(n_435), .Y(n_432) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g386 ( .A(n_380), .Y(n_386) );
OR2x2_ASAP7_75t_L g490 ( .A(n_381), .B(n_426), .Y(n_490) );
NOR2xp67_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_384), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_387), .A2(n_416), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_388), .A2(n_460), .B(n_467), .Y(n_466) );
INVx4_ASAP7_75t_L g397 ( .A(n_389), .Y(n_397) );
OAI31xp33_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_392), .A3(n_396), .B(n_398), .Y(n_390) );
INVx1_ASAP7_75t_L g448 ( .A(n_392), .Y(n_448) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g422 ( .A(n_397), .Y(n_422) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_413), .Y(n_400) );
NAND4xp25_ASAP7_75t_L g501 ( .A(n_401), .B(n_413), .C(n_432), .D(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_411), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_406), .B1(n_409), .B2(n_410), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g473 ( .A(n_405), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_406), .B(n_426), .Y(n_434) );
INVx1_ASAP7_75t_SL g447 ( .A(n_409), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_424), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_418), .B2(n_421), .Y(n_414) );
INVx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2x1_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_423), .A2(n_486), .B1(n_488), .B2(n_489), .Y(n_485) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NOR3xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_437), .C(n_443), .Y(n_430) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g502 ( .A(n_437), .Y(n_502) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI21xp33_ASAP7_75t_L g503 ( .A1(n_443), .A2(n_504), .B(n_505), .Y(n_503) );
INVxp33_ASAP7_75t_L g504 ( .A(n_444), .Y(n_504) );
AND2x2_ASAP7_75t_L g812 ( .A(n_444), .B(n_470), .Y(n_812) );
NOR2xp67_ASAP7_75t_L g444 ( .A(n_445), .B(n_452), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B1(n_449), .B2(n_451), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_449), .A2(n_472), .B(n_475), .Y(n_471) );
INVx2_ASAP7_75t_L g459 ( .A(n_450), .Y(n_459) );
NAND3xp33_ASAP7_75t_SL g452 ( .A(n_453), .B(n_457), .C(n_466), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_460), .B1(n_463), .B2(n_465), .Y(n_457) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVxp33_ASAP7_75t_SL g505 ( .A(n_470), .Y(n_505) );
NOR3x1_ASAP7_75t_L g470 ( .A(n_471), .B(n_484), .C(n_491), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_480), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_492), .B(n_495), .Y(n_491) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g814 ( .A(n_501), .Y(n_814) );
CKINVDCx11_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_673), .Y(n_509) );
NOR4xp25_ASAP7_75t_L g510 ( .A(n_511), .B(n_616), .C(n_655), .D(n_662), .Y(n_510) );
OAI221xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_537), .B1(n_574), .B2(n_583), .C(n_602), .Y(n_511) );
OR2x2_ASAP7_75t_L g746 ( .A(n_512), .B(n_608), .Y(n_746) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g661 ( .A(n_513), .B(n_586), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_513), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_SL g726 ( .A(n_513), .B(n_727), .Y(n_726) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_526), .Y(n_513) );
AND2x4_ASAP7_75t_SL g585 ( .A(n_514), .B(n_586), .Y(n_585) );
INVx3_ASAP7_75t_L g607 ( .A(n_514), .Y(n_607) );
AND2x2_ASAP7_75t_L g642 ( .A(n_514), .B(n_615), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_514), .B(n_527), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_514), .B(n_609), .Y(n_694) );
OR2x2_ASAP7_75t_L g772 ( .A(n_514), .B(n_586), .Y(n_772) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_520), .Y(n_514) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g594 ( .A(n_527), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_527), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g620 ( .A(n_527), .Y(n_620) );
OR2x2_ASAP7_75t_L g625 ( .A(n_527), .B(n_609), .Y(n_625) );
AND2x2_ASAP7_75t_L g638 ( .A(n_527), .B(n_596), .Y(n_638) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_527), .Y(n_641) );
INVx1_ASAP7_75t_L g653 ( .A(n_527), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_527), .B(n_607), .Y(n_718) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_534), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_538), .B(n_547), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g582 ( .A(n_539), .B(n_566), .Y(n_582) );
AND2x4_ASAP7_75t_L g612 ( .A(n_539), .B(n_551), .Y(n_612) );
INVx2_ASAP7_75t_L g646 ( .A(n_539), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_539), .B(n_566), .Y(n_704) );
AND2x2_ASAP7_75t_L g751 ( .A(n_539), .B(n_580), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_545), .Y(n_540) );
AOI222xp33_ASAP7_75t_L g739 ( .A1(n_547), .A2(n_611), .B1(n_654), .B2(n_714), .C1(n_740), .C2(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_559), .Y(n_548) );
AND2x2_ASAP7_75t_L g658 ( .A(n_549), .B(n_578), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_549), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g787 ( .A(n_549), .B(n_627), .Y(n_787) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_550), .A2(n_618), .B(n_622), .Y(n_617) );
AND2x2_ASAP7_75t_L g698 ( .A(n_550), .B(n_581), .Y(n_698) );
OR2x2_ASAP7_75t_L g723 ( .A(n_550), .B(n_582), .Y(n_723) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx5_ASAP7_75t_L g577 ( .A(n_551), .Y(n_577) );
AND2x2_ASAP7_75t_L g664 ( .A(n_551), .B(n_646), .Y(n_664) );
AND2x2_ASAP7_75t_L g690 ( .A(n_551), .B(n_566), .Y(n_690) );
OR2x2_ASAP7_75t_L g693 ( .A(n_551), .B(n_580), .Y(n_693) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_551), .Y(n_711) );
AND2x4_ASAP7_75t_SL g768 ( .A(n_551), .B(n_645), .Y(n_768) );
OR2x2_ASAP7_75t_L g777 ( .A(n_551), .B(n_604), .Y(n_777) );
OR2x6_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g610 ( .A(n_559), .Y(n_610) );
AOI221xp5_ASAP7_75t_SL g728 ( .A1(n_559), .A2(n_612), .B1(n_729), .B2(n_731), .C(n_732), .Y(n_728) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_566), .Y(n_559) );
OR2x2_ASAP7_75t_L g667 ( .A(n_560), .B(n_637), .Y(n_667) );
OR2x2_ASAP7_75t_L g677 ( .A(n_560), .B(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g703 ( .A(n_560), .B(n_704), .Y(n_703) );
AND2x4_ASAP7_75t_L g709 ( .A(n_560), .B(n_628), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_560), .B(n_692), .Y(n_721) );
INVx2_ASAP7_75t_L g734 ( .A(n_560), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g755 ( .A(n_560), .B(n_612), .Y(n_755) );
AND2x2_ASAP7_75t_L g759 ( .A(n_560), .B(n_581), .Y(n_759) );
AND2x2_ASAP7_75t_L g767 ( .A(n_560), .B(n_768), .Y(n_767) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g580 ( .A(n_561), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_566), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g611 ( .A(n_566), .B(n_580), .Y(n_611) );
INVx2_ASAP7_75t_L g628 ( .A(n_566), .Y(n_628) );
AND2x4_ASAP7_75t_L g645 ( .A(n_566), .B(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_566), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_578), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g757 ( .A(n_576), .B(n_579), .Y(n_757) );
AND2x4_ASAP7_75t_L g603 ( .A(n_577), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g644 ( .A(n_577), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g671 ( .A(n_577), .B(n_611), .Y(n_671) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g775 ( .A(n_579), .B(n_776), .Y(n_775) );
BUFx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g627 ( .A(n_580), .B(n_628), .Y(n_627) );
OAI21xp5_ASAP7_75t_SL g647 ( .A1(n_581), .A2(n_648), .B(n_654), .Y(n_647) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_594), .Y(n_584) );
INVx1_ASAP7_75t_SL g701 ( .A(n_585), .Y(n_701) );
AND2x2_ASAP7_75t_L g731 ( .A(n_585), .B(n_641), .Y(n_731) );
AND2x4_ASAP7_75t_L g742 ( .A(n_585), .B(n_743), .Y(n_742) );
OR2x2_ASAP7_75t_L g608 ( .A(n_586), .B(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g615 ( .A(n_586), .Y(n_615) );
AND2x4_ASAP7_75t_L g621 ( .A(n_586), .B(n_607), .Y(n_621) );
INVx2_ASAP7_75t_L g632 ( .A(n_586), .Y(n_632) );
INVx1_ASAP7_75t_L g681 ( .A(n_586), .Y(n_681) );
OR2x2_ASAP7_75t_L g702 ( .A(n_586), .B(n_686), .Y(n_702) );
OR2x2_ASAP7_75t_L g716 ( .A(n_586), .B(n_596), .Y(n_716) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_586), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_586), .B(n_638), .Y(n_788) );
OR2x6_ASAP7_75t_L g586 ( .A(n_587), .B(n_593), .Y(n_586) );
INVx1_ASAP7_75t_L g633 ( .A(n_594), .Y(n_633) );
AND2x2_ASAP7_75t_L g766 ( .A(n_594), .B(n_632), .Y(n_766) );
AND2x2_ASAP7_75t_L g791 ( .A(n_594), .B(n_621), .Y(n_791) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g609 ( .A(n_596), .Y(n_609) );
BUFx3_ASAP7_75t_L g651 ( .A(n_596), .Y(n_651) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_596), .Y(n_678) );
INVx1_ASAP7_75t_L g687 ( .A(n_596), .Y(n_687) );
AOI33xp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_605), .A3(n_610), .B1(n_611), .B2(n_612), .B3(n_613), .Y(n_602) );
AOI21x1_ASAP7_75t_SL g705 ( .A1(n_603), .A2(n_627), .B(n_689), .Y(n_705) );
INVx2_ASAP7_75t_L g735 ( .A(n_603), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_603), .B(n_734), .Y(n_741) );
AND2x2_ASAP7_75t_L g689 ( .A(n_604), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AND2x2_ASAP7_75t_L g652 ( .A(n_607), .B(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g753 ( .A(n_608), .Y(n_753) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_609), .Y(n_743) );
OAI32xp33_ASAP7_75t_L g792 ( .A1(n_610), .A2(n_612), .A3(n_788), .B1(n_793), .B2(n_795), .Y(n_792) );
AND2x2_ASAP7_75t_L g710 ( .A(n_611), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_SL g700 ( .A(n_612), .Y(n_700) );
AND2x2_ASAP7_75t_L g765 ( .A(n_612), .B(n_709), .Y(n_765) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_626), .B1(n_629), .B2(n_643), .C(n_647), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_620), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_621), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_621), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_621), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g670 ( .A(n_625), .Y(n_670) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_634), .C(n_639), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g732 ( .A1(n_631), .A2(n_693), .B1(n_733), .B2(n_736), .Y(n_732) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g636 ( .A(n_632), .Y(n_636) );
NOR2x1p5_ASAP7_75t_L g650 ( .A(n_632), .B(n_651), .Y(n_650) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_632), .Y(n_672) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI322xp33_ASAP7_75t_L g699 ( .A1(n_635), .A2(n_677), .A3(n_700), .B1(n_701), .B2(n_702), .C1(n_703), .C2(n_705), .Y(n_699) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g655 ( .A1(n_637), .A2(n_656), .B(n_657), .C(n_659), .Y(n_655) );
OR2x2_ASAP7_75t_L g747 ( .A(n_637), .B(n_701), .Y(n_747) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g654 ( .A(n_638), .B(n_642), .Y(n_654) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g660 ( .A(n_644), .B(n_661), .Y(n_660) );
INVx3_ASAP7_75t_SL g692 ( .A(n_645), .Y(n_692) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_649), .B(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_SL g696 ( .A(n_652), .Y(n_696) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_653), .Y(n_738) );
OR2x6_ASAP7_75t_SL g793 ( .A(n_656), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI211xp5_ASAP7_75t_L g783 ( .A1(n_661), .A2(n_784), .B(n_785), .C(n_792), .Y(n_783) );
O2A1O1Ixp33_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_665), .B(n_668), .C(n_672), .Y(n_662) );
OAI211xp5_ASAP7_75t_SL g674 ( .A1(n_663), .A2(n_675), .B(n_682), .C(n_706), .Y(n_674) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NOR3xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_719), .C(n_763), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_679), .Y(n_675) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_678), .Y(n_770) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g725 ( .A(n_681), .Y(n_725) );
NOR3xp33_ASAP7_75t_SL g682 ( .A(n_683), .B(n_695), .C(n_699), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_688), .B1(n_691), .B2(n_694), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g727 ( .A(n_687), .Y(n_727) );
INVxp67_ASAP7_75t_SL g794 ( .A(n_687), .Y(n_794) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_SL g780 ( .A(n_693), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
OR2x2_ASAP7_75t_L g730 ( .A(n_696), .B(n_716), .Y(n_730) );
OR2x2_ASAP7_75t_L g781 ( .A(n_696), .B(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g779 ( .A(n_704), .Y(n_779) );
OR2x2_ASAP7_75t_L g795 ( .A(n_704), .B(n_734), .Y(n_795) );
OAI21xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_710), .B(n_712), .Y(n_706) );
OAI31xp33_ASAP7_75t_L g720 ( .A1(n_707), .A2(n_721), .A3(n_722), .B(n_724), .Y(n_720) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_717), .Y(n_714) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
AND2x4_ASAP7_75t_L g752 ( .A(n_717), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND4xp25_ASAP7_75t_SL g719 ( .A(n_720), .B(n_728), .C(n_739), .D(n_744), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_727), .Y(n_762) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_748), .B1(n_752), .B2(n_754), .C(n_756), .Y(n_744) );
NAND2xp33_ASAP7_75t_SL g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g789 ( .A(n_748), .Y(n_789) );
AND2x2_ASAP7_75t_SL g748 ( .A(n_749), .B(n_751), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AOI21xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B(n_760), .Y(n_756) );
INVx1_ASAP7_75t_L g784 ( .A(n_758), .Y(n_784) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g763 ( .A(n_764), .B(n_783), .Y(n_763) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B1(n_767), .B2(n_769), .C(n_773), .Y(n_764) );
AND2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
INVx1_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
AOI21xp33_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_778), .B(n_781), .Y(n_773) );
INVxp33_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_788), .B1(n_789), .B2(n_790), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_797), .Y(n_801) );
CKINVDCx11_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
OAI21xp5_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_805), .B(n_826), .Y(n_802) );
INVx2_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
OAI21xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_809), .B(n_821), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g821 ( .A1(n_806), .A2(n_822), .B(n_823), .Y(n_821) );
INVxp67_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g822 ( .A(n_810), .Y(n_822) );
XNOR2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_815), .Y(n_810) );
NAND3x1_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .C(n_814), .Y(n_811) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g820 ( .A(n_818), .Y(n_820) );
CKINVDCx11_ASAP7_75t_R g828 ( .A(n_823), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
BUFx3_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
endmodule