module fake_ariane_1575_n_585 (n_83, n_8, n_56, n_60, n_64, n_90, n_38, n_47, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_92, n_74, n_33, n_19, n_40, n_12, n_53, n_21, n_66, n_71, n_24, n_7, n_49, n_20, n_17, n_50, n_62, n_51, n_76, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_72, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_85, n_6, n_48, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_45, n_11, n_52, n_73, n_77, n_15, n_93, n_23, n_61, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_14, n_88, n_68, n_78, n_39, n_59, n_63, n_16, n_5, n_35, n_54, n_25, n_585);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_90;
input n_38;
input n_47;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_92;
input n_74;
input n_33;
input n_19;
input n_40;
input n_12;
input n_53;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_49;
input n_20;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_72;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_85;
input n_6;
input n_48;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_93;
input n_23;
input n_61;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_14;
input n_88;
input n_68;
input n_78;
input n_39;
input n_59;
input n_63;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_585;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_119;
wire n_124;
wire n_386;
wire n_307;
wire n_516;
wire n_332;
wire n_581;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_133;
wire n_205;
wire n_341;
wire n_109;
wire n_245;
wire n_421;
wire n_96;
wire n_549;
wire n_522;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_103;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_117;
wire n_139;
wire n_524;
wire n_130;
wire n_349;
wire n_391;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_95;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_578;
wire n_152;
wire n_405;
wire n_557;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_309;
wire n_320;
wire n_115;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_481;
wire n_433;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_330;
wire n_400;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_108;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_136;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_104;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_565;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_107;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_94;
wire n_284;
wire n_448;
wire n_249;
wire n_534;
wire n_123;
wire n_212;
wire n_355;
wire n_444;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_475;
wire n_135;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_102;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_125;
wire n_577;
wire n_407;
wire n_254;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_99;
wire n_544;
wire n_216;
wire n_540;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_110;
wire n_304;
wire n_509;
wire n_583;
wire n_306;
wire n_313;
wire n_430;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_98;
wire n_375;
wire n_113;
wire n_114;
wire n_324;
wire n_337;
wire n_437;
wire n_111;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_100;
wire n_132;
wire n_147;
wire n_204;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_105;
wire n_580;
wire n_494;
wire n_131;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_101;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_112;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_118;
wire n_121;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_97;
wire n_408;
wire n_322;
wire n_251;
wire n_506;
wire n_558;
wire n_116;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_573;
wire n_127;
wire n_531;

INVx1_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_5),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_2),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVxp33_ASAP7_75t_SL g100 ( 
.A(n_25),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_72),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_12),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_49),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_6),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVxp33_ASAP7_75t_SL g109 ( 
.A(n_4),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_21),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_65),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_6),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_35),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_33),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_7),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_16),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_3),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_14),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_14),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_43),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_34),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_18),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_46),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_69),
.Y(n_134)
);

INVxp67_ASAP7_75t_SL g135 ( 
.A(n_5),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_12),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_41),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_17),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_15),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_27),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_7),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_48),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_24),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_9),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_11),
.B(n_22),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_55),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_20),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_45),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_9),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_3),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_0),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_53),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_47),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_19),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_32),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_80),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_11),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_4),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_37),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_1),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_40),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_77),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_75),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_56),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_50),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_51),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_67),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_63),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_39),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_1),
.B(n_0),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_2),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_58),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_26),
.Y(n_182)
);

NOR2x1_ASAP7_75t_L g183 ( 
.A(n_116),
.B(n_57),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_8),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_98),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

CKINVDCx11_ASAP7_75t_R g190 ( 
.A(n_129),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_105),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_113),
.B(n_13),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_118),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_29),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_104),
.B(n_30),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_150),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_105),
.A2(n_170),
.B1(n_96),
.B2(n_139),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_136),
.B(n_31),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

BUFx8_ASAP7_75t_L g204 ( 
.A(n_110),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_101),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_101),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_94),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

AND3x2_ASAP7_75t_L g209 ( 
.A(n_110),
.B(n_44),
.C(n_52),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_95),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_103),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_133),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_136),
.B(n_76),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

CKINVDCx11_ASAP7_75t_R g218 ( 
.A(n_117),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_124),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_148),
.B(n_79),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_164),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_148),
.B(n_85),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_99),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_117),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_126),
.B(n_87),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_131),
.A2(n_88),
.B1(n_89),
.B2(n_93),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_100),
.B(n_164),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_124),
.B(n_179),
.Y(n_228)
);

AND2x4_ASAP7_75t_L g229 ( 
.A(n_106),
.B(n_182),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_142),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_160),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_107),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_108),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_135),
.B(n_145),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_111),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_114),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_120),
.B(n_151),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_121),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_131),
.A2(n_165),
.B1(n_144),
.B2(n_161),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_122),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_125),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_127),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_128),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_130),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_171),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_132),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_109),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_138),
.Y(n_249)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_141),
.A2(n_153),
.B(n_178),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_134),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_143),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_147),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_155),
.Y(n_254)
);

NOR2x1_ASAP7_75t_L g255 ( 
.A(n_156),
.B(n_163),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_158),
.Y(n_256)
);

NOR2xp67_ASAP7_75t_L g257 ( 
.A(n_162),
.B(n_168),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_173),
.B(n_177),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_187),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_246),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_184),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_204),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_213),
.B(n_176),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_100),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_195),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_140),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_187),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_240),
.B(n_161),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_197),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_213),
.B(n_175),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_187),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_188),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_190),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_194),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_214),
.B(n_174),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_197),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_201),
.B(n_144),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_197),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_196),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_198),
.Y(n_285)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_197),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_190),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_228),
.B(n_137),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_203),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_228),
.B(n_137),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_218),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_208),
.Y(n_292)
);

NAND2xp33_ASAP7_75t_L g293 ( 
.A(n_197),
.B(n_199),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_234),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_185),
.B(n_112),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_185),
.B(n_216),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_189),
.Y(n_298)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_215),
.Y(n_299)
);

BUFx8_ASAP7_75t_SL g300 ( 
.A(n_205),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_215),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_214),
.B(n_181),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_217),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_217),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_205),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_210),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_250),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_231),
.B(n_109),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_206),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_231),
.B(n_134),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_217),
.Y(n_312)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_204),
.Y(n_313)
);

BUFx4f_ASAP7_75t_L g314 ( 
.A(n_313),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_225),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_313),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_263),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_267),
.A2(n_200),
.B1(n_220),
.B2(n_202),
.Y(n_319)
);

BUFx8_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_293),
.A2(n_258),
.B1(n_192),
.B2(n_221),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_307),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_230),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_222),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_300),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_259),
.Y(n_326)
);

OR2x6_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_193),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_295),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_297),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_270),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_295),
.B(n_229),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_294),
.B(n_234),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_295),
.B(n_235),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_274),
.B(n_229),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_279),
.B(n_219),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_307),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_284),
.B(n_221),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_219),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_296),
.B(n_219),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_302),
.B(n_207),
.Y(n_342)
);

OAI21xp33_ASAP7_75t_L g343 ( 
.A1(n_285),
.A2(n_258),
.B(n_238),
.Y(n_343)
);

O2A1O1Ixp5_ASAP7_75t_L g344 ( 
.A1(n_272),
.A2(n_236),
.B(n_237),
.C(n_242),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_270),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_272),
.B(n_226),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_260),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_266),
.B(n_244),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_293),
.A2(n_192),
.B1(n_250),
.B2(n_255),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_248),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_309),
.B(n_241),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_272),
.B(n_183),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_261),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_308),
.A2(n_241),
.B1(n_252),
.B2(n_253),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_292),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_275),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_312),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_312),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_275),
.Y(n_361)
);

O2A1O1Ixp5_ASAP7_75t_L g362 ( 
.A1(n_282),
.A2(n_245),
.B(n_239),
.C(n_249),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_273),
.B(n_207),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_308),
.Y(n_364)
);

NAND2x1p5_ASAP7_75t_L g365 ( 
.A(n_314),
.B(n_264),
.Y(n_365)
);

OR2x6_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_264),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_322),
.B(n_286),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_315),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_311),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_353),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_327),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_354),
.A2(n_271),
.B1(n_281),
.B2(n_248),
.Y(n_373)
);

NAND3x1_ASAP7_75t_L g374 ( 
.A(n_319),
.B(n_191),
.C(n_300),
.Y(n_374)
);

AO31x2_ASAP7_75t_L g375 ( 
.A1(n_323),
.A2(n_286),
.A3(n_282),
.B(n_303),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_352),
.A2(n_338),
.B(n_336),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_345),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_327),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_350),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_337),
.B(n_280),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_346),
.A2(n_165),
.B1(n_172),
.B2(n_257),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_314),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_317),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_318),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_354),
.B(n_280),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_325),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_326),
.Y(n_389)
);

INVx3_ASAP7_75t_SL g390 ( 
.A(n_347),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_320),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

O2A1O1Ixp33_ASAP7_75t_L g394 ( 
.A1(n_324),
.A2(n_193),
.B(n_243),
.C(n_256),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_346),
.A2(n_172),
.B1(n_273),
.B2(n_283),
.Y(n_395)
);

OR2x6_ASAP7_75t_L g396 ( 
.A(n_316),
.B(n_212),
.Y(n_396)
);

A2O1A1Ixp33_ASAP7_75t_SL g397 ( 
.A1(n_355),
.A2(n_301),
.B(n_283),
.C(n_304),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_334),
.B(n_287),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_329),
.A2(n_244),
.B1(n_211),
.B2(n_254),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_349),
.A2(n_254),
.B1(n_247),
.B2(n_232),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_321),
.B(n_301),
.Y(n_401)
);

BUFx12f_ASAP7_75t_L g402 ( 
.A(n_339),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_344),
.A2(n_283),
.B(n_301),
.Y(n_403)
);

NAND2x1p5_ASAP7_75t_L g404 ( 
.A(n_339),
.B(n_356),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_344),
.A2(n_304),
.B(n_299),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_321),
.A2(n_304),
.B1(n_223),
.B2(n_232),
.Y(n_406)
);

O2A1O1Ixp33_ASAP7_75t_SL g407 ( 
.A1(n_340),
.A2(n_341),
.B(n_348),
.C(n_342),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_333),
.B(n_233),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_343),
.B(n_277),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_332),
.B(n_206),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_357),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_361),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_363),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_358),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_349),
.B(n_277),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_358),
.Y(n_416)
);

O2A1O1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_362),
.A2(n_306),
.B(n_233),
.C(n_223),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_331),
.B(n_224),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_358),
.B(n_291),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_359),
.Y(n_420)
);

INVxp33_ASAP7_75t_L g421 ( 
.A(n_360),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_359),
.Y(n_422)
);

BUFx12f_ASAP7_75t_L g423 ( 
.A(n_359),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_360),
.A2(n_224),
.B1(n_312),
.B2(n_209),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_383),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_368),
.A2(n_218),
.B1(n_291),
.B2(n_331),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_388),
.B(n_331),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_384),
.Y(n_428)
);

CKINVDCx11_ASAP7_75t_R g429 ( 
.A(n_387),
.Y(n_429)
);

NAND3xp33_ASAP7_75t_L g430 ( 
.A(n_369),
.B(n_298),
.C(n_299),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_388),
.B(n_299),
.Y(n_431)
);

OA21x2_ASAP7_75t_L g432 ( 
.A1(n_405),
.A2(n_209),
.B(n_299),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_423),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_376),
.A2(n_297),
.B(n_298),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_382),
.B(n_298),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_386),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_402),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_416),
.Y(n_438)
);

AOI221xp5_ASAP7_75t_L g439 ( 
.A1(n_373),
.A2(n_265),
.B1(n_268),
.B2(n_415),
.C(n_392),
.Y(n_439)
);

O2A1O1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_417),
.A2(n_265),
.B(n_268),
.C(n_394),
.Y(n_440)
);

BUFx8_ASAP7_75t_L g441 ( 
.A(n_391),
.Y(n_441)
);

AO21x2_ASAP7_75t_L g442 ( 
.A1(n_401),
.A2(n_265),
.B(n_268),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_416),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_367),
.A2(n_364),
.B(n_401),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_381),
.A2(n_395),
.B1(n_400),
.B2(n_406),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_408),
.B(n_395),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_370),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_379),
.B(n_398),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_382),
.B(n_366),
.Y(n_449)
);

AO21x2_ASAP7_75t_L g450 ( 
.A1(n_407),
.A2(n_397),
.B(n_385),
.Y(n_450)
);

BUFx8_ASAP7_75t_L g451 ( 
.A(n_371),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_408),
.B(n_406),
.Y(n_452)
);

AOI222xp33_ASAP7_75t_L g453 ( 
.A1(n_372),
.A2(n_378),
.B1(n_393),
.B2(n_409),
.C1(n_410),
.C2(n_418),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_414),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_385),
.A2(n_422),
.B(n_420),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_381),
.B(n_413),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_411),
.Y(n_457)
);

AOI21x1_ASAP7_75t_L g458 ( 
.A1(n_380),
.A2(n_396),
.B(n_375),
.Y(n_458)
);

OAI21x1_ASAP7_75t_SL g459 ( 
.A1(n_419),
.A2(n_424),
.B(n_399),
.Y(n_459)
);

AO31x2_ASAP7_75t_L g460 ( 
.A1(n_375),
.A2(n_424),
.A3(n_389),
.B(n_374),
.Y(n_460)
);

OA21x2_ASAP7_75t_L g461 ( 
.A1(n_375),
.A2(n_412),
.B(n_418),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_404),
.A2(n_421),
.B(n_377),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_366),
.A2(n_396),
.B1(n_390),
.B2(n_365),
.Y(n_463)
);

OAI21x1_ASAP7_75t_L g464 ( 
.A1(n_396),
.A2(n_366),
.B(n_405),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_373),
.A2(n_228),
.B1(n_415),
.B2(n_271),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_383),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_376),
.A2(n_362),
.B(n_344),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_379),
.B(n_370),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_388),
.B(n_382),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_423),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_383),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_368),
.B(n_369),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_383),
.Y(n_474)
);

INVx6_ASAP7_75t_L g475 ( 
.A(n_423),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_368),
.B(n_369),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_373),
.A2(n_228),
.B1(n_415),
.B2(n_271),
.Y(n_477)
);

OA21x2_ASAP7_75t_L g478 ( 
.A1(n_403),
.A2(n_364),
.B(n_405),
.Y(n_478)
);

OA21x2_ASAP7_75t_L g479 ( 
.A1(n_403),
.A2(n_364),
.B(n_405),
.Y(n_479)
);

OA21x2_ASAP7_75t_L g480 ( 
.A1(n_403),
.A2(n_405),
.B(n_401),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_383),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_SL g482 ( 
.A1(n_445),
.A2(n_456),
.B1(n_459),
.B2(n_446),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_425),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_481),
.Y(n_484)
);

OAI211xp5_ASAP7_75t_L g485 ( 
.A1(n_473),
.A2(n_476),
.B(n_426),
.C(n_466),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_475),
.Y(n_486)
);

AOI21xp33_ASAP7_75t_L g487 ( 
.A1(n_445),
.A2(n_466),
.B(n_477),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_428),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_473),
.A2(n_476),
.B1(n_477),
.B2(n_467),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_448),
.B(n_469),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_439),
.A2(n_446),
.B1(n_452),
.B2(n_456),
.Y(n_491)
);

OR2x6_ASAP7_75t_L g492 ( 
.A(n_437),
.B(n_475),
.Y(n_492)
);

AO21x2_ASAP7_75t_L g493 ( 
.A1(n_444),
.A2(n_458),
.B(n_455),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_440),
.A2(n_444),
.B(n_455),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_436),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_L g496 ( 
.A1(n_475),
.A2(n_447),
.B1(n_474),
.B2(n_472),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_449),
.A2(n_470),
.B1(n_453),
.B2(n_463),
.Y(n_497)
);

AOI221xp5_ASAP7_75t_L g498 ( 
.A1(n_465),
.A2(n_439),
.B1(n_463),
.B2(n_457),
.C(n_452),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_454),
.Y(n_499)
);

OAI22xp33_ASAP7_75t_L g500 ( 
.A1(n_433),
.A2(n_471),
.B1(n_437),
.B2(n_454),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_433),
.B(n_471),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_461),
.A2(n_462),
.B1(n_435),
.B2(n_464),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_461),
.A2(n_462),
.B1(n_435),
.B2(n_480),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_480),
.A2(n_442),
.B1(n_431),
.B2(n_427),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_427),
.B(n_443),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_429),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_441),
.Y(n_507)
);

OAI221xp5_ASAP7_75t_L g508 ( 
.A1(n_440),
.A2(n_468),
.B1(n_434),
.B2(n_443),
.C(n_430),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_478),
.A2(n_479),
.B1(n_450),
.B2(n_438),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g510 ( 
.A1(n_478),
.A2(n_479),
.B1(n_450),
.B2(n_438),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_SL g511 ( 
.A1(n_441),
.A2(n_451),
.B1(n_432),
.B2(n_460),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_451),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_499),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_489),
.B(n_460),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_483),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_506),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_490),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_482),
.B(n_460),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_484),
.Y(n_519)
);

AOI221xp5_ASAP7_75t_L g520 ( 
.A1(n_487),
.A2(n_432),
.B1(n_438),
.B2(n_460),
.C(n_485),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_492),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_488),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_495),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_493),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_494),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_486),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_498),
.B(n_497),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_491),
.B(n_505),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_491),
.B(n_503),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_492),
.Y(n_530)
);

NAND4xp25_ASAP7_75t_L g531 ( 
.A(n_513),
.B(n_501),
.C(n_512),
.D(n_486),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_525),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_513),
.Y(n_533)
);

OAI31xp33_ASAP7_75t_L g534 ( 
.A1(n_527),
.A2(n_496),
.A3(n_500),
.B(n_512),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_529),
.B(n_503),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_529),
.B(n_528),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_502),
.Y(n_537)
);

NAND3xp33_ASAP7_75t_L g538 ( 
.A(n_527),
.B(n_510),
.C(n_509),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_525),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_518),
.B(n_502),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_514),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_518),
.B(n_511),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_517),
.B(n_507),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_515),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_515),
.B(n_504),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_514),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_519),
.B(n_504),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_526),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_536),
.B(n_523),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_533),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_534),
.A2(n_520),
.B1(n_522),
.B2(n_523),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_R g552 ( 
.A(n_542),
.B(n_524),
.Y(n_552)
);

NOR2x1_ASAP7_75t_L g553 ( 
.A(n_531),
.B(n_519),
.Y(n_553)
);

AND2x4_ASAP7_75t_SL g554 ( 
.A(n_548),
.B(n_530),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_536),
.B(n_522),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_544),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_541),
.B(n_521),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_555),
.B(n_544),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_550),
.B(n_544),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_554),
.B(n_557),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_549),
.B(n_539),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_553),
.B(n_539),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_554),
.B(n_535),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_556),
.B(n_532),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_561),
.B(n_532),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_564),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_560),
.Y(n_567)
);

AOI32xp33_ASAP7_75t_L g568 ( 
.A1(n_562),
.A2(n_542),
.A3(n_551),
.B1(n_537),
.B2(n_543),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_563),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_558),
.A2(n_552),
.B1(n_551),
.B2(n_537),
.Y(n_570)
);

OAI221xp5_ASAP7_75t_L g571 ( 
.A1(n_559),
.A2(n_552),
.B1(n_492),
.B2(n_538),
.C(n_547),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_567),
.B(n_541),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_566),
.B(n_565),
.Y(n_573)
);

A2O1A1Ixp33_ASAP7_75t_L g574 ( 
.A1(n_568),
.A2(n_540),
.B(n_535),
.C(n_538),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_569),
.B(n_545),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_574),
.A2(n_570),
.B1(n_571),
.B2(n_546),
.Y(n_576)
);

AOI221xp5_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_573),
.B1(n_575),
.B2(n_572),
.C(n_540),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_577),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_578),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_516),
.B(n_567),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_580),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_581),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_582),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_583),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_584),
.A2(n_526),
.B(n_508),
.Y(n_585)
);


endmodule