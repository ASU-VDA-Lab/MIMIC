module real_jpeg_7913_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

AOI21xp33_ASAP7_75t_L g28 ( 
.A1(n_3),
.A2(n_27),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_3),
.B(n_60),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_3),
.A2(n_25),
.B1(n_30),
.B2(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_3),
.B(n_49),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_3),
.A2(n_52),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_3),
.B(n_52),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_3),
.A2(n_38),
.B1(n_43),
.B2(n_135),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_3),
.A2(n_49),
.B(n_104),
.Y(n_157)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

BUFx6f_ASAP7_75t_SL g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_9),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_73),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_29),
.B1(n_49),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_10),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_85),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_85),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_11),
.A2(n_29),
.B1(n_49),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_11),
.A2(n_30),
.B1(n_56),
.B2(n_91),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_56),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_56),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_14),
.A2(n_29),
.B1(n_49),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_58),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_58),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_15),
.A2(n_36),
.B1(n_37),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_15),
.A2(n_52),
.B1(n_53),
.B2(n_64),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_111),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_110),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_93),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_20),
.B(n_93),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_67),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_44),
.B1(n_65),
.B2(n_66),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.C(n_30),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_25),
.B(n_78),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_25),
.B(n_43),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_25),
.B(n_51),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_49),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_26),
.A2(n_30),
.B(n_61),
.C(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_26),
.B(n_30),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_34),
.A2(n_39),
.B1(n_40),
.B2(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_36),
.A2(n_37),
.B1(n_76),
.B2(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_36),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_37),
.B(n_79),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_37),
.B(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_38),
.A2(n_43),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_38),
.A2(n_43),
.B1(n_118),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_38),
.A2(n_43),
.B1(n_108),
.B2(n_120),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_39),
.A2(n_40),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_59),
.C(n_62),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_45),
.A2(n_46),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_51),
.B1(n_55),
.B2(n_57),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_51),
.B1(n_57),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_47),
.A2(n_51),
.B1(n_55),
.B2(n_157),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_76),
.B(n_77),
.C(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_52),
.B(n_54),
.Y(n_105)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_53),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_62),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_87),
.B1(n_90),
.B2(n_92),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_63),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_86),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_82),
.B2(n_83),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_80),
.B2(n_81),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_75),
.B1(n_78),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_78),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_75),
.A2(n_78),
.B1(n_126),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_75),
.A2(n_78),
.B1(n_99),
.B2(n_149),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_76),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.C(n_100),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_94),
.A2(n_95),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_98),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_102),
.B(n_107),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_160),
.B(n_166),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_152),
.B(n_159),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_143),
.B(n_151),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_132),
.B(n_142),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_121),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_127),
.B2(n_131),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_131),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_125),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_127),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_137),
.B(n_141),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_136),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_144),
.B(n_145),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_148),
.C(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_153),
.B(n_154),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.CI(n_158),
.CON(n_154),
.SN(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);


endmodule