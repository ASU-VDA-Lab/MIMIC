module fake_jpeg_7271_n_95 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_95);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_95;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_25),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_26),
.Y(n_30)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_19),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_26),
.B1(n_24),
.B2(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_18),
.Y(n_28)
);

AND2x6_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_18),
.B(n_13),
.C(n_25),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_10),
.B1(n_33),
.B2(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_29),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_20),
.B(n_21),
.C(n_11),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_26),
.B1(n_33),
.B2(n_32),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_19),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx11_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_48),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_20),
.Y(n_50)
);

XOR2x2_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_53),
.Y(n_60)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_55),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_19),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_46),
.C(n_52),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_62),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_42),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_50),
.C(n_53),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_72),
.C(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_23),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_63),
.B(n_58),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_35),
.B(n_10),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_45),
.C(n_40),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_75),
.C(n_76),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_24),
.C(n_12),
.Y(n_77)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_16),
.B1(n_12),
.B2(n_15),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_79),
.B1(n_16),
.B2(n_12),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_7),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_71),
.B(n_72),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_75),
.B(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_84),
.Y(n_86)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_82),
.B(n_87),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_15),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_88),
.Y(n_91)
);

AOI322xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_16),
.A3(n_8),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_1),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_82),
.B1(n_8),
.B2(n_5),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_4),
.Y(n_93)
);

OAI21x1_ASAP7_75t_SL g92 ( 
.A1(n_90),
.A2(n_5),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_93),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_91),
.Y(n_95)
);


endmodule