module real_jpeg_33732_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_0),
.Y(n_173)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_0),
.Y(n_478)
);

AO22x1_ASAP7_75t_L g58 ( 
.A1(n_1),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_1),
.A2(n_63),
.B1(n_215),
.B2(n_218),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_1),
.A2(n_63),
.B1(n_518),
.B2(n_519),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_2),
.A2(n_73),
.B1(n_74),
.B2(n_78),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_2),
.A2(n_73),
.B1(n_225),
.B2(n_229),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_3),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_4),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_4),
.Y(n_118)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_5),
.Y(n_82)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_5),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_6),
.A2(n_182),
.B1(n_183),
.B2(n_186),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_6),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_6),
.A2(n_186),
.B1(n_276),
.B2(n_336),
.Y(n_511)
);

AO22x1_ASAP7_75t_L g175 ( 
.A1(n_7),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_8),
.Y(n_112)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_8),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_8),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_9),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_9),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_9),
.A2(n_123),
.B1(n_133),
.B2(n_136),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_9),
.A2(n_123),
.B1(n_275),
.B2(n_280),
.Y(n_274)
);

OAI22x1_ASAP7_75t_L g365 ( 
.A1(n_9),
.A2(n_123),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_10),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_11),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_11),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_11),
.A2(n_160),
.B1(n_299),
.B2(n_303),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_11),
.A2(n_160),
.B1(n_381),
.B2(n_385),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_11),
.A2(n_160),
.B1(n_471),
.B2(n_473),
.Y(n_470)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_12),
.Y(n_197)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_12),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_13),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_13),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_13),
.B(n_165),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_13),
.A2(n_295),
.B1(n_390),
.B2(n_392),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_13),
.B(n_306),
.Y(n_408)
);

OAI21xp33_ASAP7_75t_L g484 ( 
.A1(n_13),
.A2(n_180),
.B(n_419),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_14),
.A2(n_239),
.B1(n_243),
.B2(n_244),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_14),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_14),
.A2(n_243),
.B1(n_252),
.B2(n_254),
.Y(n_251)
);

AO22x1_ASAP7_75t_L g319 ( 
.A1(n_14),
.A2(n_64),
.B1(n_243),
.B2(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_15),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_16),
.A2(n_86),
.B1(n_92),
.B2(n_93),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_16),
.A2(n_92),
.B1(n_259),
.B2(n_263),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_16),
.A2(n_92),
.B1(n_336),
.B2(n_339),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_16),
.A2(n_92),
.B1(n_411),
.B2(n_414),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_499),
.Y(n_17)
);

OAI21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_325),
.B(n_495),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_265),
.B(n_307),
.Y(n_20)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_21),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_166),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_22),
.B(n_167),
.C(n_231),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.C(n_129),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_23),
.B(n_268),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_51),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_24),
.B(n_51),
.Y(n_311)
);

AOI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.A3(n_35),
.B1(n_40),
.B2(n_43),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_30),
.Y(n_302)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_34),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_34),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_34),
.Y(n_157)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_38),
.Y(n_147)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_39),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_39),
.Y(n_164)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_39),
.Y(n_262)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_40),
.Y(n_296)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_45),
.A2(n_100),
.B1(n_102),
.B2(n_106),
.Y(n_99)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_46),
.Y(n_358)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_47),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_58),
.B1(n_68),
.B2(n_72),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_52),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_52),
.A2(n_58),
.B1(n_68),
.B2(n_319),
.Y(n_318)
);

NAND2x1_ASAP7_75t_SL g364 ( 
.A(n_52),
.B(n_365),
.Y(n_364)
);

OA21x2_ASAP7_75t_L g507 ( 
.A1(n_52),
.A2(n_175),
.B(n_508),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_55),
.Y(n_185)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_55),
.Y(n_193)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_55),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_55),
.Y(n_431)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_57),
.Y(n_488)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_61),
.Y(n_182)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_66),
.Y(n_178)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_66),
.Y(n_367)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_67),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_71),
.Y(n_236)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_72),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_80),
.Y(n_413)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_82),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_82),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_82),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_83),
.A2(n_84),
.B1(n_129),
.B2(n_130),
.Y(n_268)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_97),
.B(n_119),
.Y(n_84)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_85),
.Y(n_305)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_95),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_96),
.Y(n_522)
);

OAI22x1_ASAP7_75t_L g248 ( 
.A1(n_97),
.A2(n_249),
.B1(n_250),
.B2(n_256),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_97),
.A2(n_119),
.B(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_98),
.A2(n_298),
.B1(n_305),
.B2(n_306),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_SL g316 ( 
.A(n_98),
.B(n_121),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_98),
.A2(n_120),
.B1(n_251),
.B2(n_517),
.Y(n_516)
);

AND2x4_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_109),
.Y(n_98)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_103),
.Y(n_360)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_112),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_112),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_114),
.Y(n_339)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_120),
.Y(n_256)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_121),
.Y(n_249)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_128),
.Y(n_349)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_158),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_138),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_132),
.B(n_165),
.Y(n_289)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_137),
.Y(n_294)
);

AO22x1_ASAP7_75t_L g257 ( 
.A1(n_138),
.A2(n_159),
.B1(n_165),
.B2(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_138),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_138),
.B(n_258),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_151),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_142),
.B1(n_146),
.B2(n_148),
.Y(n_139)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.Y(n_151)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_153),
.Y(n_255)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_154),
.Y(n_393)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx4f_ASAP7_75t_SL g264 ( 
.A(n_164),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_231),
.Y(n_166)
);

XOR2x2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_187),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_168),
.B(n_188),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_174),
.B1(n_180),
.B2(n_181),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_172),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_180),
.A2(n_181),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_180),
.A2(n_410),
.B(n_419),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_180),
.A2(n_410),
.B1(n_470),
.B2(n_487),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_214),
.B1(n_223),
.B2(n_224),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_214),
.B1(n_223),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_189),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_189),
.A2(n_223),
.B1(n_335),
.B2(n_380),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_L g404 ( 
.A1(n_189),
.A2(n_380),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_189),
.A2(n_223),
.B1(n_224),
.B2(n_511),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_202),
.Y(n_189)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_190),
.Y(n_287)
);

OAI22x1_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_194),
.B1(n_198),
.B2(n_200),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_197),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_207),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_207),
.Y(n_285)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_217),
.Y(n_346)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_222),
.Y(n_453)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_228),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_247),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_232),
.B(n_248),
.C(n_257),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_237),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_235),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_236),
.Y(n_420)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_238),
.Y(n_286)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_246),
.Y(n_461)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_257),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_SL g306 ( 
.A(n_256),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_256),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_266),
.B(n_497),
.C(n_498),
.Y(n_496)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.C(n_270),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_267),
.B(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_269),
.B(n_271),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_288),
.C(n_297),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_297),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_286),
.B2(n_287),
.Y(n_272)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_273),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_274),
.B(n_287),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_274),
.Y(n_405)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_279),
.Y(n_354)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_279),
.Y(n_443)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_285),
.Y(n_386)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_287),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_310),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_289),
.B(n_524),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_295),
.B(n_296),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_295),
.B(n_348),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_295),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_295),
.B(n_441),
.Y(n_440)
);

OA21x2_ASAP7_75t_R g459 ( 
.A1(n_295),
.A2(n_440),
.B(n_460),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_295),
.B(n_406),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_295),
.B(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_301),
.Y(n_518)
);

INVx3_ASAP7_75t_SL g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_302),
.Y(n_391)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_323),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_308),
.B(n_323),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.C(n_312),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_309),
.B(n_374),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_311),
.B(n_312),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_317),
.C(n_318),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_314),
.B(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_318),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_319),
.B(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_320),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_320),
.B(n_482),
.Y(n_481)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_375),
.B(n_493),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_373),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_329),
.B(n_494),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_333),
.C(n_342),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_331),
.B(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_333),
.A2(n_334),
.B1(n_342),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_340),
.B(n_341),
.Y(n_334)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

OA21x2_ASAP7_75t_SL g458 ( 
.A1(n_340),
.A2(n_341),
.B(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_342),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_361),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_343),
.B(n_361),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_347),
.B1(n_350),
.B2(n_355),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_359),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2x1_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_364),
.A2(n_470),
.B(n_474),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_SL g419 ( 
.A(n_365),
.B(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_372),
.Y(n_418)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_373),
.Y(n_494)
);

AOI21x1_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_425),
.B(n_492),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_400),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_397),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_378),
.B(n_397),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_387),
.C(n_394),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_379),
.B(n_388),
.Y(n_423)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_395),
.A2(n_396),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_424),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_421),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_421),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_407),
.C(n_409),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_404),
.B(n_408),
.Y(n_464)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_409),
.Y(n_463)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_420),
.Y(n_483)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_424),
.B(n_491),
.Y(n_490)
);

AO21x1_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_465),
.B(n_490),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_462),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_427),
.B(n_462),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_458),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_428),
.B(n_458),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_429),
.A2(n_439),
.B1(n_444),
.B2(n_449),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_432),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx6_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_454),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_486),
.C(n_489),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_480),
.B(n_485),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_479),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_479),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_484),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_525),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_502),
.B(n_503),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_505),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_513),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_507),
.A2(n_509),
.B1(n_510),
.B2(n_512),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_507),
.Y(n_512)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_523),
.Y(n_515)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);


endmodule