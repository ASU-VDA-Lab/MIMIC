module fake_jpeg_21342_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

INVx8_ASAP7_75t_SL g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_17),
.B(n_20),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_51),
.B1(n_53),
.B2(n_58),
.Y(n_70)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_64),
.Y(n_76)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_67),
.Y(n_77)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_0),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_58),
.B1(n_48),
.B2(n_59),
.Y(n_72)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_57),
.B1(n_54),
.B2(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_46),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_48),
.B(n_55),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_2),
.C(n_3),
.Y(n_91)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_90),
.Y(n_103)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_42),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_70),
.C(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_3),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_92),
.B(n_4),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_97),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_27),
.B(n_39),
.C(n_38),
.D(n_8),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_4),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_104),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_25),
.C(n_37),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_29),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_85),
.B(n_12),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_5),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_109),
.B(n_112),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_83),
.B(n_6),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_6),
.B(n_9),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_93),
.C(n_95),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_114),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_103),
.B1(n_99),
.B2(n_98),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_115),
.A2(n_116),
.B1(n_112),
.B2(n_82),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_107),
.B1(n_96),
.B2(n_113),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_117),
.B(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_10),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_11),
.B(n_28),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_31),
.B(n_34),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_36),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_40),
.Y(n_125)
);


endmodule