module fake_jpeg_25545_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_9),
.B(n_6),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_25),
.B1(n_20),
.B2(n_4),
.Y(n_33)
);

CKINVDCx12_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_3),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_5),
.B(n_8),
.Y(n_38)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_15),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_30),
.B(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_20),
.B1(n_11),
.B2(n_10),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_33),
.B1(n_39),
.B2(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_25),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_19),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_22),
.A2(n_16),
.B1(n_12),
.B2(n_15),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_42),
.B1(n_44),
.B2(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_22),
.B1(n_21),
.B2(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_28),
.B1(n_23),
.B2(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_46),
.B(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_34),
.B1(n_15),
.B2(n_16),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_47),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_53),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_34),
.C(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_42),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_52),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_44),
.B(n_15),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_64),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_14),
.B1(n_19),
.B2(n_58),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_66),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_66),
.B(n_14),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_71),
.A2(n_70),
.B(n_68),
.Y(n_72)
);


endmodule