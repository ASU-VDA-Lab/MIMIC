module fake_jpeg_20204_n_75 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_75);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_75;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_71;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_72;
wire n_49;
wire n_24;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_74;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_25;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_6),
.A2(n_9),
.B(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_14),
.B(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_46),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_27),
.B1(n_33),
.B2(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_27),
.A2(n_34),
.B1(n_24),
.B2(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_41),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_57),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_55),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_59),
.C(n_57),
.Y(n_62)
);

MAJx2_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_60),
.C(n_63),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_59),
.B(n_53),
.Y(n_65)
);

OA21x2_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_66),
.B(n_51),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_53),
.B(n_30),
.Y(n_66)
);

MAJx2_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_68),
.C(n_56),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_37),
.C(n_36),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_25),
.B(n_42),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_70),
.B(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_73),
.A2(n_72),
.B(n_52),
.C(n_49),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_54),
.Y(n_75)
);


endmodule