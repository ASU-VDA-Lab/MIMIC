module fake_jpeg_21763_n_249 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx8_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_35),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_6),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVxp67_ASAP7_75t_SL g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_14),
.B1(n_18),
.B2(n_19),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_17),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_14),
.B1(n_18),
.B2(n_27),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_37),
.B(n_32),
.C(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_54),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_14),
.B1(n_18),
.B2(n_27),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_16),
.B1(n_15),
.B2(n_20),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_31),
.A2(n_16),
.B1(n_15),
.B2(n_20),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_34),
.B(n_26),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_64),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_37),
.B1(n_32),
.B2(n_29),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_73),
.B1(n_44),
.B2(n_43),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_74),
.B1(n_44),
.B2(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_70),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_30),
.B1(n_34),
.B2(n_6),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_50),
.B1(n_51),
.B2(n_41),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_48),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_72),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_53),
.B1(n_37),
.B2(n_32),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_34),
.B1(n_30),
.B2(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_75),
.B(n_86),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_65),
.B1(n_74),
.B2(n_85),
.Y(n_96)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_90),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_72),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_94),
.B1(n_70),
.B2(n_60),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_43),
.A3(n_51),
.B1(n_17),
.B2(n_24),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_71),
.C(n_64),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_89),
.B1(n_68),
.B2(n_62),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_51),
.B1(n_41),
.B2(n_2),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_63),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_97),
.B1(n_112),
.B2(n_24),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_102),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_67),
.B(n_71),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_103),
.B(n_109),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_93),
.B1(n_77),
.B2(n_83),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_107),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_61),
.C(n_58),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_91),
.C(n_26),
.Y(n_134)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_108),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_75),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_79),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_62),
.B1(n_61),
.B2(n_39),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_128),
.B1(n_105),
.B2(n_102),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_78),
.B(n_89),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_119),
.A2(n_124),
.B(n_135),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_123),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_87),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_125),
.C(n_134),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_76),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_84),
.B(n_91),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_129),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_79),
.B1(n_39),
.B2(n_59),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_39),
.Y(n_132)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

OAI22x1_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_97),
.B1(n_112),
.B2(n_96),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_138),
.B(n_143),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_114),
.B(n_109),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_147),
.B(n_151),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_101),
.B(n_114),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_109),
.C(n_96),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_145),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_96),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_101),
.C(n_108),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_134),
.C(n_124),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_0),
.B(n_1),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_120),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_150),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_26),
.B(n_28),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_154),
.Y(n_157)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_59),
.B1(n_25),
.B2(n_23),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_155),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_161),
.B(n_162),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

NAND2xp33_ASAP7_75t_SL g164 ( 
.A(n_136),
.B(n_126),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_166),
.B1(n_139),
.B2(n_142),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_168),
.B(n_169),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_171),
.C(n_175),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_122),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_145),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_125),
.C(n_123),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_135),
.B1(n_121),
.B2(n_127),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_120),
.C(n_116),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_186),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_171),
.C(n_167),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_160),
.C(n_162),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_184),
.B(n_187),
.Y(n_197)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_140),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_191),
.B(n_176),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_144),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_176),
.Y(n_201)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_139),
.Y(n_192)
);

BUFx24_ASAP7_75t_SL g199 ( 
.A(n_192),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_205),
.C(n_147),
.Y(n_211)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_204),
.Y(n_209)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_202),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_182),
.A2(n_169),
.B1(n_165),
.B2(n_158),
.Y(n_198)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_156),
.Y(n_217)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_180),
.A2(n_158),
.B1(n_166),
.B2(n_163),
.Y(n_203)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_116),
.C(n_115),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_141),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_193),
.A2(n_178),
.B1(n_189),
.B2(n_186),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_207),
.A2(n_208),
.B(n_214),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_178),
.B1(n_141),
.B2(n_177),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_218),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_0),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_SL g214 ( 
.A1(n_199),
.A2(n_156),
.A3(n_155),
.B1(n_12),
.B2(n_13),
.C1(n_10),
.C2(n_7),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_156),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_216),
.B(n_200),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_201),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_59),
.C(n_25),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_197),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_219),
.B(n_224),
.CI(n_218),
.CON(n_229),
.SN(n_229)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_220),
.A2(n_222),
.B1(n_226),
.B2(n_1),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_21),
.B1(n_28),
.B2(n_4),
.Y(n_234)
);

OAI21x1_ASAP7_75t_SL g222 ( 
.A1(n_217),
.A2(n_200),
.B(n_9),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_8),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_7),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_227),
.B(n_228),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_229),
.B(n_234),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_213),
.A3(n_208),
.B1(n_207),
.B2(n_21),
.C1(n_10),
.C2(n_7),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_231),
.B(n_1),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_12),
.B(n_9),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_21),
.C(n_2),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_233),
.A2(n_224),
.B(n_3),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_SL g240 ( 
.A1(n_235),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_219),
.B(n_28),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_236),
.B(n_229),
.Y(n_239)
);

OAI21x1_ASAP7_75t_SL g243 ( 
.A1(n_238),
.A2(n_240),
.B(n_3),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_241),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_233),
.B(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_232),
.C(n_240),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_3),
.Y(n_246)
);

OAI321xp33_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_246),
.A3(n_244),
.B1(n_5),
.B2(n_4),
.C(n_28),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_5),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_5),
.Y(n_249)
);


endmodule