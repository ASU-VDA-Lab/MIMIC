module fake_jpeg_29081_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_8),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_56),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_58),
.Y(n_61)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_1),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_19),
.B1(n_32),
.B2(n_31),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_42),
.B1(n_48),
.B2(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_2),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_66),
.Y(n_73)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_46),
.Y(n_75)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_69),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_39),
.B1(n_50),
.B2(n_41),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_82),
.B1(n_4),
.B2(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_84),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_80),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_39),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_79),
.C(n_85),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_36),
.C(n_45),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_65),
.C(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_3),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_97),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_62),
.B(n_45),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_96),
.B(n_99),
.C(n_101),
.Y(n_106)
);

XOR2x2_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_21),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_62),
.C(n_9),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_20),
.B(n_34),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_18),
.B(n_28),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_6),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_8),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_22),
.B(n_27),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_108),
.B1(n_11),
.B2(n_87),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_24),
.C(n_14),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_16),
.C(n_17),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_112),
.A2(n_92),
.B1(n_100),
.B2(n_107),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_103),
.C(n_94),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_115),
.A2(n_116),
.B(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_117),
.B(n_113),
.Y(n_118)
);

NOR4xp25_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_106),
.C(n_114),
.D(n_102),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_114),
.C(n_106),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_95),
.Y(n_121)
);


endmodule