module fake_jpeg_24020_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_1),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_24),
.B1(n_27),
.B2(n_19),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_68),
.B1(n_19),
.B2(n_33),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_28),
.B1(n_34),
.B2(n_23),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_55),
.B1(n_28),
.B2(n_20),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_19),
.B1(n_17),
.B2(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_57),
.Y(n_104)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_18),
.B(n_22),
.C(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_64),
.B(n_18),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_25),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_40),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_35),
.B1(n_17),
.B2(n_33),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_74),
.Y(n_120)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_87),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_81),
.Y(n_121)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_84),
.Y(n_135)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_85),
.A2(n_90),
.B1(n_91),
.B2(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_98),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_89),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_47),
.B1(n_46),
.B2(n_37),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_29),
.B1(n_25),
.B2(n_23),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_106),
.B1(n_29),
.B2(n_22),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_20),
.B1(n_31),
.B2(n_35),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_100),
.B1(n_31),
.B2(n_65),
.Y(n_123)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_47),
.B1(n_41),
.B2(n_43),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_99),
.B1(n_105),
.B2(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_51),
.Y(n_98)
);

AOI222xp33_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_41),
.B1(n_44),
.B2(n_43),
.C1(n_34),
.C2(n_23),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_38),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_107),
.Y(n_131)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_56),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_29),
.B1(n_34),
.B2(n_25),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_38),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_66),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_39),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_50),
.A2(n_20),
.B1(n_35),
.B2(n_31),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_49),
.B(n_38),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_32),
.Y(n_132)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_116),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_87),
.C(n_98),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_104),
.C(n_109),
.Y(n_162)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_125),
.B(n_105),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_126),
.B1(n_100),
.B2(n_110),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_61),
.B1(n_57),
.B2(n_70),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_81),
.A2(n_39),
.B1(n_32),
.B2(n_30),
.Y(n_126)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_91),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_18),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_138),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_84),
.Y(n_138)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_145),
.B(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_140),
.B(n_78),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_149),
.B(n_151),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_78),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_72),
.B(n_86),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_152),
.A2(n_3),
.B(n_4),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_164),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_157),
.B1(n_172),
.B2(n_147),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_72),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_158),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_85),
.B1(n_99),
.B2(n_107),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_101),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_141),
.A2(n_112),
.B1(n_82),
.B2(n_79),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_163),
.B1(n_136),
.B2(n_133),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_161),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_165),
.C(n_169),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_74),
.B(n_73),
.C(n_39),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_120),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_115),
.C(n_118),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_83),
.C(n_80),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_174),
.B(n_3),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_167),
.B(n_170),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_76),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_171),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_115),
.B(n_134),
.C(n_132),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_135),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_136),
.C(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_137),
.B1(n_108),
.B2(n_113),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_116),
.Y(n_173)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_128),
.B(n_18),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_32),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_1),
.Y(n_203)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_177),
.B(n_183),
.Y(n_222)
);

AO21x2_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_137),
.B(n_103),
.Y(n_178)
);

AOI22x1_ASAP7_75t_L g229 ( 
.A1(n_178),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_179),
.A2(n_184),
.B1(n_187),
.B2(n_194),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_180),
.A2(n_191),
.B1(n_202),
.B2(n_159),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_142),
.B1(n_143),
.B2(n_130),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_142),
.A3(n_127),
.B1(n_30),
.B2(n_16),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_188),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_174),
.A2(n_127),
.B1(n_119),
.B2(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_15),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_208),
.B(n_173),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_119),
.B1(n_117),
.B2(n_93),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_154),
.A2(n_30),
.B1(n_16),
.B2(n_139),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_205),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_146),
.A2(n_30),
.B1(n_16),
.B2(n_139),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_197),
.A2(n_167),
.B1(n_170),
.B2(n_150),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_15),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_148),
.B(n_2),
.Y(n_204)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_2),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_13),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_207),
.A2(n_155),
.B(n_145),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_181),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_218),
.C(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_233),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_219),
.B1(n_223),
.B2(n_187),
.Y(n_240)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_165),
.C(n_162),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_226),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_215),
.B(n_228),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_199),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_176),
.A2(n_161),
.B(n_146),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_217),
.A2(n_220),
.B(n_225),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_169),
.C(n_171),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_178),
.A2(n_164),
.B1(n_175),
.B2(n_150),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_176),
.A2(n_3),
.B(n_4),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_159),
.C(n_5),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g225 ( 
.A(n_178),
.B(n_193),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_4),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_208),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_196),
.B(n_13),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_236),
.B1(n_202),
.B2(n_205),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_178),
.Y(n_231)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_231),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_182),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_232),
.Y(n_249)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_190),
.A2(n_13),
.B(n_6),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_240),
.A2(n_259),
.B(n_255),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_231),
.A2(n_192),
.B1(n_188),
.B2(n_190),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_243),
.A2(n_253),
.B1(n_256),
.B2(n_224),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_257),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_247),
.A2(n_259),
.B1(n_241),
.B2(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_213),
.B(n_200),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_193),
.Y(n_252)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_235),
.B1(n_219),
.B2(n_211),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_211),
.A2(n_197),
.B1(n_194),
.B2(n_177),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_203),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_258),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_204),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_224),
.A2(n_180),
.B1(n_191),
.B2(n_185),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_198),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_214),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_262),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_239),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_266),
.B(n_13),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_272),
.C(n_273),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_275),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_238),
.A2(n_225),
.B1(n_230),
.B2(n_229),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_270),
.B1(n_5),
.B2(n_7),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_225),
.B1(n_229),
.B2(n_222),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_234),
.C(n_221),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_215),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_212),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_277),
.B1(n_280),
.B2(n_256),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_243),
.B(n_234),
.C(n_209),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_279),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_233),
.C(n_220),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_255),
.A2(n_236),
.B(n_6),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_282),
.Y(n_304)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_258),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_279),
.B(n_272),
.Y(n_306)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_291),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_264),
.A2(n_249),
.B1(n_254),
.B2(n_252),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_245),
.B1(n_244),
.B2(n_227),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_226),
.B1(n_7),
.B2(n_8),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_294),
.A2(n_295),
.B1(n_280),
.B2(n_271),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_5),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_9),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_274),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_303),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_265),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_306),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_293),
.Y(n_302)
);

OAI22x1_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_284),
.B1(n_292),
.B2(n_281),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_265),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_285),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_282),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_310),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_290),
.C(n_296),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_311),
.A2(n_315),
.B(n_318),
.Y(n_327)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_274),
.B1(n_295),
.B2(n_266),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_297),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_304),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_283),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_320),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_268),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_303),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_322),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_299),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_325),
.B(n_273),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_288),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_311),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_329),
.B(n_330),
.Y(n_332)
);

NAND4xp25_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_314),
.C(n_317),
.D(n_267),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_324),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_328),
.B(n_323),
.Y(n_334)
);

AOI321xp33_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_332),
.A3(n_333),
.B1(n_321),
.B2(n_12),
.C(n_11),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_9),
.B(n_10),
.Y(n_336)
);

NOR3xp33_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_9),
.C(n_10),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_10),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_11),
.B1(n_12),
.B2(n_293),
.Y(n_339)
);


endmodule