module fake_jpeg_14718_n_183 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_38),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_20),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_30),
.B1(n_15),
.B2(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_18),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_15),
.A2(n_2),
.B(n_4),
.Y(n_44)
);

AND2x4_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_5),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_56),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_20),
.B1(n_19),
.B2(n_18),
.Y(n_78)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_50),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_19),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_57),
.B(n_44),
.Y(n_70)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_58),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_68),
.Y(n_94)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_73),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_32),
.B(n_31),
.C(n_21),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_39),
.B(n_22),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_24),
.B(n_32),
.Y(n_102)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_80),
.B1(n_21),
.B2(n_6),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_16),
.B1(n_60),
.B2(n_36),
.Y(n_80)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_40),
.B1(n_34),
.B2(n_38),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_40),
.B1(n_62),
.B2(n_38),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_22),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_42),
.Y(n_106)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_83),
.B(n_38),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_85),
.Y(n_105)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_16),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_90),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_28),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_55),
.B1(n_53),
.B2(n_34),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_95),
.B(n_84),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_25),
.B1(n_31),
.B2(n_24),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_102),
.B(n_88),
.Y(n_113)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_66),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_103),
.B1(n_104),
.B2(n_110),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_76),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_81),
.C(n_72),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_106),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_40),
.B1(n_62),
.B2(n_38),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_42),
.B1(n_7),
.B2(n_8),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_112),
.B(n_116),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_122),
.B(n_91),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_114),
.B(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_82),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_5),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_127),
.C(n_128),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_83),
.C(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_125),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_67),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_79),
.C(n_73),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_139),
.B1(n_117),
.B2(n_110),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_121),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_133),
.B(n_135),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_100),
.B(n_95),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_124),
.C(n_118),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_146),
.C(n_152),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_128),
.C(n_127),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_117),
.B1(n_104),
.B2(n_111),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_154),
.B1(n_141),
.B2(n_79),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_129),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_113),
.C(n_98),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_130),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_92),
.B1(n_103),
.B2(n_97),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_143),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_161),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_148),
.B(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_134),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_142),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_163),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_152),
.C(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_158),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_101),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_173),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_168),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_156),
.B(n_144),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_136),
.C(n_11),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_136),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_66),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_166),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_10),
.B(n_11),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_177),
.C(n_176),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_74),
.A3(n_85),
.B1(n_13),
.B2(n_14),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_10),
.Y(n_183)
);


endmodule