module fake_jpeg_2064_n_315 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_4),
.B(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_46),
.Y(n_137)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_57),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_4),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_68),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

NOR3xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_86),
.C(n_30),
.Y(n_108)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx2_ASAP7_75t_SL g113 ( 
.A(n_67),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_21),
.B(n_4),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_21),
.B(n_5),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_79),
.Y(n_114)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_6),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_80),
.Y(n_116)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_6),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_45),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_40),
.Y(n_123)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_6),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_87),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_28),
.C(n_42),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_89),
.B(n_93),
.C(n_127),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_28),
.B1(n_25),
.B2(n_42),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_92),
.A2(n_106),
.B1(n_110),
.B2(n_117),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_25),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_49),
.A2(n_23),
.B1(n_44),
.B2(n_33),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_56),
.A2(n_30),
.B1(n_43),
.B2(n_41),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_62),
.A2(n_23),
.B1(n_44),
.B2(n_33),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_54),
.A2(n_43),
.B1(n_41),
.B2(n_40),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_88),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_125),
.B(n_131),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_50),
.A2(n_63),
.B1(n_60),
.B2(n_35),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_128),
.A2(n_130),
.B1(n_138),
.B2(n_137),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_61),
.A2(n_35),
.B1(n_34),
.B2(n_11),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_46),
.B(n_34),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_70),
.A2(n_7),
.B1(n_10),
.B2(n_12),
.Y(n_134)
);

AOI222xp33_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_108),
.C2(n_138),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_46),
.B(n_7),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_69),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_79),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_139),
.B(n_140),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_69),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_75),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_142),
.B(n_159),
.Y(n_198)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_144),
.Y(n_210)
);

OR2x2_ASAP7_75t_SL g145 ( 
.A(n_133),
.B(n_67),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_127),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_158),
.Y(n_190)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_133),
.A2(n_79),
.B1(n_75),
.B2(n_67),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_149),
.B1(n_162),
.B2(n_176),
.Y(n_187)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_121),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_156),
.Y(n_189)
);

INVx2_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_15),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_161),
.Y(n_204)
);

INVx3_ASAP7_75t_SL g161 ( 
.A(n_100),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_117),
.A2(n_106),
.B1(n_110),
.B2(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_166),
.Y(n_211)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_170),
.Y(n_182)
);

OR2x4_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_116),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_168),
.A2(n_145),
.B(n_163),
.C(n_149),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g169 ( 
.A1(n_128),
.A2(n_124),
.B1(n_112),
.B2(n_132),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_143),
.B1(n_161),
.B2(n_155),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_107),
.B(n_94),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_172),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_103),
.Y(n_172)
);

AO22x1_ASAP7_75t_SL g173 ( 
.A1(n_112),
.A2(n_132),
.B1(n_96),
.B2(n_111),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_177),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_151),
.Y(n_207)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_100),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_180),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_124),
.A2(n_111),
.B1(n_102),
.B2(n_95),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_179),
.A2(n_154),
.B1(n_177),
.B2(n_146),
.Y(n_203)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_95),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_129),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_207),
.C(n_196),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_162),
.B(n_164),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_186),
.A2(n_188),
.B(n_209),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_102),
.B(n_122),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_141),
.A2(n_113),
.B1(n_168),
.B2(n_173),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_199),
.B1(n_188),
.B2(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_194),
.B(n_182),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_203),
.B1(n_206),
.B2(n_189),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_169),
.B1(n_153),
.B2(n_144),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_148),
.B(n_152),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_209),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_157),
.B1(n_156),
.B2(n_151),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_168),
.CI(n_145),
.CON(n_209),
.SN(n_209)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_213),
.A2(n_222),
.B1(n_223),
.B2(n_234),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_187),
.A2(n_201),
.B1(n_191),
.B2(n_181),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_197),
.B(n_202),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_181),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_218),
.B(n_221),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_193),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_216),
.B(n_231),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_194),
.B(n_185),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_208),
.Y(n_244)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

AO221x1_ASAP7_75t_L g254 ( 
.A1(n_219),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.C(n_233),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_182),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_225),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_184),
.B1(n_195),
.B2(n_196),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_223),
.A2(n_208),
.B1(n_205),
.B2(n_212),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_226),
.B1(n_233),
.B2(n_227),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_184),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_200),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_202),
.C(n_190),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_234),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_190),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_190),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_210),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_235),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_183),
.B(n_210),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_236),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_203),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_238),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_239),
.A2(n_249),
.B(n_238),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_251),
.B1(n_227),
.B2(n_228),
.Y(n_265)
);

OA21x2_ASAP7_75t_SL g269 ( 
.A1(n_244),
.A2(n_228),
.B(n_254),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_217),
.Y(n_245)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_248),
.Y(n_258)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_222),
.Y(n_250)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_213),
.A2(n_224),
.B1(n_231),
.B2(n_215),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_252),
.A2(n_245),
.B1(n_244),
.B2(n_247),
.Y(n_271)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_229),
.B(n_215),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_256),
.A2(n_263),
.B(n_270),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_225),
.C(n_220),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_262),
.C(n_266),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_232),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_261),
.B(n_242),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_229),
.C(n_227),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_238),
.A2(n_252),
.B(n_240),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_243),
.B1(n_255),
.B2(n_250),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_219),
.C(n_228),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_241),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_243),
.B1(n_246),
.B2(n_248),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_270),
.A2(n_245),
.B(n_254),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_266),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_279),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_258),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_257),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_257),
.B1(n_264),
.B2(n_259),
.Y(n_290)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_290),
.B1(n_273),
.B2(n_263),
.Y(n_294)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_260),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_286),
.B(n_271),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_262),
.C(n_256),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_276),
.C(n_279),
.Y(n_299)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_296),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_277),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_276),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_298),
.C(n_299),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_269),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_288),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_264),
.A3(n_288),
.B1(n_291),
.B2(n_289),
.C1(n_280),
.C2(n_274),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_302),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_305),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_299),
.B(n_295),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_297),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_307),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_296),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_300),
.B(n_290),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_310),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_311),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_308),
.B1(n_267),
.B2(n_259),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_314),
.A2(n_313),
.B(n_272),
.Y(n_315)
);


endmodule