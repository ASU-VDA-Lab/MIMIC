module fake_jpeg_571_n_130 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_14),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_51),
.Y(n_55)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_46),
.B1(n_39),
.B2(n_40),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_53),
.B(n_33),
.C(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_59),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_74),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_51),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_73),
.Y(n_80)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_70),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_44),
.C(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_64),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_54),
.B(n_66),
.C(n_69),
.Y(n_79)
);

MAJx3_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_35),
.C(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_39),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_62),
.B(n_54),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_78),
.B(n_79),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_72),
.B(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_12),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_1),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_58),
.B1(n_20),
.B2(n_21),
.Y(n_101)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_93),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_57),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

HAxp5_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_38),
.CON(n_92),
.SN(n_92)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_6),
.B(n_8),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_1),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_18),
.Y(n_96)
);

FAx1_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_102),
.CI(n_8),
.CON(n_115),
.SN(n_115)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_99),
.B(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_31),
.B1(n_22),
.B2(n_23),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_13),
.C(n_30),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_15),
.Y(n_114)
);

AOI221xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_107),
.B1(n_111),
.B2(n_114),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_113),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_115),
.A2(n_92),
.B1(n_102),
.B2(n_9),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_91),
.C(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_116),
.B(n_119),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_109),
.A2(n_101),
.B1(n_11),
.B2(n_24),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_120),
.A2(n_105),
.B1(n_110),
.B2(n_104),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_121),
.A2(n_122),
.B1(n_118),
.B2(n_113),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

NOR2xp67_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_116),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_125),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_106),
.B(n_120),
.C(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_10),
.Y(n_130)
);


endmodule