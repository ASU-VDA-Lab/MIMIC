module real_aes_3205_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_1103, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_1103;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_1064;
wire n_540;
wire n_1075;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_923;
wire n_1034;
wire n_894;
wire n_952;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_932;
wire n_399;
wire n_1021;
wire n_700;
wire n_948;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_1078;
wire n_495;
wire n_1072;
wire n_892;
wire n_370;
wire n_994;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_1053;
wire n_976;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_1081;
wire n_1084;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_1100;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1014;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_1083;
wire n_727;
wire n_397;
wire n_749;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_314;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_1090;
wire n_456;
wire n_359;
wire n_717;
wire n_982;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_371;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_1045;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_601;
wire n_500;
wire n_1101;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
wire n_429;
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_0), .A2(n_295), .B1(n_583), .B2(n_584), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_1), .A2(n_129), .B1(n_448), .B2(n_454), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_2), .A2(n_198), .B1(n_456), .B2(n_457), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_3), .B(n_375), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_4), .A2(n_237), .B1(n_424), .B2(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_5), .A2(n_280), .B1(n_496), .B2(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g738 ( .A(n_6), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_7), .A2(n_245), .B1(n_692), .B2(n_693), .C(n_694), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_8), .A2(n_255), .B1(n_356), .B2(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g922 ( .A(n_9), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g1089 ( .A1(n_10), .A2(n_84), .B1(n_740), .B2(n_1090), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_11), .A2(n_175), .B1(n_456), .B2(n_457), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g1063 ( .A1(n_12), .A2(n_190), .B1(n_451), .B2(n_1064), .Y(n_1063) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_13), .B(n_332), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_14), .A2(n_257), .B1(n_482), .B2(n_483), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_15), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_16), .A2(n_234), .B1(n_492), .B2(n_678), .Y(n_696) );
AOI21xp33_ASAP7_75t_L g1073 ( .A1(n_17), .A2(n_558), .B(n_1074), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_18), .A2(n_91), .B1(n_488), .B2(n_542), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_19), .A2(n_34), .B1(n_482), .B2(n_483), .Y(n_724) );
INVx1_ASAP7_75t_L g367 ( .A(n_20), .Y(n_367) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_21), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_22), .A2(n_88), .B1(n_854), .B2(n_856), .Y(n_853) );
INVx1_ASAP7_75t_L g578 ( .A(n_23), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g1096 ( .A1(n_24), .A2(n_289), .B1(n_413), .B2(n_584), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_25), .A2(n_36), .B1(n_453), .B2(n_454), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_26), .A2(n_117), .B1(n_495), .B2(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g668 ( .A(n_27), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_28), .A2(n_127), .B1(n_488), .B2(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g1075 ( .A(n_29), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_30), .A2(n_195), .B1(n_465), .B2(n_470), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_31), .B(n_460), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_32), .A2(n_147), .B1(n_403), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_33), .A2(n_160), .B1(n_542), .B2(n_588), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g561 ( .A1(n_35), .A2(n_291), .B1(n_462), .B2(n_463), .C(n_562), .Y(n_561) );
AO22x1_ASAP7_75t_L g323 ( .A1(n_37), .A2(n_54), .B1(n_324), .B2(n_348), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_38), .A2(n_784), .B(n_786), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_39), .A2(n_169), .B1(n_349), .B2(n_678), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_40), .A2(n_204), .B1(n_839), .B2(n_843), .Y(n_924) );
INVx1_ASAP7_75t_L g801 ( .A(n_41), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_42), .A2(n_98), .B1(n_418), .B2(n_482), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_43), .A2(n_51), .B1(n_628), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_44), .A2(n_93), .B1(n_469), .B2(n_470), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_45), .A2(n_148), .B1(n_425), .B2(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_46), .A2(n_297), .B1(n_450), .B2(n_451), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_47), .A2(n_122), .B1(n_413), .B2(n_483), .Y(n_703) );
INVx1_ASAP7_75t_L g882 ( .A(n_48), .Y(n_882) );
AO22x1_ASAP7_75t_L g562 ( .A1(n_49), .A2(n_69), .B1(n_470), .B2(n_537), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_50), .A2(n_214), .B1(n_572), .B2(n_573), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_52), .A2(n_251), .B1(n_462), .B2(n_470), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_53), .B(n_389), .Y(n_620) );
OA22x2_ASAP7_75t_L g347 ( .A1(n_55), .A2(n_137), .B1(n_332), .B2(n_346), .Y(n_347) );
INVx1_ASAP7_75t_L g362 ( .A(n_55), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g1067 ( .A1(n_56), .A2(n_97), .B1(n_434), .B2(n_765), .Y(n_1067) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_57), .A2(n_66), .B1(n_369), .B2(n_375), .C(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_58), .A2(n_258), .B1(n_542), .B2(n_588), .Y(n_1098) );
AOI221x1_ASAP7_75t_L g751 ( .A1(n_59), .A2(n_224), .B1(n_531), .B2(n_543), .C(n_752), .Y(n_751) );
INVxp67_ASAP7_75t_L g721 ( .A(n_60), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_61), .A2(n_128), .B1(n_488), .B2(n_489), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_62), .A2(n_307), .B1(n_403), .B2(n_413), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g1070 ( .A1(n_63), .A2(n_115), .B1(n_356), .B2(n_755), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_64), .A2(n_281), .B1(n_462), .B2(n_470), .Y(n_797) );
INVx1_ASAP7_75t_L g345 ( .A(n_65), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g363 ( .A1(n_65), .A2(n_137), .B(n_364), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_65), .B(n_156), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_67), .A2(n_264), .B1(n_433), .B2(n_437), .Y(n_432) );
INVx1_ASAP7_75t_L g636 ( .A(n_68), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_70), .A2(n_95), .B1(n_425), .B2(n_586), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_71), .A2(n_150), .B1(n_622), .B2(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g773 ( .A(n_72), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_73), .A2(n_186), .B1(n_447), .B2(n_453), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_74), .A2(n_200), .B1(n_447), .B2(n_448), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g748 ( .A(n_75), .B(n_749), .C(n_753), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_75), .A2(n_753), .B1(n_758), .B2(n_1103), .Y(n_768) );
OAI21xp5_ASAP7_75t_L g769 ( .A1(n_75), .A2(n_749), .B(n_763), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_76), .A2(n_143), .B1(n_456), .B2(n_457), .Y(n_455) );
AOI21xp33_ASAP7_75t_L g464 ( .A1(n_77), .A2(n_465), .B(n_466), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_78), .A2(n_81), .B1(n_403), .B2(n_605), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_79), .A2(n_174), .B1(n_424), .B2(n_429), .Y(n_423) );
INVx1_ASAP7_75t_L g832 ( .A(n_80), .Y(n_832) );
AND2x4_ASAP7_75t_L g840 ( .A(n_80), .B(n_232), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_82), .A2(n_180), .B1(n_403), .B2(n_590), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_83), .A2(n_87), .B1(n_450), .B2(n_451), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_85), .A2(n_201), .B1(n_496), .B2(n_692), .Y(n_782) );
AOI21xp33_ASAP7_75t_L g799 ( .A1(n_86), .A2(n_537), .B(n_800), .Y(n_799) );
XNOR2x2_ASAP7_75t_L g657 ( .A(n_88), .B(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_89), .A2(n_102), .B1(n_453), .B2(n_454), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_90), .A2(n_288), .B1(n_349), .B2(n_619), .Y(n_1069) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_92), .A2(n_138), .B1(n_379), .B2(n_462), .Y(n_527) );
INVx1_ASAP7_75t_L g645 ( .A(n_94), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_96), .A2(n_218), .B1(n_488), .B2(n_489), .Y(n_776) );
INVx1_ASAP7_75t_L g830 ( .A(n_99), .Y(n_830) );
AND2x4_ASAP7_75t_L g835 ( .A(n_99), .B(n_815), .Y(n_835) );
INVx1_ASAP7_75t_SL g855 ( .A(n_99), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_100), .A2(n_304), .B1(n_542), .B2(n_543), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_101), .A2(n_103), .B1(n_425), .B2(n_586), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_104), .A2(n_286), .B1(n_492), .B2(n_493), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g591 ( .A(n_105), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_106), .A2(n_125), .B1(n_828), .B2(n_893), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_107), .A2(n_254), .B1(n_462), .B2(n_463), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_108), .A2(n_134), .B1(n_479), .B2(n_480), .Y(n_478) );
XNOR2x1_ASAP7_75t_L g793 ( .A(n_109), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g880 ( .A(n_110), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_111), .A2(n_196), .B1(n_522), .B2(n_524), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_112), .A2(n_263), .B1(n_492), .B2(n_631), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_113), .A2(n_142), .B1(n_403), .B2(n_413), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_114), .A2(n_149), .B1(n_451), .B2(n_453), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_116), .A2(n_290), .B1(n_607), .B2(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g617 ( .A(n_118), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_119), .B(n_558), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_120), .A2(n_303), .B1(n_625), .B2(n_692), .Y(n_735) );
NAND2xp33_ASAP7_75t_L g750 ( .A(n_121), .B(n_418), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_123), .A2(n_299), .B1(n_450), .B2(n_454), .Y(n_1066) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_124), .A2(n_152), .B1(n_425), .B2(n_526), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_126), .A2(n_194), .B1(n_599), .B2(n_601), .Y(n_598) );
INVx1_ASAP7_75t_L g467 ( .A(n_130), .Y(n_467) );
XNOR2x1_ASAP7_75t_L g475 ( .A(n_131), .B(n_476), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_132), .A2(n_225), .B1(n_403), .B2(n_413), .Y(n_687) );
INVx1_ASAP7_75t_L g787 ( .A(n_133), .Y(n_787) );
CKINVDCx6p67_ASAP7_75t_R g833 ( .A(n_135), .Y(n_833) );
INVx1_ASAP7_75t_L g339 ( .A(n_136), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_136), .B(n_187), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_136), .B(n_360), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_137), .B(n_242), .Y(n_395) );
AND2x2_ASAP7_75t_L g752 ( .A(n_139), .B(n_523), .Y(n_752) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_140), .A2(n_248), .B1(n_463), .B2(n_465), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_141), .A2(n_146), .B1(n_493), .B2(n_506), .Y(n_714) );
AOI21xp33_ASAP7_75t_L g666 ( .A1(n_144), .A2(n_558), .B(n_667), .Y(n_666) );
XNOR2x1_ASAP7_75t_L g518 ( .A(n_145), .B(n_519), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_151), .A2(n_284), .B1(n_858), .B2(n_859), .Y(n_863) );
INVx1_ASAP7_75t_L g1060 ( .A(n_151), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_151), .A2(n_1081), .B1(n_1083), .B2(n_1100), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_153), .A2(n_309), .B1(n_492), .B2(n_625), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_154), .B(n_389), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_155), .A2(n_179), .B1(n_542), .B2(n_543), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_156), .B(n_331), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_157), .A2(n_182), .B1(n_496), .B2(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_158), .A2(n_181), .B1(n_727), .B2(n_728), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g857 ( .A1(n_159), .A2(n_246), .B1(n_858), .B2(n_859), .Y(n_857) );
INVx1_ASAP7_75t_L g663 ( .A(n_161), .Y(n_663) );
INVx1_ASAP7_75t_L g504 ( .A(n_162), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_163), .A2(n_230), .B1(n_418), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_164), .A2(n_269), .B1(n_425), .B2(n_526), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_165), .A2(n_221), .B1(n_572), .B2(n_573), .Y(n_1094) );
INVx1_ASAP7_75t_L g837 ( .A(n_166), .Y(n_837) );
INVx1_ASAP7_75t_L g471 ( .A(n_167), .Y(n_471) );
OA22x2_ASAP7_75t_L g550 ( .A1(n_168), .A2(n_551), .B1(n_563), .B2(n_564), .Y(n_550) );
INVx1_ASAP7_75t_L g564 ( .A(n_168), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_168), .A2(n_261), .B1(n_828), .B2(n_849), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_170), .A2(n_173), .B1(n_379), .B2(n_389), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_171), .B(n_1072), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_172), .A2(n_287), .B1(n_413), .B2(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_176), .A2(n_216), .B1(n_603), .B2(n_604), .Y(n_602) );
AOI21xp33_ASAP7_75t_L g643 ( .A1(n_177), .A2(n_469), .B(n_644), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_178), .A2(n_235), .B1(n_425), .B2(n_430), .Y(n_1065) );
AOI22xp5_ASAP7_75t_L g862 ( .A1(n_183), .A2(n_294), .B1(n_854), .B2(n_856), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_184), .A2(n_240), .B1(n_843), .B2(n_867), .Y(n_891) );
AOI21x1_ASAP7_75t_SL g498 ( .A1(n_185), .A2(n_499), .B(n_503), .Y(n_498) );
INVx1_ASAP7_75t_L g343 ( .A(n_187), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_188), .A2(n_308), .B1(n_450), .B2(n_451), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_189), .A2(n_203), .B1(n_847), .B2(n_867), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_191), .A2(n_210), .B1(n_456), .B2(n_457), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_192), .A2(n_282), .B1(n_674), .B2(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g507 ( .A(n_193), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_197), .A2(n_274), .B1(n_448), .B2(n_454), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_199), .A2(n_302), .B1(n_447), .B2(n_448), .Y(n_647) );
INVx1_ASAP7_75t_L g354 ( .A(n_202), .Y(n_354) );
INVx1_ASAP7_75t_L g711 ( .A(n_205), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_206), .A2(n_215), .B1(n_447), .B2(n_463), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_207), .A2(n_271), .B1(n_640), .B2(n_761), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_208), .A2(n_296), .B1(n_590), .B2(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_209), .A2(n_300), .B1(n_572), .B2(n_680), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_211), .A2(n_276), .B1(n_496), .B2(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_212), .A2(n_228), .B1(n_828), .B2(n_849), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_213), .A2(n_278), .B1(n_413), .B2(n_417), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_217), .A2(n_233), .B1(n_584), .B2(n_586), .Y(n_686) );
INVx1_ASAP7_75t_L g539 ( .A(n_219), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_220), .B(n_570), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_222), .A2(n_250), .B1(n_402), .B2(n_408), .Y(n_401) );
AOI221xp5_ASAP7_75t_SL g557 ( .A1(n_223), .A2(n_266), .B1(n_465), .B2(n_558), .C(n_559), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g1099 ( .A1(n_226), .A2(n_305), .B1(n_403), .B2(n_728), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_227), .A2(n_239), .B1(n_482), .B2(n_483), .Y(n_777) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_229), .A2(n_253), .B1(n_627), .B2(n_629), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_231), .A2(n_247), .B1(n_839), .B2(n_847), .Y(n_846) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_232), .Y(n_817) );
AND2x4_ASAP7_75t_L g831 ( .A(n_232), .B(n_832), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_236), .A2(n_256), .B1(n_698), .B2(n_734), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_238), .A2(n_277), .B1(n_425), .B2(n_524), .Y(n_766) );
INVx1_ASAP7_75t_L g695 ( .A(n_241), .Y(n_695) );
INVx1_ASAP7_75t_L g337 ( .A(n_242), .Y(n_337) );
INVxp67_ASAP7_75t_L g388 ( .A(n_242), .Y(n_388) );
AOI21xp33_ASAP7_75t_L g736 ( .A1(n_243), .A2(n_492), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_244), .B(n_369), .Y(n_1091) );
INVxp67_ASAP7_75t_R g841 ( .A(n_249), .Y(n_841) );
INVx2_ASAP7_75t_L g815 ( .A(n_252), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_259), .A2(n_272), .B1(n_590), .B2(n_727), .Y(n_778) );
OAI22x1_ASAP7_75t_L g441 ( .A1(n_260), .A2(n_442), .B1(n_443), .B2(n_472), .Y(n_441) );
INVx1_ASAP7_75t_L g472 ( .A(n_260), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_262), .A2(n_293), .B1(n_542), .B2(n_588), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_265), .A2(n_283), .B1(n_533), .B2(n_535), .C(n_538), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_267), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_268), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_270), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g700 ( .A(n_273), .Y(n_700) );
AOI21xp33_ASAP7_75t_SL g613 ( .A1(n_275), .A2(n_614), .B(n_616), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_279), .A2(n_306), .B1(n_450), .B2(n_465), .Y(n_803) );
OAI22x1_ASAP7_75t_L g594 ( .A1(n_285), .A2(n_595), .B1(n_596), .B2(n_632), .Y(n_594) );
INVx1_ASAP7_75t_L g632 ( .A(n_285), .Y(n_632) );
AOI22x1_ASAP7_75t_L g652 ( .A1(n_285), .A2(n_595), .B1(n_596), .B2(n_632), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g1083 ( .A1(n_292), .A2(n_1084), .B1(n_1085), .B2(n_1086), .Y(n_1083) );
CKINVDCx5p33_ASAP7_75t_R g1084 ( .A(n_292), .Y(n_1084) );
INVx1_ASAP7_75t_L g373 ( .A(n_298), .Y(n_373) );
INVx1_ASAP7_75t_L g923 ( .A(n_301), .Y(n_923) );
XNOR2x1_ASAP7_75t_L g683 ( .A(n_310), .B(n_684), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g574 ( .A1(n_311), .A2(n_575), .B(n_577), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_809), .B(n_818), .Y(n_312) );
XNOR2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_545), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B1(n_513), .B2(n_544), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_473), .B(n_511), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_318), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
XNOR2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_441), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_399), .Y(n_321) );
NOR3xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_353), .C(n_372), .Y(n_322) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g698 ( .A(n_325), .Y(n_698) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g493 ( .A(n_326), .Y(n_493) );
INVx2_ASAP7_75t_L g755 ( .A(n_326), .Y(n_755) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_327), .Y(n_572) );
BUFx3_ASAP7_75t_L g631 ( .A(n_327), .Y(n_631) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_340), .Y(n_327) );
AND2x4_ASAP7_75t_L g350 ( .A(n_328), .B(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g436 ( .A(n_328), .B(n_427), .Y(n_436) );
AND2x4_ASAP7_75t_L g456 ( .A(n_328), .B(n_427), .Y(n_456) );
AND2x4_ASAP7_75t_L g462 ( .A(n_328), .B(n_340), .Y(n_462) );
AND2x4_ASAP7_75t_L g465 ( .A(n_328), .B(n_351), .Y(n_465) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_334), .Y(n_328) );
INVx2_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
AND2x2_ASAP7_75t_L g382 ( .A(n_329), .B(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g405 ( .A(n_329), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g416 ( .A(n_329), .B(n_407), .Y(n_416) );
AND2x4_ASAP7_75t_L g329 ( .A(n_330), .B(n_333), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_331), .B(n_337), .Y(n_336) );
INVxp67_ASAP7_75t_L g360 ( .A(n_331), .Y(n_360) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp33_ASAP7_75t_L g338 ( .A(n_332), .B(n_339), .Y(n_338) );
NAND2xp33_ASAP7_75t_L g342 ( .A(n_332), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g346 ( .A(n_332), .Y(n_346) );
INVx1_ASAP7_75t_L g364 ( .A(n_332), .Y(n_364) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_332), .Y(n_384) );
NAND3xp33_ASAP7_75t_L g397 ( .A(n_333), .B(n_359), .C(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g365 ( .A(n_334), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g407 ( .A(n_335), .Y(n_407) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
AND2x2_ASAP7_75t_L g377 ( .A(n_340), .B(n_365), .Y(n_377) );
AND2x2_ASAP7_75t_L g404 ( .A(n_340), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g414 ( .A(n_340), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g450 ( .A(n_340), .B(n_405), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_340), .B(n_421), .Y(n_451) );
AND2x2_ASAP7_75t_L g523 ( .A(n_340), .B(n_405), .Y(n_523) );
AND2x2_ASAP7_75t_L g537 ( .A(n_340), .B(n_365), .Y(n_537) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_347), .Y(n_340) );
INVx1_ASAP7_75t_L g352 ( .A(n_341), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_343), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g387 ( .A1(n_345), .A2(n_364), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g351 ( .A(n_347), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g386 ( .A(n_347), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g428 ( .A(n_347), .Y(n_428) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_350), .Y(n_492) );
INVx1_ASAP7_75t_L g576 ( .A(n_350), .Y(n_576) );
BUFx3_ASAP7_75t_L g628 ( .A(n_350), .Y(n_628) );
AND2x4_ASAP7_75t_L g371 ( .A(n_351), .B(n_365), .Y(n_371) );
AND2x2_ASAP7_75t_L g469 ( .A(n_351), .B(n_365), .Y(n_469) );
AND2x4_ASAP7_75t_L g427 ( .A(n_352), .B(n_428), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_367), .B2(n_368), .Y(n_353) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx3_ASAP7_75t_L g497 ( .A(n_357), .Y(n_497) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_357), .Y(n_625) );
AND2x4_ASAP7_75t_L g357 ( .A(n_358), .B(n_365), .Y(n_357) );
AND2x4_ASAP7_75t_L g411 ( .A(n_358), .B(n_405), .Y(n_411) );
AND2x4_ASAP7_75t_L g420 ( .A(n_358), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g448 ( .A(n_358), .B(n_421), .Y(n_448) );
AND2x4_ASAP7_75t_L g454 ( .A(n_358), .B(n_405), .Y(n_454) );
AND2x4_ASAP7_75t_L g470 ( .A(n_358), .B(n_365), .Y(n_470) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_363), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
AND2x2_ASAP7_75t_L g440 ( .A(n_365), .B(n_427), .Y(n_440) );
AND2x4_ASAP7_75t_L g457 ( .A(n_365), .B(n_427), .Y(n_457) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g495 ( .A(n_370), .Y(n_495) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g534 ( .A(n_371), .Y(n_534) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_371), .Y(n_558) );
BUFx3_ASAP7_75t_L g570 ( .A(n_371), .Y(n_570) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_371), .Y(n_623) );
BUFx8_ASAP7_75t_SL g692 ( .A(n_371), .Y(n_692) );
OAI21xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B(n_378), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx3_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g693 ( .A(n_376), .Y(n_693) );
INVx2_ASAP7_75t_L g1072 ( .A(n_376), .Y(n_1072) );
INVx2_ASAP7_75t_L g1090 ( .A(n_376), .Y(n_1090) );
INVx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g460 ( .A(n_377), .Y(n_460) );
INVx2_ASAP7_75t_L g502 ( .A(n_377), .Y(n_502) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g506 ( .A(n_380), .Y(n_506) );
INVx4_ASAP7_75t_L g678 ( .A(n_380), .Y(n_678) );
INVx2_ASAP7_75t_L g734 ( .A(n_380), .Y(n_734) );
INVx5_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_L g573 ( .A(n_381), .Y(n_573) );
BUFx4f_ASAP7_75t_L g619 ( .A(n_381), .Y(n_619) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_386), .Y(n_381) );
AND2x2_ASAP7_75t_L g463 ( .A(n_382), .B(n_386), .Y(n_463) );
AND2x4_ASAP7_75t_L g789 ( .A(n_382), .B(n_386), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g393 ( .A(n_384), .Y(n_393) );
INVx4_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_390), .B(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g1074 ( .A(n_390), .B(n_1075), .Y(n_1074) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx4_ASAP7_75t_L g579 ( .A(n_391), .Y(n_579) );
INVx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_392), .Y(n_510) );
AO21x2_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B(n_397), .Y(n_392) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_394), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
NOR2x1_ASAP7_75t_L g399 ( .A(n_400), .B(n_422), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_412), .Y(n_400) );
BUFx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx8_ASAP7_75t_L g486 ( .A(n_404), .Y(n_486) );
AND2x4_ASAP7_75t_L g426 ( .A(n_405), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g453 ( .A(n_405), .B(n_427), .Y(n_453) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g480 ( .A(n_410), .Y(n_480) );
INVx2_ASAP7_75t_SL g526 ( .A(n_410), .Y(n_526) );
INVx4_ASAP7_75t_L g590 ( .A(n_410), .Y(n_590) );
INVx2_ASAP7_75t_L g611 ( .A(n_410), .Y(n_611) );
INVx4_ASAP7_75t_L g675 ( .A(n_410), .Y(n_675) );
INVx4_ASAP7_75t_L g706 ( .A(n_410), .Y(n_706) );
INVx2_ASAP7_75t_L g728 ( .A(n_410), .Y(n_728) );
INVx8_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_414), .Y(n_524) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_414), .Y(n_583) );
BUFx12f_ASAP7_75t_L g605 ( .A(n_414), .Y(n_605) );
AND2x4_ASAP7_75t_L g447 ( .A(n_415), .B(n_427), .Y(n_447) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g421 ( .A(n_416), .Y(n_421) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx5_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx3_ASAP7_75t_L g584 ( .A(n_419), .Y(n_584) );
INVx2_ASAP7_75t_L g1064 ( .A(n_419), .Y(n_1064) );
INVx6_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx12f_ASAP7_75t_L g483 ( .A(n_420), .Y(n_483) );
AND2x4_ASAP7_75t_L g431 ( .A(n_421), .B(n_427), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_432), .Y(n_422) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx12f_ASAP7_75t_L g479 ( .A(n_425), .Y(n_479) );
BUFx12f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_426), .Y(n_674) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_426), .Y(n_727) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g600 ( .A(n_430), .Y(n_600) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_431), .Y(n_482) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_431), .Y(n_531) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_431), .Y(n_586) );
BUFx4f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g588 ( .A(n_435), .Y(n_588) );
INVx1_ASAP7_75t_L g607 ( .A(n_435), .Y(n_607) );
INVx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_436), .Y(n_488) );
BUFx12f_ASAP7_75t_L g543 ( .A(n_436), .Y(n_543) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx5_ASAP7_75t_L g489 ( .A(n_440), .Y(n_489) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_440), .Y(n_542) );
BUFx3_ASAP7_75t_L g765 ( .A(n_440), .Y(n_765) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
XOR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_471), .Y(n_443) );
NOR2xp67_ASAP7_75t_L g444 ( .A(n_445), .B(n_458), .Y(n_444) );
NAND4xp25_ASAP7_75t_L g445 ( .A(n_446), .B(n_449), .C(n_452), .D(n_455), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .C(n_464), .D(n_468), .Y(n_458) );
BUFx3_ASAP7_75t_L g615 ( .A(n_460), .Y(n_615) );
INVx2_ASAP7_75t_L g785 ( .A(n_460), .Y(n_785) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g512 ( .A(n_475), .Y(n_512) );
NAND4xp75_ASAP7_75t_SL g476 ( .A(n_477), .B(n_484), .C(n_490), .D(n_498), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_481), .Y(n_477) );
BUFx3_ASAP7_75t_L g601 ( .A(n_483), .Y(n_601) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_494), .Y(n_490) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g680 ( .A(n_497), .Y(n_680) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g665 ( .A(n_501), .Y(n_665) );
INVx2_ASAP7_75t_L g732 ( .A(n_501), .Y(n_732) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g640 ( .A(n_502), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B1(n_507), .B2(n_508), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_510), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_510), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g670 ( .A(n_510), .Y(n_670) );
INVx1_ASAP7_75t_L g740 ( .A(n_510), .Y(n_740) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_510), .Y(n_762) );
INVx1_ASAP7_75t_L g544 ( .A(n_513), .Y(n_544) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NOR2x1_ASAP7_75t_L g519 ( .A(n_520), .B(n_529), .Y(n_519) );
NAND4xp25_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .C(n_527), .D(n_528), .Y(n_520) );
BUFx4f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_523), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .C(n_541), .Y(n_529) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
BUFx2_ASAP7_75t_SL g608 ( .A(n_542), .Y(n_608) );
XNOR2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_654), .Y(n_545) );
XOR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_593), .Y(n_546) );
BUFx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OA22x2_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_565), .B1(n_566), .B2(n_592), .Y(n_549) );
INVx2_ASAP7_75t_L g592 ( .A(n_550), .Y(n_592) );
INVx1_ASAP7_75t_L g563 ( .A(n_551), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_557), .C(n_561), .Y(n_551) );
AND4x1_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .C(n_555), .D(n_556), .Y(n_552) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
XNOR2x1_ASAP7_75t_L g566 ( .A(n_567), .B(n_591), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_581), .Y(n_567) );
NAND4xp25_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .C(n_574), .D(n_580), .Y(n_568) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g1093 ( .A(n_576), .Y(n_1093) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_579), .B(n_645), .Y(n_644) );
INVx4_ASAP7_75t_L g713 ( .A(n_579), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_579), .B(n_801), .Y(n_800) );
NAND4xp25_ASAP7_75t_L g581 ( .A(n_582), .B(n_585), .C(n_587), .D(n_589), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_591), .A2(n_827), .B1(n_833), .B2(n_834), .Y(n_826) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_633), .B1(n_652), .B2(n_653), .Y(n_593) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_612), .Y(n_596) );
NAND4xp25_ASAP7_75t_SL g597 ( .A(n_598), .B(n_602), .C(n_606), .D(n_609), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_621), .C(n_626), .Y(n_612) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI21xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B(n_620), .Y(n_616) );
INVx2_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
BUFx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_632), .A2(n_834), .B1(n_879), .B2(n_880), .Y(n_878) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g653 ( .A(n_635), .Y(n_653) );
AO21x2_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B(n_651), .Y(n_635) );
NOR3xp33_ASAP7_75t_SL g651 ( .A(n_636), .B(n_638), .C(n_646), .Y(n_651) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_646), .Y(n_637) );
NAND4xp75_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .C(n_642), .D(n_643), .Y(n_638) );
NAND4xp25_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .C(n_649), .D(n_650), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B1(n_716), .B2(n_717), .Y(n_654) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
XNOR2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_681), .Y(n_656) );
NAND4xp75_ASAP7_75t_L g658 ( .A(n_659), .B(n_662), .C(n_671), .D(n_676), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
OA21x2_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_669), .B(n_695), .Y(n_694) );
INVx3_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVxp67_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
XNOR2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_699), .Y(n_682) );
NOR2x1_ASAP7_75t_L g684 ( .A(n_685), .B(n_690), .Y(n_684) );
NAND4xp25_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .C(n_688), .D(n_689), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_696), .C(n_697), .Y(n_690) );
XNOR2x1_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
NOR2x1_ASAP7_75t_L g701 ( .A(n_702), .B(n_708), .Y(n_701) );
NAND4xp25_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .C(n_705), .D(n_707), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_714), .C(n_715), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_770), .B1(n_771), .B2(n_808), .Y(n_717) );
INVx1_ASAP7_75t_L g808 ( .A(n_718), .Y(n_808) );
INVx2_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
XOR2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_747), .Y(n_719) );
OAI21xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B(n_741), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_721), .B(n_733), .Y(n_744) );
NOR2xp67_ASAP7_75t_L g722 ( .A(n_723), .B(n_730), .Y(n_722) );
INVx1_ASAP7_75t_L g742 ( .A(n_723), .Y(n_742) );
NAND4xp25_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .C(n_726), .D(n_729), .Y(n_723) );
NAND4xp25_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .C(n_735), .D(n_736), .Y(n_730) );
INVx1_ASAP7_75t_L g745 ( .A(n_731), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_735), .B(n_736), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .C(n_746), .Y(n_743) );
AO21x2_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_757), .B(n_767), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g753 ( .A(n_754), .B(n_756), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_763), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND2x1_ASAP7_75t_SL g763 ( .A(n_764), .B(n_766), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OA22x2_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_791), .B1(n_792), .B2(n_807), .Y(n_771) );
INVx1_ASAP7_75t_L g807 ( .A(n_772), .Y(n_807) );
XNOR2x1_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
NOR2x1_ASAP7_75t_L g774 ( .A(n_775), .B(n_780), .Y(n_774) );
NAND4xp25_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .C(n_778), .D(n_779), .Y(n_775) );
NAND3xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .C(n_783), .Y(n_780) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
OAI21xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_788), .B(n_790), .Y(n_786) );
INVx4_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NOR2x1_ASAP7_75t_L g794 ( .A(n_795), .B(n_802), .Y(n_794) );
NAND4xp25_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .C(n_798), .D(n_799), .Y(n_795) );
NAND4xp25_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .C(n_805), .D(n_806), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
BUFx10_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NAND3xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_816), .C(n_817), .Y(n_812) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_813), .B(n_1078), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_813), .B(n_1079), .Y(n_1082) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
OA21x2_ASAP7_75t_L g1100 ( .A1(n_814), .A2(n_855), .B(n_1101), .Y(n_1100) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g829 ( .A(n_815), .B(n_830), .Y(n_829) );
AND3x4_ASAP7_75t_L g854 ( .A(n_815), .B(n_831), .C(n_855), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g1078 ( .A(n_816), .B(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_817), .Y(n_1079) );
OAI221xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_1051), .B1(n_1053), .B2(n_1076), .C(n_1080), .Y(n_818) );
AOI211xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_964), .B(n_1012), .C(n_1037), .Y(n_819) );
NAND5xp2_ASAP7_75t_L g820 ( .A(n_821), .B(n_899), .C(n_928), .D(n_937), .E(n_957), .Y(n_820) );
NOR3xp33_ASAP7_75t_SL g821 ( .A(n_822), .B(n_869), .C(n_887), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_824), .B(n_850), .Y(n_823) );
INVx1_ASAP7_75t_L g949 ( .A(n_824), .Y(n_949) );
AOI221xp5_ASAP7_75t_L g965 ( .A1(n_824), .A2(n_966), .B1(n_968), .B2(n_969), .C(n_970), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_824), .B(n_896), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_824), .B(n_876), .Y(n_1031) );
AND2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_844), .Y(n_824) );
AND2x2_ASAP7_75t_L g886 ( .A(n_825), .B(n_845), .Y(n_886) );
INVx2_ASAP7_75t_L g903 ( .A(n_825), .Y(n_903) );
INVx3_ASAP7_75t_L g910 ( .A(n_825), .Y(n_910) );
OR2x2_ASAP7_75t_L g939 ( .A(n_825), .B(n_845), .Y(n_939) );
NOR2xp33_ASAP7_75t_L g956 ( .A(n_825), .B(n_877), .Y(n_956) );
OR2x2_ASAP7_75t_L g825 ( .A(n_826), .B(n_836), .Y(n_825) );
OAI221xp5_ASAP7_75t_L g921 ( .A1(n_827), .A2(n_834), .B1(n_922), .B2(n_923), .C(n_924), .Y(n_921) );
INVx3_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AND2x4_ASAP7_75t_L g828 ( .A(n_829), .B(n_831), .Y(n_828) );
AND2x4_ASAP7_75t_L g839 ( .A(n_829), .B(n_840), .Y(n_839) );
AND2x2_ASAP7_75t_L g858 ( .A(n_829), .B(n_840), .Y(n_858) );
AND2x2_ASAP7_75t_L g867 ( .A(n_829), .B(n_840), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_831), .B(n_835), .Y(n_834) );
AND2x4_ASAP7_75t_L g849 ( .A(n_831), .B(n_835), .Y(n_849) );
AND2x4_ASAP7_75t_L g856 ( .A(n_831), .B(n_835), .Y(n_856) );
AND2x4_ASAP7_75t_L g843 ( .A(n_835), .B(n_840), .Y(n_843) );
AND2x2_ASAP7_75t_L g847 ( .A(n_835), .B(n_840), .Y(n_847) );
AND2x2_ASAP7_75t_L g859 ( .A(n_835), .B(n_840), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B1(n_841), .B2(n_842), .Y(n_836) );
INVx3_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g1101 ( .A(n_840), .Y(n_1101) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
BUFx2_ASAP7_75t_L g1052 ( .A(n_843), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_844), .B(n_889), .Y(n_888) );
INVx3_ASAP7_75t_L g919 ( .A(n_844), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_844), .B(n_890), .Y(n_1029) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_844), .B(n_890), .Y(n_1050) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
AND2x2_ASAP7_75t_L g909 ( .A(n_845), .B(n_910), .Y(n_909) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_845), .B(n_890), .Y(n_1025) );
AND2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_848), .Y(n_845) );
O2A1O1Ixp33_ASAP7_75t_L g973 ( .A1(n_850), .A2(n_963), .B(n_974), .C(n_976), .Y(n_973) );
AOI222xp33_ASAP7_75t_L g1022 ( .A1(n_850), .A2(n_1023), .B1(n_1025), .B2(n_1026), .C1(n_1027), .C2(n_1030), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_850), .B(n_876), .Y(n_1024) );
AND2x2_ASAP7_75t_L g850 ( .A(n_851), .B(n_860), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_851), .B(n_871), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_851), .B(n_873), .Y(n_931) );
AND2x2_ASAP7_75t_SL g936 ( .A(n_851), .B(n_906), .Y(n_936) );
NOR2xp33_ASAP7_75t_L g960 ( .A(n_851), .B(n_961), .Y(n_960) );
AND2x2_ASAP7_75t_L g967 ( .A(n_851), .B(n_876), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_851), .B(n_877), .Y(n_986) );
AND2x2_ASAP7_75t_L g998 ( .A(n_851), .B(n_864), .Y(n_998) );
A2O1A1Ixp33_ASAP7_75t_L g1032 ( .A1(n_851), .A2(n_1033), .B(n_1034), .C(n_1035), .Y(n_1032) );
CKINVDCx6p67_ASAP7_75t_R g851 ( .A(n_852), .Y(n_851) );
AND2x2_ASAP7_75t_L g898 ( .A(n_852), .B(n_860), .Y(n_898) );
AND2x2_ASAP7_75t_L g905 ( .A(n_852), .B(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g914 ( .A(n_852), .Y(n_914) );
OR2x2_ASAP7_75t_L g983 ( .A(n_852), .B(n_861), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_852), .B(n_873), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_852), .B(n_968), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_852), .B(n_861), .Y(n_1042) );
AND2x2_ASAP7_75t_L g852 ( .A(n_853), .B(n_857), .Y(n_852) );
INVx1_ASAP7_75t_L g879 ( .A(n_854), .Y(n_879) );
INVx2_ASAP7_75t_SL g894 ( .A(n_856), .Y(n_894) );
INVx1_ASAP7_75t_L g885 ( .A(n_858), .Y(n_885) );
INVx1_ASAP7_75t_L g883 ( .A(n_859), .Y(n_883) );
INVx1_ASAP7_75t_L g1010 ( .A(n_860), .Y(n_1010) );
OR2x2_ASAP7_75t_L g1033 ( .A(n_860), .B(n_906), .Y(n_1033) );
AND2x2_ASAP7_75t_L g860 ( .A(n_861), .B(n_864), .Y(n_860) );
AND2x2_ASAP7_75t_L g871 ( .A(n_861), .B(n_865), .Y(n_871) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_861), .Y(n_874) );
AND2x4_ASAP7_75t_SL g861 ( .A(n_862), .B(n_863), .Y(n_861) );
AND2x2_ASAP7_75t_L g873 ( .A(n_864), .B(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g912 ( .A(n_864), .Y(n_912) );
NOR2xp33_ASAP7_75t_L g940 ( .A(n_864), .B(n_913), .Y(n_940) );
AND2x2_ASAP7_75t_L g955 ( .A(n_864), .B(n_913), .Y(n_955) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
AND2x2_ASAP7_75t_L g906 ( .A(n_865), .B(n_874), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_868), .Y(n_865) );
AOI21xp33_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_872), .B(n_875), .Y(n_869) );
INVx1_ASAP7_75t_L g1018 ( .A(n_870), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_870), .B(n_1045), .Y(n_1044) );
AND2x2_ASAP7_75t_L g951 ( .A(n_871), .B(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g961 ( .A(n_871), .Y(n_961) );
AND2x2_ASAP7_75t_L g968 ( .A(n_871), .B(n_877), .Y(n_968) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_871), .B(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
AND2x2_ASAP7_75t_L g947 ( .A(n_873), .B(n_877), .Y(n_947) );
OAI321xp33_ASAP7_75t_L g985 ( .A1(n_873), .A2(n_911), .A3(n_950), .B1(n_984), .B2(n_986), .C(n_987), .Y(n_985) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_873), .B(n_952), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_874), .B(n_913), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_876), .B(n_886), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g916 ( .A(n_876), .B(n_917), .Y(n_916) );
AND2x2_ASAP7_75t_L g952 ( .A(n_876), .B(n_913), .Y(n_952) );
NOR2x1p5_ASAP7_75t_L g982 ( .A(n_876), .B(n_983), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_876), .B(n_919), .Y(n_996) );
INVx1_ASAP7_75t_L g1007 ( .A(n_876), .Y(n_1007) );
NOR2xp33_ASAP7_75t_L g1048 ( .A(n_876), .B(n_910), .Y(n_1048) );
CKINVDCx6p67_ASAP7_75t_R g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g897 ( .A(n_877), .Y(n_897) );
AND2x2_ASAP7_75t_L g904 ( .A(n_877), .B(n_905), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_877), .B(n_940), .Y(n_975) );
NOR2xp33_ASAP7_75t_L g988 ( .A(n_877), .B(n_910), .Y(n_988) );
NOR2xp33_ASAP7_75t_L g1009 ( .A(n_877), .B(n_1010), .Y(n_1009) );
OR2x6_ASAP7_75t_SL g877 ( .A(n_878), .B(n_881), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_882), .A2(n_883), .B1(n_884), .B2(n_885), .Y(n_881) );
INVx1_ASAP7_75t_L g971 ( .A(n_886), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_886), .B(n_890), .Y(n_1036) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_895), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_888), .B(n_896), .Y(n_929) );
INVx1_ASAP7_75t_L g1043 ( .A(n_888), .Y(n_1043) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_889), .B(n_927), .Y(n_926) );
INVx2_ASAP7_75t_L g944 ( .A(n_889), .Y(n_944) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_889), .Y(n_989) );
INVx3_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g933 ( .A(n_890), .Y(n_933) );
AND2x2_ASAP7_75t_L g963 ( .A(n_890), .B(n_938), .Y(n_963) );
AND2x4_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
INVx2_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_896), .B(n_898), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_896), .B(n_909), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_896), .B(n_936), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_896), .B(n_955), .Y(n_1017) );
INVx3_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g1045 ( .A(n_898), .Y(n_1045) );
OAI21xp33_ASAP7_75t_L g899 ( .A1(n_900), .A2(n_907), .B(n_925), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_904), .Y(n_901) );
INVx2_ASAP7_75t_L g969 ( .A(n_902), .Y(n_969) );
BUFx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_903), .B(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g992 ( .A(n_903), .Y(n_992) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_903), .B(n_1020), .Y(n_1019) );
NOR2xp33_ASAP7_75t_L g1041 ( .A(n_903), .B(n_1042), .Y(n_1041) );
AND2x2_ASAP7_75t_L g966 ( .A(n_906), .B(n_967), .Y(n_966) );
OAI221xp5_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_911), .B1(n_915), .B2(n_918), .C(n_920), .Y(n_907) );
INVx1_ASAP7_75t_L g999 ( .A(n_909), .Y(n_999) );
O2A1O1Ixp33_ASAP7_75t_L g1013 ( .A1(n_909), .A2(n_1014), .B(n_1018), .C(n_1019), .Y(n_1013) );
INVx1_ASAP7_75t_L g981 ( .A(n_910), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_910), .B(n_944), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_910), .B(n_951), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_911), .B(n_931), .Y(n_930) );
NOR2xp33_ASAP7_75t_L g976 ( .A(n_911), .B(n_977), .Y(n_976) );
O2A1O1Ixp33_ASAP7_75t_L g1005 ( .A1(n_911), .A2(n_1006), .B(n_1008), .C(n_1011), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_912), .B(n_913), .Y(n_911) );
AND2x2_ASAP7_75t_L g993 ( .A(n_913), .B(n_947), .Y(n_993) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g1015 ( .A(n_916), .B(n_1016), .Y(n_1015) );
OAI22xp33_ASAP7_75t_L g995 ( .A1(n_917), .A2(n_996), .B1(n_997), .B2(n_999), .Y(n_995) );
NOR2xp33_ASAP7_75t_L g953 ( .A(n_918), .B(n_954), .Y(n_953) );
OAI221xp5_ASAP7_75t_L g970 ( .A1(n_918), .A2(n_927), .B1(n_959), .B2(n_971), .C(n_972), .Y(n_970) );
INVx3_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_919), .A2(n_946), .B1(n_948), .B2(n_950), .Y(n_945) );
INVx1_ASAP7_75t_L g984 ( .A(n_919), .Y(n_984) );
OAI221xp5_ASAP7_75t_L g1037 ( .A1(n_919), .A2(n_942), .B1(n_1038), .B2(n_1039), .C(n_1040), .Y(n_1037) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
BUFx3_ASAP7_75t_L g927 ( .A(n_921), .Y(n_927) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_930), .B1(n_932), .B2(n_934), .Y(n_928) );
INVx1_ASAP7_75t_L g1011 ( .A(n_932), .Y(n_1011) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
AOI311xp33_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_940), .A3(n_941), .B(n_945), .C(n_953), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_940), .B(n_956), .Y(n_972) );
OAI211xp5_ASAP7_75t_L g1012 ( .A1(n_941), .A2(n_1013), .B(n_1022), .C(n_1032), .Y(n_1012) );
INVx3_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_942), .B(n_949), .Y(n_948) );
INVx3_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_943), .B(n_1048), .Y(n_1047) );
INVx3_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_951), .B(n_992), .Y(n_1039) );
AOI21xp33_ASAP7_75t_L g1049 ( .A1(n_954), .A2(n_1002), .B(n_1050), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_955), .B(n_956), .Y(n_954) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_959), .B(n_962), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
NAND5xp2_ASAP7_75t_L g964 ( .A(n_965), .B(n_973), .C(n_978), .D(n_990), .E(n_994), .Y(n_964) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_977), .B(n_1047), .Y(n_1046) );
A2O1A1Ixp33_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_984), .B(n_985), .C(n_989), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_981), .B(n_982), .Y(n_980) );
INVx1_ASAP7_75t_L g1021 ( .A(n_986), .Y(n_1021) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g1000 ( .A(n_989), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_991), .B(n_993), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_992), .B(n_1028), .Y(n_1027) );
AOI221xp5_ASAP7_75t_L g994 ( .A1(n_995), .A2(n_1000), .B1(n_1001), .B2(n_1003), .C(n_1005), .Y(n_994) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
CKINVDCx14_ASAP7_75t_R g1006 ( .A(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVxp67_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
AOI221xp5_ASAP7_75t_L g1040 ( .A1(n_1041), .A2(n_1043), .B1(n_1044), .B2(n_1046), .C(n_1049), .Y(n_1040) );
CKINVDCx5p33_ASAP7_75t_R g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVxp67_ASAP7_75t_SL g1057 ( .A(n_1058), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
XNOR2x1_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1061), .Y(n_1059) );
NOR2x1_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1068), .Y(n_1061) );
NAND4xp25_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1065), .C(n_1066), .D(n_1067), .Y(n_1062) );
NAND4xp25_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1070), .C(n_1071), .D(n_1073), .Y(n_1068) );
CKINVDCx16_ASAP7_75t_R g1076 ( .A(n_1077), .Y(n_1076) );
BUFx2_ASAP7_75t_SL g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
HB1xp67_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
NOR2x1_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1095), .Y(n_1087) );
NAND4xp25_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1091), .C(n_1092), .D(n_1094), .Y(n_1088) );
NAND4xp25_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1097), .C(n_1098), .D(n_1099), .Y(n_1095) );
endmodule