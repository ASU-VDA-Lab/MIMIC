module fake_jpeg_1952_n_249 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_218;
wire n_63;
wire n_92;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_1),
.B(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_8),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_50),
.Y(n_72)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_59),
.Y(n_82)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_20),
.B(n_21),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_0),
.Y(n_88)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_64),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_29),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_33),
.Y(n_66)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_65),
.B(n_3),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_66),
.B(n_88),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_98),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_36),
.B1(n_35),
.B2(n_17),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_84),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_25),
.B1(n_17),
.B2(n_31),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_62),
.B1(n_43),
.B2(n_57),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_83),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_24),
.B1(n_31),
.B2(n_27),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_41),
.A2(n_27),
.B1(n_24),
.B2(n_25),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_37),
.B1(n_23),
.B2(n_21),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_100),
.B1(n_57),
.B2(n_7),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_23),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_7),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_5),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_39),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_5),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_95),
.B(n_42),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_47),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_49),
.A2(n_6),
.B1(n_7),
.B2(n_12),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_102),
.B(n_104),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_103),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_52),
.C(n_48),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_71),
.Y(n_135)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_118),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_45),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_70),
.B(n_15),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_12),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_123),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_13),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_14),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_127),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_77),
.B(n_57),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_93),
.Y(n_142)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_80),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_132),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_142),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_107),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_102),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_89),
.B1(n_101),
.B2(n_71),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_141),
.A2(n_153),
.B1(n_158),
.B2(n_112),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_96),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_108),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_105),
.A2(n_128),
.B1(n_110),
.B2(n_120),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_121),
.A2(n_89),
.B1(n_101),
.B2(n_96),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_127),
.B1(n_106),
.B2(n_114),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_171),
.B1(n_141),
.B2(n_158),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_160),
.B(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_135),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_163),
.C(n_167),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_117),
.C(n_113),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_165),
.A2(n_151),
.B1(n_134),
.B2(n_150),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_116),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_177),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_118),
.C(n_122),
.Y(n_170)
);

OAI21x1_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_172),
.B(n_148),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_114),
.B1(n_119),
.B2(n_115),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_129),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_174),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_124),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_86),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_136),
.A2(n_81),
.B1(n_93),
.B2(n_86),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_90),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_183),
.A2(n_197),
.B1(n_171),
.B2(n_178),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_185),
.B(n_194),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_150),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_186),
.A2(n_136),
.B(n_90),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_151),
.B(n_144),
.C(n_152),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_195),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_193),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_170),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_157),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_174),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_198),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_145),
.C(n_149),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_204),
.A2(n_211),
.B(n_212),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_205),
.B(n_209),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_163),
.B1(n_164),
.B2(n_168),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_183),
.A2(n_145),
.B1(n_156),
.B2(n_149),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_190),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_184),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_138),
.Y(n_211)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_186),
.C(n_187),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_220),
.C(n_221),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_191),
.C(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_195),
.C(n_189),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_200),
.B1(n_206),
.B2(n_187),
.Y(n_223)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_207),
.B1(n_201),
.B2(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_229),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_199),
.B(n_212),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_225),
.B(n_227),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_204),
.C(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_218),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_228),
.B(n_214),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_235),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_219),
.C(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_227),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_226),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_232),
.B(n_138),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_241),
.A2(n_234),
.B1(n_136),
.B2(n_81),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_125),
.Y(n_245)
);

AOI221xp5_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_246),
.B1(n_243),
.B2(n_74),
.C(n_92),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_237),
.C(n_103),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_68),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_248),
.B(n_92),
.Y(n_249)
);


endmodule