module fake_jpeg_18828_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx10_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

HAxp5_ASAP7_75t_SL g12 ( 
.A(n_5),
.B(n_1),
.CON(n_12),
.SN(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_16),
.B(n_24),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_SL g18 ( 
.A(n_7),
.B(n_4),
.C(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_22),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_19)
);

OAI22x1_ASAP7_75t_L g31 ( 
.A1(n_19),
.A2(n_10),
.B1(n_13),
.B2(n_9),
.Y(n_31)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_14),
.B1(n_10),
.B2(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_11),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_12),
.C(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_24),
.Y(n_33)
);

BUFx12f_ASAP7_75t_SL g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_38),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_16),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_10),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_31),
.B1(n_28),
.B2(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_42),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_17),
.B1(n_20),
.B2(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_46),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

NOR4xp25_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_43),
.C(n_29),
.D(n_23),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_47),
.B(n_36),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_49),
.C(n_47),
.Y(n_51)
);


endmodule