module fake_jpeg_12863_n_574 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_574);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_574;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_53),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_55),
.B(n_69),
.Y(n_126)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_56),
.Y(n_149)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_64),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_68),
.B(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_18),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_28),
.B(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_72),
.B(n_83),
.Y(n_140)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_87),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_77),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_32),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_34),
.B(n_49),
.Y(n_113)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_34),
.A2(n_16),
.B(n_14),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_28),
.B(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_86),
.B(n_48),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_31),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_93),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_96),
.Y(n_109)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_24),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

INVx11_ASAP7_75t_SL g106 ( 
.A(n_33),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_36),
.B1(n_33),
.B2(n_37),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_107),
.A2(n_70),
.B1(n_89),
.B2(n_75),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_106),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_112),
.B(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_113),
.A2(n_47),
.B1(n_46),
.B2(n_45),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_81),
.A2(n_36),
.B1(n_49),
.B2(n_41),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_116),
.A2(n_123),
.B(n_167),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_56),
.A2(n_50),
.B(n_39),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_118),
.B(n_165),
.Y(n_213)
);

INVx2_ASAP7_75t_R g121 ( 
.A(n_85),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_121),
.B(n_54),
.Y(n_205)
);

INVx6_ASAP7_75t_SL g122 ( 
.A(n_79),
.Y(n_122)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_122),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_63),
.A2(n_52),
.B1(n_49),
.B2(n_41),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_41),
.C(n_52),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_124),
.B(n_48),
.C(n_39),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_34),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_134),
.B(n_136),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_59),
.B(n_25),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_90),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_163),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_92),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_61),
.B(n_25),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_94),
.B(n_24),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_168),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_71),
.A2(n_42),
.B1(n_38),
.B2(n_37),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_171),
.Y(n_269)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_173),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_177),
.Y(n_287)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_179),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_116),
.A2(n_84),
.B1(n_67),
.B2(n_78),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_180),
.A2(n_232),
.B1(n_100),
.B2(n_101),
.Y(n_265)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_126),
.B(n_94),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_182),
.B(n_185),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_183),
.B(n_188),
.Y(n_238)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_184),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_46),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_186),
.Y(n_270)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_187),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_158),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_109),
.A2(n_73),
.B1(n_37),
.B2(n_22),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_189),
.Y(n_279)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_190),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_191),
.A2(n_196),
.B1(n_151),
.B2(n_143),
.Y(n_283)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_192),
.Y(n_286)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_133),
.Y(n_193)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_193),
.Y(n_273)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_194),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_107),
.A2(n_77),
.B1(n_104),
.B2(n_95),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_196),
.A2(n_169),
.B1(n_160),
.B2(n_151),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_43),
.C(n_26),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_40),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_198),
.B(n_206),
.Y(n_252)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_135),
.Y(n_200)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_200),
.Y(n_276)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_201),
.Y(n_267)
);

BUFx4f_ASAP7_75t_SL g202 ( 
.A(n_149),
.Y(n_202)
);

INVx13_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_109),
.A2(n_22),
.B1(n_38),
.B2(n_42),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_203),
.A2(n_212),
.B1(n_215),
.B2(n_222),
.Y(n_242)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_138),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_204),
.B(n_207),
.Y(n_256)
);

NAND2xp33_ASAP7_75t_SL g243 ( 
.A(n_205),
.B(n_43),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_40),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_211),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_141),
.Y(n_209)
);

INVx13_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_210),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_111),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_152),
.A2(n_22),
.B1(n_38),
.B2(n_42),
.Y(n_212)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_214),
.B(n_217),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_154),
.A2(n_39),
.B1(n_50),
.B2(n_96),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_118),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_216),
.B(n_218),
.Y(n_277)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_120),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_130),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_219),
.B(n_220),
.Y(n_284)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_120),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_147),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_221),
.B(n_226),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_128),
.A2(n_50),
.B1(n_97),
.B2(n_98),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_170),
.A2(n_105),
.B1(n_102),
.B2(n_88),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_223),
.A2(n_167),
.B(n_123),
.Y(n_237)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_128),
.Y(n_224)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_128),
.Y(n_225)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_108),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_127),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_227),
.Y(n_246)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_146),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_229),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_145),
.B(n_47),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_230),
.B(n_114),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_143),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_231),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_110),
.B1(n_162),
.B2(n_161),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_234),
.A2(n_247),
.B1(n_214),
.B2(n_178),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_237),
.A2(n_243),
.B(n_191),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_195),
.B(n_205),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_240),
.A2(n_241),
.B(n_262),
.C(n_228),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_121),
.B(n_45),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_199),
.A2(n_110),
.B1(n_162),
.B2(n_161),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_248),
.B(n_271),
.C(n_280),
.Y(n_292)
);

NAND2x1_ASAP7_75t_L g249 ( 
.A(n_195),
.B(n_108),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_249),
.Y(n_289)
);

AOI32xp33_ASAP7_75t_L g250 ( 
.A1(n_176),
.A2(n_26),
.A3(n_129),
.B1(n_125),
.B2(n_117),
.Y(n_250)
);

AOI32xp33_ASAP7_75t_L g312 ( 
.A1(n_250),
.A2(n_228),
.A3(n_177),
.B1(n_211),
.B2(n_231),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_259),
.A2(n_283),
.B1(n_2),
.B2(n_3),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_197),
.A2(n_117),
.B(n_114),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_174),
.B(n_0),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_263),
.B(n_268),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_193),
.B(n_129),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_175),
.B(n_125),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_282),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_223),
.B(n_1),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_200),
.B(n_169),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_204),
.B(n_160),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_282),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_236),
.B(n_202),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_288),
.B(n_290),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_238),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_291),
.Y(n_353)
);

OR2x2_ASAP7_75t_SL g293 ( 
.A(n_240),
.B(n_192),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_293),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_295),
.A2(n_316),
.B(n_281),
.Y(n_372)
);

BUFx8_ASAP7_75t_L g296 ( 
.A(n_239),
.Y(n_296)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_296),
.Y(n_368)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_297),
.Y(n_363)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_298),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_236),
.B(n_202),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_299),
.B(n_301),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_300),
.B(n_304),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_256),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_245),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_233),
.B(n_219),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_303),
.B(n_309),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_173),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_262),
.B(n_207),
.C(n_229),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_281),
.C(n_260),
.Y(n_342)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_306),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_249),
.A2(n_209),
.B(n_217),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_307),
.A2(n_286),
.B(n_281),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_254),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_329),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_233),
.B(n_187),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_311),
.B(n_315),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_312),
.A2(n_328),
.B1(n_286),
.B2(n_269),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_279),
.A2(n_224),
.B1(n_225),
.B2(n_177),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_314),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_248),
.B(n_190),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_279),
.A2(n_180),
.B1(n_211),
.B2(n_220),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_235),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_323),
.Y(n_344)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_244),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_318),
.B(n_319),
.Y(n_378)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_244),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_265),
.A2(n_201),
.B1(n_227),
.B2(n_231),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_320),
.B(n_321),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_237),
.A2(n_227),
.B1(n_171),
.B2(n_3),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_249),
.B(n_1),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_322),
.B(n_330),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_235),
.Y(n_324)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_324),
.Y(n_354)
);

AND2x6_ASAP7_75t_L g325 ( 
.A(n_251),
.B(n_11),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_327),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_252),
.B(n_2),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_326),
.B(n_334),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g327 ( 
.A(n_277),
.B(n_11),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_266),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_241),
.B(n_2),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_271),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_332),
.B(n_333),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_255),
.B(n_11),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_263),
.B(n_4),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_271),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_335),
.B(n_336),
.Y(n_365)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_266),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g337 ( 
.A(n_243),
.B(n_4),
.CI(n_5),
.CON(n_337),
.SN(n_337)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_337),
.B(n_287),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_292),
.B(n_280),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_338),
.B(n_340),
.C(n_342),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_292),
.B(n_270),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_308),
.A2(n_242),
.B1(n_259),
.B2(n_270),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_341),
.B(n_366),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_304),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_343),
.B(n_339),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_256),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_345),
.B(n_348),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_294),
.B(n_256),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_356),
.A2(n_307),
.B(n_322),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_362),
.A2(n_379),
.B(n_295),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_364),
.A2(n_310),
.B1(n_327),
.B2(n_337),
.Y(n_408)
);

OAI32xp33_ASAP7_75t_L g366 ( 
.A1(n_294),
.A2(n_273),
.A3(n_276),
.B1(n_257),
.B2(n_278),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_289),
.B(n_295),
.C(n_291),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_295),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_371),
.B(n_380),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_372),
.A2(n_375),
.B(n_380),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_300),
.Y(n_373)
);

INVx13_ASAP7_75t_L g419 ( 
.A(n_373),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_308),
.A2(n_253),
.B1(n_260),
.B2(n_276),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_376),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_289),
.A2(n_287),
.B(n_246),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_328),
.A2(n_253),
.B1(n_273),
.B2(n_261),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_316),
.A2(n_257),
.B1(n_267),
.B2(n_264),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_320),
.Y(n_400)
);

OA21x2_ASAP7_75t_L g379 ( 
.A1(n_321),
.A2(n_267),
.B(n_245),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_293),
.A2(n_246),
.B(n_264),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_403),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_355),
.B(n_309),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_383),
.B(n_388),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_385),
.A2(n_384),
.B(n_375),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_368),
.Y(n_386)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_386),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_387),
.B(n_389),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_378),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_331),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_363),
.Y(n_390)
);

BUFx5_ASAP7_75t_L g442 ( 
.A(n_390),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_360),
.B(n_333),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_391),
.B(n_392),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_347),
.B(n_323),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_344),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_393),
.B(n_402),
.Y(n_446)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_363),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_395),
.Y(n_436)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_396),
.Y(n_429)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_359),
.Y(n_397)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_373),
.A2(n_335),
.B1(n_332),
.B2(n_302),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_399),
.A2(n_367),
.B1(n_372),
.B2(n_369),
.Y(n_421)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_401),
.B(n_406),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_317),
.Y(n_402)
);

INVx5_ASAP7_75t_SL g403 ( 
.A(n_346),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_359),
.Y(n_404)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_404),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_345),
.C(n_342),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_SL g407 ( 
.A(n_370),
.B(n_330),
.C(n_325),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_407),
.A2(n_410),
.B(n_412),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_408),
.A2(n_351),
.B1(n_353),
.B2(n_381),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_365),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_409),
.B(n_411),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_358),
.A2(n_341),
.B1(n_364),
.B2(n_357),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_365),
.B(n_324),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_362),
.A2(n_296),
.B(n_297),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_352),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_414),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_352),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_356),
.B(n_296),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_R g427 ( 
.A(n_416),
.B(n_350),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_362),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_417),
.B(n_379),
.Y(n_439)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_361),
.Y(n_418)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_418),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_R g479 ( 
.A(n_420),
.B(n_427),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_421),
.A2(n_394),
.B1(n_398),
.B2(n_419),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_340),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_444),
.C(n_415),
.Y(n_457)
);

OAI22x1_ASAP7_75t_L g475 ( 
.A1(n_425),
.A2(n_354),
.B1(n_368),
.B2(n_337),
.Y(n_475)
);

AO21x1_ASAP7_75t_L g428 ( 
.A1(n_417),
.A2(n_370),
.B(n_369),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_428),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_431),
.B(n_415),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_381),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_432),
.B(n_445),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_384),
.A2(n_371),
.B(n_357),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_452),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_437),
.A2(n_379),
.B1(n_350),
.B2(n_377),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_353),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_438),
.Y(n_480)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_439),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_412),
.A2(n_346),
.B(n_350),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_385),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_409),
.B(n_348),
.Y(n_443)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_443),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_405),
.B(n_338),
.C(n_361),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_393),
.B(n_354),
.Y(n_445)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_397),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_453),
.B(n_457),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_451),
.A2(n_408),
.B1(n_396),
.B2(n_410),
.Y(n_454)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_454),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_SL g456 ( 
.A(n_451),
.B(n_387),
.C(n_416),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_456),
.B(n_458),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_SL g458 ( 
.A(n_425),
.B(n_416),
.C(n_407),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_460),
.A2(n_433),
.B(n_450),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_435),
.A2(n_394),
.B1(n_414),
.B2(n_413),
.Y(n_461)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_461),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_431),
.B(n_399),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_476),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_463),
.A2(n_429),
.B1(n_427),
.B2(n_438),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_444),
.B(n_419),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_466),
.C(n_468),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_422),
.B(n_398),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_435),
.B(n_395),
.Y(n_467)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_467),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_421),
.B(n_400),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_424),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_469),
.B(n_473),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_441),
.A2(n_403),
.B1(n_418),
.B2(n_404),
.Y(n_470)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_470),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_442),
.Y(n_472)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_472),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_314),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_474),
.A2(n_477),
.B1(n_438),
.B2(n_429),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_475),
.B(n_481),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_447),
.A2(n_376),
.B1(n_374),
.B2(n_390),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_425),
.B(n_443),
.C(n_420),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_478),
.B(n_453),
.C(n_462),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_441),
.B(n_424),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_485),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_486),
.B(n_492),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_457),
.B(n_423),
.C(n_437),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_487),
.B(n_488),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_423),
.C(n_440),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_480),
.B(n_426),
.Y(n_489)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_489),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_428),
.C(n_426),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_491),
.B(n_498),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_459),
.B(n_446),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_493),
.B(n_504),
.Y(n_519)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_494),
.Y(n_515)
);

NOR2x1_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_439),
.Y(n_497)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_497),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_468),
.B(n_428),
.C(n_446),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_447),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_499),
.B(n_452),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_500),
.A2(n_449),
.B1(n_448),
.B2(n_434),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_455),
.B(n_390),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_485),
.A2(n_471),
.B(n_479),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g535 ( 
.A1(n_506),
.A2(n_501),
.B(n_495),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_502),
.A2(n_479),
.B(n_474),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_509),
.B(n_512),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_483),
.B(n_463),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_510),
.B(n_524),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_483),
.B(n_475),
.C(n_430),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_511),
.B(n_520),
.Y(n_528)
);

BUFx12f_ASAP7_75t_SL g512 ( 
.A(n_488),
.Y(n_512)
);

OAI21xp33_ASAP7_75t_L g513 ( 
.A1(n_503),
.A2(n_448),
.B(n_430),
.Y(n_513)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_513),
.Y(n_526)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_518),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_477),
.Y(n_520)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_522),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_490),
.B(n_449),
.C(n_436),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_523),
.B(n_498),
.C(n_499),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_491),
.B(n_434),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_497),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_517),
.A2(n_496),
.B1(n_502),
.B2(n_505),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_525),
.A2(n_527),
.B1(n_269),
.B2(n_278),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_515),
.A2(n_484),
.B1(n_500),
.B2(n_489),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_529),
.B(n_530),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_523),
.B(n_490),
.C(n_486),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_532),
.B(n_534),
.Y(n_543)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_522),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_535),
.A2(n_507),
.B(n_521),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_520),
.B(n_494),
.C(n_482),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_537),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_516),
.B(n_482),
.C(n_472),
.Y(n_537)
);

FAx1_ASAP7_75t_SL g538 ( 
.A(n_506),
.B(n_442),
.CI(n_298),
.CON(n_538),
.SN(n_538)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_538),
.B(n_513),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_SL g549 ( 
.A(n_539),
.B(n_514),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_541),
.A2(n_545),
.B(n_546),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_531),
.A2(n_521),
.B1(n_519),
.B2(n_511),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_544),
.B(n_536),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_540),
.A2(n_508),
.B(n_512),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_540),
.A2(n_514),
.B(n_510),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_537),
.B(n_526),
.Y(n_547)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_547),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_549),
.B(n_552),
.C(n_535),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_550),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_551),
.B(n_538),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_529),
.A2(n_258),
.B(n_306),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_554),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_543),
.B(n_532),
.C(n_528),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_556),
.Y(n_562)
);

AOI31xp67_ASAP7_75t_L g558 ( 
.A1(n_542),
.A2(n_525),
.A3(n_538),
.B(n_527),
.Y(n_558)
);

AOI322xp5_ASAP7_75t_L g561 ( 
.A1(n_558),
.A2(n_547),
.A3(n_533),
.B1(n_550),
.B2(n_551),
.C1(n_548),
.C2(n_539),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_560),
.B(n_258),
.Y(n_563)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_561),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_563),
.B(n_559),
.C(n_557),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_565),
.B(n_272),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_564),
.B(n_560),
.C(n_555),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_566),
.B(n_562),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_568),
.B(n_569),
.C(n_567),
.Y(n_570)
);

AOI322xp5_ASAP7_75t_L g571 ( 
.A1(n_570),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_571),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_572)
);

BUFx24_ASAP7_75t_SL g573 ( 
.A(n_572),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_573),
.A2(n_7),
.B1(n_10),
.B2(n_567),
.Y(n_574)
);


endmodule