module fake_jpeg_11990_n_464 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_464);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_464;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_46),
.Y(n_154)
);

HAxp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_0),
.CON(n_47),
.SN(n_47)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_47),
.B(n_62),
.Y(n_123)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_49),
.Y(n_155)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_50),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_51),
.Y(n_139)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_52),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_56),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_59),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_11),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx2_ASAP7_75t_SL g121 ( 
.A(n_71),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_16),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_93),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_24),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_80),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_0),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_95),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_35),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_96),
.B(n_98),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_17),
.B(n_1),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_99),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_17),
.B(n_3),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_49),
.A2(n_41),
.B1(n_35),
.B2(n_25),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_122),
.A2(n_148),
.B1(n_26),
.B2(n_14),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_41),
.B1(n_20),
.B2(n_34),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_144),
.B1(n_22),
.B2(n_39),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_84),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_135),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_84),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_62),
.B(n_20),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_149),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_80),
.A2(n_41),
.B1(n_34),
.B2(n_25),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_47),
.A2(n_19),
.B1(n_95),
.B2(n_94),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_42),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_83),
.B(n_39),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_23),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_154),
.Y(n_157)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_110),
.B(n_96),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_166),
.C(n_192),
.Y(n_221)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_133),
.A2(n_19),
.B1(n_18),
.B2(n_38),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_162),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_208)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

BUFx4f_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_164),
.Y(n_227)
);

BUFx12_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_165),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_38),
.C(n_18),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_148),
.B1(n_87),
.B2(n_76),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_200),
.B1(n_103),
.B2(n_68),
.Y(n_209)
);

INVx4_ASAP7_75t_SL g169 ( 
.A(n_127),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_169),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_66),
.B1(n_57),
.B2(n_54),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_185),
.B1(n_193),
.B2(n_67),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_28),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_180),
.Y(n_215)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_131),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_178),
.Y(n_202)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_175),
.Y(n_229)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_176),
.Y(n_231)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_119),
.B1(n_155),
.B2(n_115),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_108),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_107),
.B(n_28),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_127),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_183),
.Y(n_211)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_133),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_117),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_190),
.C(n_197),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_132),
.A2(n_88),
.B1(n_82),
.B2(n_74),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_189),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_124),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_100),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_22),
.B(n_14),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_145),
.A2(n_73),
.B1(n_70),
.B2(n_69),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_103),
.A2(n_19),
.B1(n_26),
.B2(n_13),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_198),
.Y(n_219)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_137),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_113),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_113),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_105),
.B1(n_115),
.B2(n_138),
.Y(n_201)
);

AO21x2_ASAP7_75t_L g240 ( 
.A1(n_201),
.A2(n_230),
.B(n_163),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_102),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_204),
.B(n_216),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_199),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_209),
.A2(n_223),
.B1(n_161),
.B2(n_141),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_159),
.B(n_104),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_220),
.B1(n_228),
.B2(n_199),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_174),
.A2(n_140),
.B1(n_119),
.B2(n_139),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_168),
.A2(n_140),
.B1(n_139),
.B2(n_150),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_177),
.A2(n_166),
.B1(n_172),
.B2(n_178),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_150),
.B1(n_134),
.B2(n_155),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_171),
.B(n_106),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_232),
.B(n_118),
.Y(n_250)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_244),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_180),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_236),
.B(n_246),
.Y(n_261)
);

AO21x1_ASAP7_75t_L g281 ( 
.A1(n_237),
.A2(n_205),
.B(n_224),
.Y(n_281)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_238),
.Y(n_272)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_239),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_243),
.B1(n_247),
.B2(n_251),
.Y(n_266)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_242),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_204),
.A2(n_198),
.B1(n_195),
.B2(n_51),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_203),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_226),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_254),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_167),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_212),
.A2(n_179),
.B1(n_176),
.B2(n_188),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_157),
.B(n_191),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_248),
.A2(n_255),
.B(n_208),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_250),
.B(n_222),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_187),
.B1(n_158),
.B2(n_160),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_196),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_259),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_221),
.A2(n_142),
.B(n_126),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_209),
.A2(n_100),
.B(n_154),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_257),
.B1(n_218),
.B2(n_207),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_109),
.B1(n_129),
.B2(n_141),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_260),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_175),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_217),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_238),
.B(n_215),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_263),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_265),
.A2(n_273),
.B1(n_240),
.B2(n_206),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_239),
.B(n_215),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_275),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_280),
.B(n_275),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_220),
.B1(n_205),
.B2(n_207),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_246),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_276),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_205),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_247),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_206),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_235),
.B(n_258),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_282),
.Y(n_299)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_222),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_284),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_213),
.C(n_210),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_251),
.Y(n_285)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_259),
.B(n_210),
.Y(n_286)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

OAI22x1_ASAP7_75t_SL g288 ( 
.A1(n_280),
.A2(n_241),
.B1(n_240),
.B2(n_237),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_288),
.A2(n_290),
.B1(n_300),
.B2(n_301),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_255),
.B1(n_252),
.B2(n_240),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_SL g325 ( 
.A1(n_292),
.A2(n_283),
.B(n_282),
.C(n_269),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_253),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_293),
.A2(n_295),
.B(n_262),
.C(n_302),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_248),
.B(n_250),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_294),
.A2(n_309),
.B(n_264),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_266),
.A2(n_240),
.B1(n_257),
.B2(n_245),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_296),
.A2(n_298),
.B1(n_265),
.B2(n_285),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_243),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_283),
.C(n_286),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_266),
.A2(n_240),
.B1(n_243),
.B2(n_260),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_281),
.A2(n_240),
.B1(n_260),
.B2(n_254),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_270),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_311),
.Y(n_324)
);

OAI22x1_ASAP7_75t_SL g306 ( 
.A1(n_273),
.A2(n_244),
.B1(n_242),
.B2(n_225),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_306),
.A2(n_276),
.B1(n_277),
.B2(n_272),
.Y(n_322)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_271),
.A2(n_225),
.B(n_229),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_310),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_279),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_267),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_274),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_309),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_327),
.Y(n_354)
);

AO21x1_ASAP7_75t_L g353 ( 
.A1(n_315),
.A2(n_325),
.B(n_229),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_316),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_292),
.A2(n_269),
.B(n_267),
.Y(n_317)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_317),
.B(n_333),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_319),
.A2(n_290),
.B1(n_300),
.B2(n_288),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_289),
.A2(n_272),
.B1(n_277),
.B2(n_284),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_320),
.A2(n_189),
.B1(n_152),
.B2(n_129),
.Y(n_363)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_321),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_322),
.A2(n_326),
.B1(n_303),
.B2(n_312),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_323),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_296),
.A2(n_261),
.B1(n_278),
.B2(n_263),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_313),
.Y(n_327)
);

NAND3xp33_ASAP7_75t_L g328 ( 
.A(n_295),
.B(n_268),
.C(n_262),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_335),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_284),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_332),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_289),
.A2(n_287),
.B(n_227),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_305),
.B(n_299),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_334),
.B(n_336),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_291),
.B(n_169),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_293),
.B(n_165),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g337 ( 
.A(n_294),
.B(n_165),
.CI(n_214),
.CON(n_337),
.SN(n_337)
);

FAx1_ASAP7_75t_SL g358 ( 
.A(n_337),
.B(n_214),
.CI(n_37),
.CON(n_358),
.SN(n_358)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_299),
.B(n_146),
.Y(n_338)
);

XOR2x2_ASAP7_75t_L g342 ( 
.A(n_338),
.B(n_336),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_304),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_231),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_297),
.C(n_291),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_340),
.B(n_350),
.C(n_352),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_342),
.B(n_349),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_318),
.A2(n_298),
.B1(n_303),
.B2(n_311),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_343),
.A2(n_345),
.B1(n_363),
.B2(n_331),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_344),
.A2(n_361),
.B1(n_189),
.B2(n_214),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_318),
.A2(n_322),
.B1(n_330),
.B2(n_324),
.Y(n_348)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_348),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_SL g349 ( 
.A(n_320),
.B(n_307),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_307),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_310),
.C(n_306),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_353),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_330),
.A2(n_254),
.B1(n_227),
.B2(n_231),
.Y(n_355)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_355),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_358),
.A2(n_14),
.B(n_13),
.Y(n_382)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_360),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_314),
.A2(n_189),
.B1(n_186),
.B2(n_182),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_164),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_346),
.C(n_325),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_SL g364 ( 
.A(n_359),
.B(n_324),
.C(n_315),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_341),
.Y(n_397)
);

FAx1_ASAP7_75t_SL g368 ( 
.A(n_351),
.B(n_316),
.CI(n_325),
.CON(n_368),
.SN(n_368)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_342),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_353),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_372),
.A2(n_374),
.B1(n_382),
.B2(n_3),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_340),
.B(n_325),
.C(n_317),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_381),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_343),
.A2(n_331),
.B1(n_333),
.B2(n_337),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_347),
.A2(n_337),
.B1(n_152),
.B2(n_64),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_375),
.A2(n_377),
.B1(n_378),
.B2(n_341),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_344),
.A2(n_60),
.B1(n_53),
.B2(n_63),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_354),
.Y(n_379)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_357),
.Y(n_380)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_380),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_346),
.B(n_13),
.C(n_26),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_350),
.C(n_356),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_384),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_23),
.C(n_37),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_341),
.C(n_349),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_SL g407 ( 
.A(n_385),
.B(n_389),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_387),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_362),
.Y(n_388)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_388),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_390),
.A2(n_369),
.B1(n_374),
.B2(n_382),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_361),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_393),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_341),
.C(n_358),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_398),
.C(n_399),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_376),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_372),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_369),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_402),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_358),
.C(n_37),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_376),
.B(n_3),
.C(n_4),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_401),
.Y(n_415)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_367),
.Y(n_403)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_403),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_408),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_406),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_384),
.C(n_381),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_368),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_411),
.A2(n_392),
.B(n_399),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_368),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_412),
.B(n_413),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_395),
.A2(n_377),
.B1(n_378),
.B2(n_24),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_3),
.C(n_4),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_414),
.B(n_416),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_4),
.C(n_5),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_411),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_420),
.B(n_423),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_385),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_424),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_389),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_400),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_425),
.B(n_427),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_401),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_404),
.B(n_398),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_428),
.B(n_431),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_24),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_407),
.B(n_24),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_414),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_419),
.A2(n_24),
.B1(n_44),
.B2(n_6),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_433),
.B(n_405),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_426),
.A2(n_419),
.B(n_415),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_SL g445 ( 
.A(n_434),
.B(n_439),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_410),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_436),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_418),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_437),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_421),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_440),
.B(n_444),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_441),
.B(n_432),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_SL g444 ( 
.A(n_423),
.B(n_416),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_445),
.A2(n_4),
.B(n_5),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_446),
.B(n_447),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_429),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_413),
.Y(n_450)
);

OAI21x1_ASAP7_75t_SL g452 ( 
.A1(n_450),
.A2(n_438),
.B(n_44),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_452),
.A2(n_454),
.B(n_455),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_449),
.A2(n_438),
.B(n_5),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_449),
.A2(n_4),
.B(n_5),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_456),
.Y(n_458)
);

AOI321xp33_ASAP7_75t_L g457 ( 
.A1(n_453),
.A2(n_451),
.A3(n_448),
.B1(n_8),
.B2(n_9),
.C(n_7),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_457),
.A2(n_6),
.B(n_7),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_460),
.A2(n_461),
.B(n_7),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_459),
.B(n_458),
.C(n_8),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_462),
.A2(n_7),
.B(n_8),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_463),
.A2(n_9),
.B(n_437),
.Y(n_464)
);


endmodule