module fake_netlist_1_12378_n_31 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_31);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g13 ( .A(n_11), .B(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
BUFx6f_ASAP7_75t_SL g19 ( .A(n_18), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_15), .B(n_0), .Y(n_20) );
AOI22xp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_14), .B1(n_17), .B2(n_13), .Y(n_21) );
AOI221xp5_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_13), .B1(n_16), .B2(n_3), .C(n_5), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_19), .B1(n_2), .B2(n_3), .Y(n_23) );
OAI21xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_22), .B(n_19), .Y(n_24) );
HAxp5_ASAP7_75t_SL g25 ( .A(n_24), .B(n_1), .CON(n_25), .SN(n_25) );
AOI221xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_2), .B1(n_5), .B2(n_6), .C(n_7), .Y(n_26) );
INVxp67_ASAP7_75t_SL g27 ( .A(n_25), .Y(n_27) );
BUFx2_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_26), .B(n_25), .Y(n_29) );
INVx1_ASAP7_75t_SL g30 ( .A(n_28), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_29), .B1(n_8), .B2(n_9), .Y(n_31) );
endmodule