module fake_jpeg_18013_n_375 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_375);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_375;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_11),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx2_ASAP7_75t_SL g100 ( 
.A(n_39),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g114 ( 
.A(n_41),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_50),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_6),
.B(n_12),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_52),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_6),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_60),
.Y(n_101)
);

HAxp5_ASAP7_75t_SL g60 ( 
.A(n_20),
.B(n_7),
.CON(n_60),
.SN(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_63),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_7),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_7),
.C(n_12),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_74)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_29),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_68),
.B1(n_19),
.B2(n_28),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_29),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_16),
.B1(n_18),
.B2(n_34),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_70),
.A2(n_72),
.B1(n_77),
.B2(n_80),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_18),
.B1(n_34),
.B2(n_57),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_10),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_18),
.B1(n_20),
.B2(n_31),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_31),
.B1(n_14),
.B2(n_30),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_78),
.A2(n_79),
.B1(n_86),
.B2(n_97),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_59),
.B1(n_65),
.B2(n_62),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_14),
.B1(n_33),
.B2(n_32),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_14),
.B1(n_33),
.B2(n_32),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_81),
.A2(n_85),
.B1(n_90),
.B2(n_96),
.Y(n_126)
);

BUFx2_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g147 ( 
.A(n_82),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_36),
.B1(n_30),
.B2(n_35),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_36),
.B1(n_19),
.B2(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_21),
.B1(n_35),
.B2(n_7),
.Y(n_90)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_19),
.B1(n_26),
.B2(n_35),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_95),
.B1(n_103),
.B2(n_109),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_61),
.B1(n_52),
.B2(n_53),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_21),
.B1(n_5),
.B2(n_8),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_40),
.A2(n_68),
.B1(n_67),
.B2(n_64),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_38),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_8),
.B1(n_9),
.B2(n_13),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_108),
.B1(n_110),
.B2(n_0),
.Y(n_136)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_107),
.B(n_75),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_47),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_41),
.A2(n_37),
.B1(n_28),
.B2(n_9),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_50),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_51),
.A2(n_4),
.B1(n_10),
.B2(n_5),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_112),
.A2(n_115),
.B1(n_3),
.B2(n_109),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_56),
.A2(n_4),
.B1(n_10),
.B2(n_37),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_28),
.Y(n_149)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_53),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_123),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_45),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_43),
.C(n_42),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_124),
.B(n_159),
.Y(n_170)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_76),
.B(n_37),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_128),
.B(n_144),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_130),
.A2(n_133),
.B1(n_132),
.B2(n_131),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_131),
.B(n_141),
.Y(n_194)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_92),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_136),
.A2(n_164),
.B1(n_165),
.B2(n_147),
.Y(n_201)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_76),
.A2(n_28),
.B1(n_37),
.B2(n_39),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_146),
.B(n_151),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_74),
.A2(n_37),
.B(n_1),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_142),
.A2(n_156),
.B(n_114),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_58),
.B(n_28),
.C(n_2),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_143),
.A2(n_148),
.B(n_100),
.C(n_114),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_0),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_101),
.A2(n_28),
.B1(n_58),
.B2(n_2),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_69),
.A2(n_84),
.B(n_89),
.C(n_83),
.Y(n_148)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_89),
.B(n_58),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_150),
.B(n_152),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_69),
.A2(n_58),
.B(n_1),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_84),
.B(n_0),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_95),
.B(n_3),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_154),
.B(n_86),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_155),
.A2(n_164),
.B1(n_161),
.B2(n_121),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_112),
.A2(n_103),
.B(n_94),
.C(n_116),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_162),
.Y(n_197)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_113),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_137),
.Y(n_208)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_106),
.B(n_107),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_75),
.B(n_107),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_102),
.A2(n_99),
.B1(n_71),
.B2(n_118),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_75),
.B(n_91),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_166),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_99),
.A2(n_117),
.B1(n_93),
.B2(n_92),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_167),
.A2(n_114),
.B1(n_125),
.B2(n_132),
.Y(n_188)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_169),
.Y(n_206)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_100),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_180),
.B(n_209),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_120),
.A2(n_92),
.B1(n_102),
.B2(n_114),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_193),
.B1(n_199),
.B2(n_202),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_191),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_186),
.A2(n_195),
.B(n_212),
.Y(n_216)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_123),
.A2(n_114),
.B(n_128),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_187),
.A2(n_182),
.B(n_200),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_188),
.A2(n_203),
.B1(n_205),
.B2(n_183),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_142),
.A2(n_144),
.B(n_145),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_119),
.B(n_129),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_191),
.A2(n_201),
.B1(n_207),
.B2(n_211),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_126),
.A2(n_156),
.B1(n_124),
.B2(n_138),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_130),
.B(n_151),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_208),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_156),
.A2(n_140),
.B1(n_146),
.B2(n_130),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_196),
.A2(n_171),
.B1(n_211),
.B2(n_175),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_143),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_156),
.A2(n_160),
.B1(n_153),
.B2(n_127),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_159),
.B1(n_135),
.B2(n_134),
.Y(n_202)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_147),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_210),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_134),
.A2(n_135),
.B1(n_133),
.B2(n_158),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_133),
.B(n_168),
.Y(n_209)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_133),
.B(n_157),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_139),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_216),
.A2(n_220),
.B(n_229),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_217),
.B(n_223),
.Y(n_276)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_225),
.B(n_215),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_186),
.A2(n_170),
.B(n_209),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_227),
.B(n_228),
.Y(n_277)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_230),
.A2(n_240),
.B1(n_215),
.B2(n_235),
.Y(n_269)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_175),
.B(n_170),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_178),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_193),
.A2(n_199),
.B1(n_202),
.B2(n_176),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_235),
.B1(n_238),
.B2(n_242),
.Y(n_254)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_171),
.A2(n_188),
.B1(n_196),
.B2(n_207),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_192),
.B(n_190),
.C(n_206),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_236),
.B(n_246),
.C(n_245),
.Y(n_283)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_198),
.A2(n_192),
.B1(n_180),
.B2(n_185),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_181),
.A2(n_182),
.B1(n_190),
.B2(n_206),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_243),
.A2(n_252),
.B(n_174),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_244),
.A2(n_245),
.B1(n_225),
.B2(n_247),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_203),
.A2(n_214),
.B1(n_197),
.B2(n_179),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_194),
.B(n_172),
.C(n_205),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_184),
.Y(n_247)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_247),
.Y(n_281)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_249),
.Y(n_259)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_183),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_250),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_172),
.A2(n_183),
.B(n_178),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_263),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_255),
.B(n_256),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_210),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_258),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_178),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_174),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_264),
.A2(n_266),
.B(n_272),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_237),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_265),
.B(n_255),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_229),
.A2(n_174),
.B(n_251),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_246),
.B1(n_252),
.B2(n_239),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_222),
.B(n_221),
.Y(n_271)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_219),
.A2(n_220),
.B1(n_242),
.B2(n_230),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_266),
.Y(n_299)
);

A2O1A1O1Ixp25_ASAP7_75t_L g279 ( 
.A1(n_216),
.A2(n_238),
.B(n_219),
.C(n_218),
.D(n_233),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_283),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_243),
.A2(n_221),
.B(n_218),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_261),
.B(n_278),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_248),
.B1(n_249),
.B2(n_217),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_223),
.A2(n_227),
.B1(n_228),
.B2(n_218),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_258),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_260),
.B(n_236),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_293),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_288),
.A2(n_282),
.B1(n_262),
.B2(n_267),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_241),
.Y(n_289)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_289),
.Y(n_318)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_299),
.B1(n_309),
.B2(n_269),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_260),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_263),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_297),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_257),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_301),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_259),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_264),
.B(n_261),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_302),
.A2(n_304),
.B(n_305),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_276),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_303),
.A2(n_306),
.B1(n_281),
.B2(n_270),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_280),
.B(n_278),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_268),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_254),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_262),
.C(n_256),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_272),
.C(n_259),
.Y(n_308)
);

NOR3xp33_ASAP7_75t_SL g328 ( 
.A(n_308),
.B(n_296),
.C(n_286),
.Y(n_328)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_268),
.Y(n_309)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_274),
.A2(n_284),
.B(n_267),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_310),
.A2(n_275),
.B1(n_281),
.B2(n_306),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_323),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_254),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_312),
.B(n_314),
.C(n_320),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_313),
.A2(n_315),
.B1(n_316),
.B2(n_321),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_282),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_298),
.A2(n_293),
.B1(n_287),
.B2(n_292),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_298),
.A2(n_287),
.B1(n_289),
.B2(n_305),
.Y(n_316)
);

AOI22x1_ASAP7_75t_L g321 ( 
.A1(n_291),
.A2(n_277),
.B1(n_275),
.B2(n_270),
.Y(n_321)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_322),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_296),
.A2(n_304),
.B1(n_302),
.B2(n_294),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_324),
.A2(n_329),
.B1(n_330),
.B2(n_321),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_328),
.B(n_303),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_300),
.A2(n_309),
.B1(n_290),
.B2(n_307),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_290),
.A2(n_282),
.B1(n_288),
.B2(n_299),
.Y(n_330)
);

OAI32xp33_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_303),
.A3(n_326),
.B1(n_321),
.B2(n_318),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_332),
.B(n_335),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_327),
.B(n_317),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_333),
.B(n_343),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_329),
.C(n_314),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_337),
.B(n_339),
.C(n_336),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_312),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_315),
.Y(n_340)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_340),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_326),
.Y(n_341)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_341),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_325),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_342),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_318),
.Y(n_343)
);

NAND2x1_ASAP7_75t_SL g345 ( 
.A(n_319),
.B(n_323),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_344),
.A2(n_313),
.B1(n_319),
.B2(n_328),
.Y(n_346)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_346),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_350),
.C(n_355),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_336),
.C(n_339),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_331),
.Y(n_352)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_352),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_334),
.C(n_338),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_334),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_356),
.B(n_359),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_348),
.A2(n_331),
.B(n_345),
.Y(n_358)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_358),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_338),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_352),
.A2(n_353),
.B(n_355),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_362),
.A2(n_351),
.B(n_347),
.Y(n_364)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_364),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_360),
.B(n_354),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_366),
.B(n_362),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_363),
.B(n_356),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_367),
.B(n_368),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_365),
.Y(n_371)
);

AOI21x1_ASAP7_75t_L g372 ( 
.A1(n_371),
.A2(n_359),
.B(n_353),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_346),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_370),
.B(n_357),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_361),
.Y(n_375)
);


endmodule