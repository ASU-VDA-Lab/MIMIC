module fake_netlist_6_1055_n_1361 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_341, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_350, n_78, n_84, n_142, n_143, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_353, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_348, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1361);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_341;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1361;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_595;
wire n_627;
wire n_524;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_1339;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_312),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_350),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_354),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_16),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_127),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_145),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_188),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_216),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_153),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_102),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_175),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_162),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_220),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_141),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_116),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_325),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_208),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_225),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_26),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_44),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_88),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_337),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_192),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_9),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_255),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_55),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_273),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_300),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_244),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_151),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_194),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_146),
.B(n_68),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_206),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_72),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_306),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_253),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_128),
.B(n_310),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_321),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_143),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_15),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_355),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_259),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_169),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_251),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_56),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_357),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_129),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_101),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_295),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_241),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_156),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_254),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_66),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_120),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_237),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_261),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_21),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_103),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_289),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_327),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_316),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_223),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_270),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_187),
.Y(n_424)
);

INVxp33_ASAP7_75t_SL g425 ( 
.A(n_274),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_200),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_214),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_122),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_150),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_28),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_213),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_330),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_328),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_101),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_313),
.Y(n_435)
);

BUFx10_ASAP7_75t_L g436 ( 
.A(n_191),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_222),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_120),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_185),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_263),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_89),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_299),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_335),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_93),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_155),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_163),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_344),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_320),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_15),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_256),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_301),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_36),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_249),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_236),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_277),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_116),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_154),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_288),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_82),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_278),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_358),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_158),
.B(n_103),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_34),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_28),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_4),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_331),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_30),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_83),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_250),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_215),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_33),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_196),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_L g473 ( 
.A(n_233),
.B(n_189),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_56),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_55),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_69),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_343),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_359),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_179),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_314),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_180),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_198),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_235),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_102),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_135),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_304),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_78),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_130),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_182),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_164),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_37),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_49),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_266),
.B(n_58),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_177),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_134),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_67),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_81),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_230),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_49),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_157),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_193),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_190),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_342),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_12),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_257),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_39),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_272),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_34),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_293),
.Y(n_509)
);

CKINVDCx14_ASAP7_75t_R g510 ( 
.A(n_160),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_115),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_292),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_323),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_23),
.Y(n_514)
);

INVxp33_ASAP7_75t_L g515 ( 
.A(n_176),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_58),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_248),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_205),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_152),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_186),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_227),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_159),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_207),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_76),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_67),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_61),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_147),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_115),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_276),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_229),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_51),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_352),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_113),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_356),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_29),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_226),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_307),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_100),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_329),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_231),
.Y(n_540)
);

OAI22x1_ASAP7_75t_SL g541 ( 
.A1(n_430),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_541)
);

OA22x2_ASAP7_75t_L g542 ( 
.A1(n_384),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_431),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_438),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_456),
.Y(n_545)
);

INVx6_ASAP7_75t_L g546 ( 
.A(n_436),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_438),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_492),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_456),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_447),
.B(n_3),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_456),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_481),
.B(n_3),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_431),
.Y(n_553)
);

OA21x2_ASAP7_75t_L g554 ( 
.A1(n_444),
.A2(n_4),
.B(n_5),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_475),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_431),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_475),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_481),
.B(n_5),
.Y(n_558)
);

CKINVDCx11_ASAP7_75t_R g559 ( 
.A(n_491),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_502),
.B(n_362),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_384),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_431),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_475),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_469),
.B(n_6),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_533),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_469),
.B(n_6),
.Y(n_566)
);

BUFx8_ASAP7_75t_L g567 ( 
.A(n_412),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_533),
.Y(n_568)
);

OA21x2_ASAP7_75t_L g569 ( 
.A1(n_444),
.A2(n_7),
.B(n_8),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_515),
.B(n_7),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_SL g571 ( 
.A1(n_506),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_533),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_378),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_502),
.B(n_10),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_379),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_470),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_416),
.B(n_521),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_470),
.B(n_11),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_499),
.B(n_11),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_380),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_368),
.A2(n_137),
.B(n_136),
.Y(n_581)
);

OAI21x1_ASAP7_75t_L g582 ( 
.A1(n_368),
.A2(n_139),
.B(n_138),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_526),
.Y(n_583)
);

CKINVDCx16_ASAP7_75t_R g584 ( 
.A(n_385),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_386),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_394),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_375),
.B(n_12),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_363),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_405),
.Y(n_589)
);

BUFx12f_ASAP7_75t_L g590 ( 
.A(n_436),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_499),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_364),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_408),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_433),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_433),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_369),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_433),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_399),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_598)
);

AOI22x1_ASAP7_75t_SL g599 ( 
.A1(n_511),
.A2(n_18),
.B1(n_14),
.B2(n_17),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_413),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_415),
.B(n_17),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_414),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_418),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_428),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_409),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_441),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_449),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_459),
.Y(n_608)
);

OA21x2_ASAP7_75t_L g609 ( 
.A1(n_465),
.A2(n_19),
.B(n_20),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_374),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_534),
.B(n_22),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_381),
.A2(n_142),
.B(n_140),
.Y(n_612)
);

OA21x2_ASAP7_75t_L g613 ( 
.A1(n_474),
.A2(n_22),
.B(n_23),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_487),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_534),
.Y(n_615)
);

CKINVDCx11_ASAP7_75t_R g616 ( 
.A(n_538),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_488),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_401),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_401),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_545),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_545),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_565),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_568),
.Y(n_623)
);

NAND3xp33_ASAP7_75t_L g624 ( 
.A(n_577),
.B(n_560),
.C(n_570),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_572),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_565),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_549),
.Y(n_627)
);

BUFx10_ASAP7_75t_L g628 ( 
.A(n_577),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_549),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_SL g630 ( 
.A(n_579),
.B(n_493),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_551),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_546),
.B(n_425),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_551),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_543),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_555),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_555),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_584),
.B(n_393),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_596),
.B(n_424),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_610),
.B(n_510),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_576),
.B(n_478),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_618),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_559),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_557),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_546),
.B(n_482),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_588),
.B(n_397),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_576),
.B(n_432),
.Y(n_646)
);

INVxp33_ASAP7_75t_L g647 ( 
.A(n_561),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_615),
.B(n_508),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_542),
.B(n_392),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_L g650 ( 
.A(n_552),
.B(n_462),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_563),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_L g652 ( 
.A(n_558),
.B(n_400),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_563),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_618),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_615),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_618),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_592),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_618),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_L g659 ( 
.A1(n_542),
.A2(n_467),
.B1(n_476),
.B2(n_464),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_619),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_583),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_583),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_619),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_570),
.B(n_389),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_619),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_573),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_666),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_SL g668 ( 
.A1(n_647),
.A2(n_574),
.B1(n_605),
.B2(n_598),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_658),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_634),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_656),
.Y(n_671)
);

NOR3xp33_ASAP7_75t_L g672 ( 
.A(n_624),
.B(n_571),
.C(n_601),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_634),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_649),
.A2(n_564),
.B1(n_566),
.B2(n_550),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_623),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_625),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_638),
.B(n_546),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_622),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_626),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_640),
.B(n_591),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_657),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_649),
.A2(n_564),
.B1(n_566),
.B2(n_550),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_649),
.A2(n_611),
.B1(n_578),
.B2(n_609),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_660),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_639),
.B(n_590),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_664),
.B(n_590),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_649),
.A2(n_611),
.B1(n_578),
.B2(n_609),
.Y(n_687)
);

OAI221xp5_ASAP7_75t_L g688 ( 
.A1(n_630),
.A2(n_587),
.B1(n_593),
.B2(n_575),
.C(n_586),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_644),
.B(n_567),
.Y(n_689)
);

BUFx5_ASAP7_75t_L g690 ( 
.A(n_627),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_626),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_620),
.B(n_543),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_620),
.B(n_543),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_650),
.A2(n_372),
.B1(n_402),
.B2(n_360),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_640),
.B(n_561),
.Y(n_695)
);

OR2x6_ASAP7_75t_L g696 ( 
.A(n_655),
.B(n_593),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_632),
.B(n_567),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_665),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_655),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_621),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_648),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_648),
.B(n_544),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_646),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_647),
.B(n_547),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_641),
.B(n_597),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_621),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_637),
.Y(n_707)
);

AO221x1_ASAP7_75t_L g708 ( 
.A1(n_659),
.A2(n_504),
.B1(n_366),
.B2(n_367),
.C(n_365),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_629),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_628),
.B(n_454),
.Y(n_710)
);

OAI221xp5_ASAP7_75t_L g711 ( 
.A1(n_652),
.A2(n_602),
.B1(n_603),
.B2(n_589),
.C(n_580),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_629),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_628),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_652),
.A2(n_613),
.B1(n_609),
.B2(n_569),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_641),
.B(n_562),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_628),
.B(n_477),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_631),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_641),
.B(n_594),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_654),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_645),
.B(n_485),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_633),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_654),
.B(n_530),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_663),
.B(n_543),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_635),
.B(n_553),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_663),
.A2(n_503),
.B1(n_370),
.B2(n_371),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_SL g726 ( 
.A(n_642),
.B(n_417),
.C(n_407),
.Y(n_726)
);

INVxp33_ASAP7_75t_L g727 ( 
.A(n_661),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_661),
.A2(n_434),
.B1(n_463),
.B2(n_452),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_680),
.B(n_548),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_718),
.A2(n_634),
.B(n_653),
.Y(n_730)
);

NAND2x1_ASAP7_75t_L g731 ( 
.A(n_719),
.B(n_634),
.Y(n_731)
);

OAI21xp5_ASAP7_75t_L g732 ( 
.A1(n_683),
.A2(n_582),
.B(n_581),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_672),
.A2(n_612),
.B(n_473),
.C(n_435),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_702),
.Y(n_734)
);

BUFx12f_ASAP7_75t_L g735 ( 
.A(n_696),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_704),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_703),
.B(n_636),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_SL g738 ( 
.A(n_694),
.B(n_642),
.C(n_471),
.Y(n_738)
);

OAI21xp5_ASAP7_75t_L g739 ( 
.A1(n_687),
.A2(n_613),
.B(n_569),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_681),
.B(n_559),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_702),
.Y(n_741)
);

AOI21x1_ASAP7_75t_L g742 ( 
.A1(n_723),
.A2(n_651),
.B(n_643),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_699),
.B(n_701),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_682),
.B(n_377),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_717),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_696),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_688),
.B(n_616),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_695),
.B(n_727),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_686),
.B(n_388),
.Y(n_749)
);

AO21x2_ASAP7_75t_L g750 ( 
.A1(n_722),
.A2(n_373),
.B(n_361),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_705),
.A2(n_556),
.B(n_553),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_678),
.B(n_435),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_679),
.B(n_437),
.Y(n_753)
);

INVx3_ASAP7_75t_SL g754 ( 
.A(n_696),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_691),
.B(n_437),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_670),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_675),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_714),
.A2(n_448),
.B1(n_455),
.B2(n_445),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_685),
.A2(n_676),
.B(n_725),
.C(n_671),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_710),
.B(n_606),
.Y(n_760)
);

OAI321xp33_ASAP7_75t_L g761 ( 
.A1(n_711),
.A2(n_528),
.A3(n_531),
.B1(n_516),
.B2(n_614),
.C(n_383),
.Y(n_761)
);

CKINVDCx10_ASAP7_75t_R g762 ( 
.A(n_668),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_670),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_698),
.Y(n_764)
);

O2A1O1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_728),
.A2(n_600),
.B(n_604),
.C(n_585),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_707),
.B(n_662),
.Y(n_766)
);

O2A1O1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_720),
.A2(n_600),
.B(n_604),
.C(n_585),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_669),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_689),
.B(n_391),
.Y(n_769)
);

NOR3xp33_ASAP7_75t_L g770 ( 
.A(n_716),
.B(n_726),
.C(n_697),
.Y(n_770)
);

INVx11_ASAP7_75t_L g771 ( 
.A(n_708),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_684),
.B(n_468),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_700),
.A2(n_455),
.B1(n_505),
.B2(n_448),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_706),
.A2(n_613),
.B(n_569),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_692),
.A2(n_595),
.B(n_662),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_690),
.B(n_376),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_692),
.A2(n_724),
.B(n_693),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_709),
.B(n_607),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_712),
.A2(n_387),
.B(n_390),
.C(n_382),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_724),
.A2(n_406),
.B(n_395),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_721),
.A2(n_398),
.B1(n_403),
.B2(n_396),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_673),
.A2(n_420),
.B(n_419),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_703),
.B(n_422),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_703),
.B(n_423),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_715),
.A2(n_427),
.B(n_426),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_683),
.A2(n_554),
.B(n_451),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_674),
.A2(n_453),
.B1(n_457),
.B2(n_450),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_672),
.A2(n_461),
.B(n_466),
.C(n_458),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_672),
.B(n_404),
.Y(n_789)
);

OAI21xp33_ASAP7_75t_SL g790 ( 
.A1(n_683),
.A2(n_483),
.B(n_480),
.Y(n_790)
);

NOR2x1_ASAP7_75t_L g791 ( 
.A(n_685),
.B(n_554),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_703),
.B(n_486),
.Y(n_792)
);

AOI33xp33_ASAP7_75t_L g793 ( 
.A1(n_695),
.A2(n_608),
.A3(n_617),
.B1(n_541),
.B2(n_501),
.B3(n_490),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_703),
.B(n_498),
.Y(n_794)
);

AND2x6_ASAP7_75t_L g795 ( 
.A(n_677),
.B(n_500),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_699),
.B(n_507),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_713),
.B(n_410),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_715),
.A2(n_519),
.B(n_518),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_683),
.A2(n_529),
.B(n_527),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_703),
.B(n_532),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_667),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_715),
.A2(n_421),
.B(n_411),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_703),
.B(n_484),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_683),
.A2(n_439),
.B(n_429),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_696),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_672),
.A2(n_442),
.B1(n_443),
.B2(n_440),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_703),
.B(n_446),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_703),
.B(n_460),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_672),
.B(n_472),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_672),
.A2(n_497),
.B1(n_514),
.B2(n_496),
.Y(n_810)
);

CKINVDCx10_ASAP7_75t_R g811 ( 
.A(n_696),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_SL g812 ( 
.A(n_713),
.B(n_479),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_667),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_703),
.B(n_489),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_683),
.A2(n_495),
.B(n_494),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_703),
.B(n_509),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_703),
.B(n_524),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_715),
.A2(n_513),
.B(n_512),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_672),
.B(n_517),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_703),
.B(n_525),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_715),
.A2(n_522),
.B(n_520),
.Y(n_821)
);

NOR2x1_ASAP7_75t_SL g822 ( 
.A(n_758),
.B(n_144),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_745),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_SL g824 ( 
.A1(n_770),
.A2(n_599),
.B(n_535),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_748),
.B(n_786),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_739),
.A2(n_536),
.B(n_523),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_734),
.B(n_537),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_734),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_766),
.B(n_539),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_799),
.B(n_540),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_791),
.A2(n_733),
.B(n_790),
.Y(n_831)
);

BUFx10_ASAP7_75t_L g832 ( 
.A(n_740),
.Y(n_832)
);

AO31x2_ASAP7_75t_L g833 ( 
.A1(n_788),
.A2(n_26),
.A3(n_24),
.B(n_25),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_734),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_803),
.B(n_24),
.C(n_25),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_774),
.A2(n_149),
.B(n_148),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_811),
.Y(n_837)
);

OAI21x1_ASAP7_75t_L g838 ( 
.A1(n_742),
.A2(n_730),
.B(n_731),
.Y(n_838)
);

INVx5_ASAP7_75t_L g839 ( 
.A(n_735),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_817),
.B(n_820),
.Y(n_840)
);

AND3x4_ASAP7_75t_L g841 ( 
.A(n_743),
.B(n_27),
.C(n_29),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_736),
.B(n_27),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_783),
.B(n_784),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_768),
.A2(n_353),
.B(n_161),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_756),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_807),
.B(n_30),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_729),
.Y(n_847)
);

OR2x6_ASAP7_75t_L g848 ( 
.A(n_805),
.B(n_31),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_743),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_754),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_792),
.B(n_31),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_789),
.A2(n_819),
.B(n_809),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_776),
.A2(n_815),
.B(n_804),
.Y(n_853)
);

AO21x1_ASAP7_75t_L g854 ( 
.A1(n_787),
.A2(n_32),
.B(n_33),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_808),
.B(n_165),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_746),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_806),
.A2(n_36),
.B(n_32),
.C(n_35),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_794),
.B(n_35),
.Y(n_858)
);

NOR2xp67_ASAP7_75t_L g859 ( 
.A(n_738),
.B(n_166),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_759),
.A2(n_168),
.B1(n_170),
.B2(n_167),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_760),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_778),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_814),
.A2(n_172),
.B1(n_173),
.B2(n_171),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_800),
.B(n_37),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_756),
.Y(n_865)
);

CKINVDCx11_ASAP7_75t_R g866 ( 
.A(n_811),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_737),
.A2(n_178),
.B(n_174),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_763),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_816),
.B(n_181),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_801),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_757),
.B(n_812),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_813),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_L g873 ( 
.A(n_810),
.B(n_38),
.C(n_40),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_SL g874 ( 
.A1(n_763),
.A2(n_184),
.B(n_183),
.Y(n_874)
);

AOI221x1_ASAP7_75t_L g875 ( 
.A1(n_785),
.A2(n_221),
.B1(n_349),
.B2(n_348),
.C(n_346),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_764),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_796),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_750),
.B(n_41),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_797),
.B(n_41),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_752),
.Y(n_880)
);

AO31x2_ASAP7_75t_L g881 ( 
.A1(n_773),
.A2(n_44),
.A3(n_42),
.B(n_43),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_750),
.B(n_42),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_795),
.B(n_772),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_771),
.Y(n_884)
);

INVx5_ASAP7_75t_L g885 ( 
.A(n_795),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_753),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_755),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_795),
.B(n_43),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_795),
.B(n_45),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_798),
.A2(n_197),
.B(n_195),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_744),
.B(n_199),
.Y(n_891)
);

AOI211x1_ASAP7_75t_L g892 ( 
.A1(n_780),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_747),
.A2(n_202),
.B1(n_203),
.B2(n_201),
.Y(n_893)
);

OAI21x1_ASAP7_75t_L g894 ( 
.A1(n_775),
.A2(n_351),
.B(n_204),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_802),
.A2(n_210),
.B(n_209),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_767),
.Y(n_896)
);

OAI21x1_ASAP7_75t_L g897 ( 
.A1(n_751),
.A2(n_345),
.B(n_212),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_818),
.A2(n_217),
.B(n_211),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_821),
.A2(n_219),
.B(n_218),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_749),
.A2(n_239),
.B1(n_341),
.B2(n_340),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_781),
.B(n_224),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_769),
.Y(n_902)
);

AOI221x1_ASAP7_75t_L g903 ( 
.A1(n_782),
.A2(n_238),
.B1(n_339),
.B2(n_338),
.C(n_336),
.Y(n_903)
);

AO31x2_ASAP7_75t_L g904 ( 
.A1(n_779),
.A2(n_48),
.A3(n_50),
.B(n_51),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_765),
.B(n_793),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_761),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_762),
.A2(n_232),
.B(n_228),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_762),
.B(n_48),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_748),
.B(n_50),
.Y(n_909)
);

AO31x2_ASAP7_75t_L g910 ( 
.A1(n_733),
.A2(n_52),
.A3(n_53),
.B(n_54),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_748),
.B(n_57),
.Y(n_911)
);

AOI221x1_ASAP7_75t_L g912 ( 
.A1(n_788),
.A2(n_245),
.B1(n_334),
.B2(n_333),
.C(n_332),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_748),
.B(n_59),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_739),
.A2(n_240),
.B(n_234),
.Y(n_914)
);

BUFx8_ASAP7_75t_L g915 ( 
.A(n_805),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_799),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_741),
.B(n_242),
.Y(n_917)
);

INVx4_ASAP7_75t_L g918 ( 
.A(n_734),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_778),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_748),
.B(n_60),
.Y(n_920)
);

BUFx4_ASAP7_75t_SL g921 ( 
.A(n_805),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_739),
.A2(n_246),
.B(n_243),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_811),
.Y(n_923)
);

OAI21x1_ASAP7_75t_SL g924 ( 
.A1(n_799),
.A2(n_252),
.B(n_247),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_811),
.Y(n_925)
);

AOI211x1_ASAP7_75t_L g926 ( 
.A1(n_799),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_778),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_778),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_739),
.A2(n_260),
.B(n_258),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_741),
.B(n_262),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_734),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_741),
.B(n_264),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_811),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_811),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_786),
.A2(n_326),
.B1(n_324),
.B2(n_322),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_778),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_SL g937 ( 
.A1(n_739),
.A2(n_319),
.B(n_318),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_741),
.B(n_265),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_739),
.A2(n_317),
.B(n_315),
.Y(n_939)
);

OAI21xp33_ASAP7_75t_SL g940 ( 
.A1(n_739),
.A2(n_64),
.B(n_65),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_754),
.Y(n_941)
);

OAI21xp33_ASAP7_75t_L g942 ( 
.A1(n_810),
.A2(n_65),
.B(n_66),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_748),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_786),
.A2(n_311),
.B1(n_309),
.B2(n_308),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_734),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_734),
.Y(n_946)
);

AOI222xp33_ASAP7_75t_L g947 ( 
.A1(n_840),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.C1(n_73),
.C2(n_74),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_853),
.A2(n_846),
.B(n_929),
.C(n_922),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_866),
.Y(n_949)
);

AO31x2_ASAP7_75t_L g950 ( 
.A1(n_822),
.A2(n_70),
.A3(n_71),
.B(n_73),
.Y(n_950)
);

NAND3xp33_ASAP7_75t_L g951 ( 
.A(n_873),
.B(n_74),
.C(n_75),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_825),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_871),
.A2(n_305),
.B1(n_303),
.B2(n_302),
.Y(n_953)
);

OAI221xp5_ASAP7_75t_L g954 ( 
.A1(n_861),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.C(n_78),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_943),
.B(n_77),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_941),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_917),
.B(n_267),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_843),
.B(n_79),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_939),
.A2(n_298),
.B(n_297),
.Y(n_959)
);

AO21x2_ASAP7_75t_L g960 ( 
.A1(n_852),
.A2(n_296),
.B(n_294),
.Y(n_960)
);

OR2x6_ASAP7_75t_L g961 ( 
.A(n_918),
.B(n_828),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_850),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_886),
.B(n_79),
.Y(n_963)
);

AO21x2_ASAP7_75t_L g964 ( 
.A1(n_883),
.A2(n_291),
.B(n_290),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_884),
.B(n_268),
.Y(n_965)
);

NOR2xp67_ASAP7_75t_L g966 ( 
.A(n_884),
.B(n_269),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_847),
.B(n_80),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_SL g968 ( 
.A1(n_891),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_849),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_917),
.B(n_281),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_830),
.A2(n_287),
.B(n_286),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_911),
.B(n_84),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_880),
.A2(n_285),
.B1(n_284),
.B2(n_283),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_914),
.A2(n_282),
.B(n_280),
.Y(n_974)
);

AO21x2_ASAP7_75t_L g975 ( 
.A1(n_836),
.A2(n_279),
.B(n_275),
.Y(n_975)
);

O2A1O1Ixp5_ASAP7_75t_L g976 ( 
.A1(n_826),
.A2(n_271),
.B(n_86),
.C(n_87),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_828),
.Y(n_977)
);

INVx6_ASAP7_75t_L g978 ( 
.A(n_915),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_940),
.A2(n_85),
.B(n_86),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_842),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_872),
.Y(n_981)
);

NAND2x1p5_ASAP7_75t_L g982 ( 
.A(n_834),
.B(n_87),
.Y(n_982)
);

NOR2xp67_ASAP7_75t_L g983 ( 
.A(n_839),
.B(n_88),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_834),
.B(n_89),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_829),
.B(n_90),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_887),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_942),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_823),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_SL g989 ( 
.A(n_837),
.B(n_94),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_SL g990 ( 
.A1(n_891),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_862),
.B(n_95),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_885),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_919),
.B(n_97),
.Y(n_993)
);

NAND2x1p5_ASAP7_75t_L g994 ( 
.A(n_834),
.B(n_98),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_927),
.B(n_99),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_SL g996 ( 
.A1(n_916),
.A2(n_901),
.B(n_855),
.C(n_869),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_931),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_876),
.Y(n_998)
);

NOR2x1_ASAP7_75t_SL g999 ( 
.A(n_885),
.B(n_133),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_845),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_928),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_844),
.A2(n_104),
.B(n_105),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_936),
.B(n_106),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_885),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_845),
.Y(n_1005)
);

NAND2x1p5_ASAP7_75t_L g1006 ( 
.A(n_931),
.B(n_107),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_905),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_937),
.A2(n_898),
.B(n_895),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_894),
.A2(n_109),
.B(n_110),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_896),
.A2(n_111),
.B(n_112),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_851),
.B(n_111),
.Y(n_1011)
);

AO21x2_ASAP7_75t_L g1012 ( 
.A1(n_924),
.A2(n_133),
.B(n_113),
.Y(n_1012)
);

OR2x6_ASAP7_75t_L g1013 ( 
.A(n_931),
.B(n_112),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_858),
.B(n_864),
.Y(n_1014)
);

CKINVDCx6p67_ASAP7_75t_R g1015 ( 
.A(n_839),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_877),
.B(n_114),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_910),
.Y(n_1017)
);

NOR2xp67_ASAP7_75t_L g1018 ( 
.A(n_839),
.B(n_117),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_899),
.A2(n_118),
.B(n_119),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_897),
.A2(n_121),
.B(n_122),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_SL g1021 ( 
.A1(n_857),
.A2(n_123),
.B(n_124),
.C(n_125),
.Y(n_1021)
);

CKINVDCx6p67_ASAP7_75t_R g1022 ( 
.A(n_856),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_SL g1023 ( 
.A1(n_854),
.A2(n_123),
.B(n_124),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_909),
.A2(n_125),
.B(n_126),
.C(n_127),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_930),
.B(n_126),
.Y(n_1025)
);

AO31x2_ASAP7_75t_L g1026 ( 
.A1(n_912),
.A2(n_128),
.A3(n_129),
.B(n_130),
.Y(n_1026)
);

NAND3xp33_ASAP7_75t_L g1027 ( 
.A(n_835),
.B(n_131),
.C(n_132),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_865),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_906),
.A2(n_913),
.B(n_920),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_946),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_902),
.B(n_832),
.Y(n_1031)
);

OAI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_888),
.A2(n_889),
.B1(n_824),
.B2(n_882),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_926),
.A2(n_932),
.B1(n_930),
.B2(n_938),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_879),
.B(n_938),
.Y(n_1034)
);

OA21x2_ASAP7_75t_L g1035 ( 
.A1(n_878),
.A2(n_875),
.B(n_890),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_915),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_832),
.B(n_827),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_848),
.B(n_908),
.Y(n_1038)
);

BUFx2_ASAP7_75t_SL g1039 ( 
.A(n_868),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_868),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_859),
.A2(n_893),
.B(n_907),
.C(n_867),
.Y(n_1041)
);

AO21x2_ASAP7_75t_L g1042 ( 
.A1(n_863),
.A2(n_900),
.B(n_870),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_921),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_848),
.B(n_833),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_923),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_841),
.A2(n_892),
.B1(n_903),
.B2(n_934),
.Y(n_1046)
);

AO21x2_ASAP7_75t_L g1047 ( 
.A1(n_874),
.A2(n_904),
.B(n_881),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_925),
.B(n_933),
.Y(n_1048)
);

CKINVDCx16_ASAP7_75t_R g1049 ( 
.A(n_941),
.Y(n_1049)
);

CKINVDCx14_ASAP7_75t_R g1050 ( 
.A(n_866),
.Y(n_1050)
);

AO21x2_ASAP7_75t_L g1051 ( 
.A1(n_853),
.A2(n_831),
.B(n_922),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_853),
.A2(n_825),
.B(n_831),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_917),
.B(n_930),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_838),
.A2(n_777),
.B(n_732),
.Y(n_1054)
);

NAND2x1p5_ASAP7_75t_L g1055 ( 
.A(n_918),
.B(n_945),
.Y(n_1055)
);

OA21x2_ASAP7_75t_L g1056 ( 
.A1(n_831),
.A2(n_853),
.B(n_922),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_861),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_838),
.A2(n_777),
.B(n_732),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_853),
.A2(n_825),
.B(n_831),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_853),
.A2(n_840),
.B(n_846),
.C(n_922),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_853),
.A2(n_739),
.B(n_831),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_849),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_828),
.Y(n_1063)
);

AO32x2_ASAP7_75t_L g1064 ( 
.A1(n_935),
.A2(n_758),
.A3(n_944),
.B1(n_787),
.B2(n_860),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_SL g1065 ( 
.A(n_884),
.Y(n_1065)
);

AO21x2_ASAP7_75t_L g1066 ( 
.A1(n_853),
.A2(n_831),
.B(n_922),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_861),
.B(n_748),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_850),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_838),
.A2(n_777),
.B(n_732),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_853),
.A2(n_825),
.B(n_831),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_969),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_952),
.B(n_1014),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_1057),
.Y(n_1073)
);

INVxp33_ASAP7_75t_L g1074 ( 
.A(n_1067),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_SL g1075 ( 
.A1(n_989),
.A2(n_954),
.B1(n_1010),
.B2(n_1033),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_1062),
.B(n_1001),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_958),
.B(n_985),
.Y(n_1077)
);

BUFx4f_ASAP7_75t_SL g1078 ( 
.A(n_956),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_961),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_1039),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_1028),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_962),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_961),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_1068),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_1022),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_977),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_988),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_955),
.B(n_1053),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_1053),
.B(n_1063),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_980),
.B(n_981),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_997),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_SL g1092 ( 
.A(n_949),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_967),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_998),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_1050),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_947),
.A2(n_987),
.B1(n_979),
.B2(n_1007),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_1060),
.B(n_1034),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1030),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1008),
.A2(n_1061),
.B(n_948),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_991),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_978),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1003),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_972),
.B(n_1025),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1025),
.B(n_993),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_963),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_952),
.B(n_1052),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_1011),
.B(n_1049),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_1044),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1054),
.A2(n_1058),
.B(n_1069),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_1040),
.Y(n_1110)
);

INVxp67_ASAP7_75t_SL g1111 ( 
.A(n_1059),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1070),
.B(n_1051),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_995),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1017),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1017),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_957),
.B(n_970),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1038),
.B(n_1031),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1016),
.B(n_1013),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1013),
.B(n_968),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_1000),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1019),
.A2(n_959),
.B(n_1056),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1005),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1055),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_978),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_951),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1021),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1066),
.B(n_1029),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1027),
.Y(n_1128)
);

INVxp67_ASAP7_75t_L g1129 ( 
.A(n_1023),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_999),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_990),
.B(n_1046),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_999),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1032),
.B(n_1056),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_1036),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1048),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1041),
.B(n_996),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_982),
.B(n_1006),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_986),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_984),
.B(n_994),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_950),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1037),
.B(n_1045),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1043),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1047),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_965),
.B(n_966),
.Y(n_1144)
);

INVx6_ASAP7_75t_L g1145 ( 
.A(n_1049),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_SL g1146 ( 
.A1(n_1048),
.A2(n_953),
.B1(n_1004),
.B2(n_992),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1020),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1015),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_1065),
.Y(n_1149)
);

CKINVDCx6p67_ASAP7_75t_R g1150 ( 
.A(n_1065),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1042),
.A2(n_1035),
.B1(n_975),
.B2(n_1012),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1107),
.B(n_960),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1104),
.B(n_1018),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1103),
.B(n_983),
.Y(n_1154)
);

INVx5_ASAP7_75t_L g1155 ( 
.A(n_1081),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1074),
.B(n_1024),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_1084),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1074),
.B(n_1012),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1116),
.B(n_964),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1084),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_1071),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_1071),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1088),
.B(n_1026),
.Y(n_1163)
);

INVxp67_ASAP7_75t_L g1164 ( 
.A(n_1073),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1097),
.B(n_1026),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1117),
.B(n_1009),
.Y(n_1166)
);

NOR2x1_ASAP7_75t_L g1167 ( 
.A(n_1072),
.B(n_973),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_1076),
.B(n_971),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1113),
.B(n_1077),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1077),
.B(n_974),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1116),
.B(n_976),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1097),
.B(n_1002),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1131),
.B(n_1064),
.Y(n_1173)
);

INVxp67_ASAP7_75t_SL g1174 ( 
.A(n_1136),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1087),
.B(n_1064),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1105),
.B(n_1108),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1100),
.B(n_1102),
.Y(n_1177)
);

BUFx2_ASAP7_75t_R g1178 ( 
.A(n_1095),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_1082),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1114),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1115),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1118),
.B(n_1093),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1093),
.B(n_1141),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1125),
.B(n_1128),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1119),
.B(n_1137),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1090),
.B(n_1086),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1139),
.B(n_1094),
.Y(n_1187)
);

OR2x6_ASAP7_75t_L g1188 ( 
.A(n_1145),
.B(n_1136),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1124),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1143),
.Y(n_1190)
);

CKINVDCx14_ASAP7_75t_R g1191 ( 
.A(n_1095),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1106),
.B(n_1111),
.Y(n_1192)
);

OR2x2_ASAP7_75t_SL g1193 ( 
.A(n_1145),
.B(n_1079),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1143),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_1086),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_SL g1196 ( 
.A1(n_1096),
.A2(n_1075),
.B(n_1099),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1091),
.B(n_1106),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1075),
.B(n_1138),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1133),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1096),
.B(n_1080),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_1110),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1098),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1147),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1079),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1091),
.B(n_1120),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1080),
.B(n_1112),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1133),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1122),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1083),
.B(n_1142),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1146),
.A2(n_1099),
.B1(n_1126),
.B2(n_1121),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1112),
.B(n_1089),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1089),
.B(n_1083),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1165),
.B(n_1140),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1188),
.B(n_1159),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1195),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_1186),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1180),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1181),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1193),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1190),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1169),
.B(n_1145),
.Y(n_1221)
);

INVxp67_ASAP7_75t_SL g1222 ( 
.A(n_1195),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1200),
.B(n_1129),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1189),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1173),
.B(n_1127),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1163),
.B(n_1151),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1175),
.B(n_1151),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1199),
.B(n_1207),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1203),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1203),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1175),
.B(n_1121),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1177),
.B(n_1078),
.Y(n_1232)
);

INVxp33_ASAP7_75t_L g1233 ( 
.A(n_1183),
.Y(n_1233)
);

NAND2xp33_ASAP7_75t_R g1234 ( 
.A(n_1188),
.B(n_1132),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1159),
.B(n_1130),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1176),
.B(n_1184),
.Y(n_1236)
);

INVxp33_ASAP7_75t_L g1237 ( 
.A(n_1187),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1176),
.B(n_1078),
.Y(n_1238)
);

NOR2x1_ASAP7_75t_L g1239 ( 
.A(n_1206),
.B(n_1170),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1167),
.B(n_1144),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1160),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1198),
.B(n_1123),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1158),
.B(n_1109),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1204),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1220),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1229),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1239),
.B(n_1192),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1229),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1216),
.B(n_1211),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1244),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1231),
.B(n_1190),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1230),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1235),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1228),
.B(n_1194),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1230),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1236),
.B(n_1196),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1223),
.B(n_1197),
.Y(n_1257)
);

AND2x2_ASAP7_75t_SL g1258 ( 
.A(n_1214),
.B(n_1210),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1227),
.B(n_1172),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1240),
.A2(n_1156),
.B1(n_1210),
.B2(n_1171),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1232),
.B(n_1179),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1227),
.B(n_1172),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1226),
.B(n_1194),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1226),
.B(n_1225),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1225),
.B(n_1152),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1220),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1233),
.B(n_1161),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1213),
.B(n_1166),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1245),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1266),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1249),
.B(n_1215),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1264),
.B(n_1243),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1246),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1251),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1247),
.B(n_1222),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1246),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1248),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1260),
.A2(n_1240),
.B1(n_1219),
.B2(n_1214),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1248),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1253),
.B(n_1214),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1252),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1264),
.B(n_1243),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1263),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1258),
.A2(n_1234),
.B1(n_1144),
.B2(n_1159),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1255),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1257),
.B(n_1217),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1252),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1265),
.B(n_1241),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1251),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1258),
.A2(n_1174),
.B(n_1237),
.C(n_1234),
.Y(n_1290)
);

OAI211xp5_ASAP7_75t_L g1291 ( 
.A1(n_1256),
.A2(n_1242),
.B(n_1164),
.C(n_1221),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1273),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1284),
.A2(n_1261),
.B1(n_1253),
.B2(n_1259),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1276),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1288),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1277),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1290),
.A2(n_1237),
.B1(n_1250),
.B2(n_1174),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1279),
.Y(n_1298)
);

INVxp33_ASAP7_75t_L g1299 ( 
.A(n_1271),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1281),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1285),
.Y(n_1301)
);

AOI32xp33_ASAP7_75t_L g1302 ( 
.A1(n_1269),
.A2(n_1262),
.A3(n_1259),
.B1(n_1263),
.B2(n_1268),
.Y(n_1302)
);

AOI222xp33_ASAP7_75t_L g1303 ( 
.A1(n_1291),
.A2(n_1182),
.B1(n_1153),
.B2(n_1154),
.C1(n_1185),
.C2(n_1162),
.Y(n_1303)
);

INVxp67_ASAP7_75t_L g1304 ( 
.A(n_1270),
.Y(n_1304)
);

O2A1O1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1290),
.A2(n_1212),
.B(n_1168),
.C(n_1267),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1287),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1285),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1272),
.B(n_1262),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1292),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1308),
.B(n_1282),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1297),
.A2(n_1278),
.B1(n_1280),
.B2(n_1275),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1294),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1296),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1299),
.B(n_1274),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_1298),
.Y(n_1315)
);

AOI221x1_ASAP7_75t_L g1316 ( 
.A1(n_1312),
.A2(n_1297),
.B1(n_1313),
.B2(n_1314),
.C(n_1306),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1311),
.B(n_1305),
.C(n_1303),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1315),
.A2(n_1305),
.B(n_1309),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1309),
.A2(n_1303),
.B(n_1286),
.Y(n_1319)
);

AOI222xp33_ASAP7_75t_L g1320 ( 
.A1(n_1310),
.A2(n_1304),
.B1(n_1283),
.B2(n_1238),
.C1(n_1274),
.C2(n_1289),
.Y(n_1320)
);

NOR3x1_ASAP7_75t_L g1321 ( 
.A(n_1317),
.B(n_1101),
.C(n_1148),
.Y(n_1321)
);

NAND4xp25_ASAP7_75t_L g1322 ( 
.A(n_1316),
.B(n_1293),
.C(n_1302),
.D(n_1209),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1319),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1318),
.B(n_1295),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1320),
.B(n_1280),
.Y(n_1325)
);

NOR3x1_ASAP7_75t_L g1326 ( 
.A(n_1317),
.B(n_1085),
.C(n_1157),
.Y(n_1326)
);

NOR3x1_ASAP7_75t_L g1327 ( 
.A(n_1317),
.B(n_1157),
.C(n_1178),
.Y(n_1327)
);

NOR3xp33_ASAP7_75t_L g1328 ( 
.A(n_1317),
.B(n_1191),
.C(n_1149),
.Y(n_1328)
);

NOR2x1_ASAP7_75t_L g1329 ( 
.A(n_1322),
.B(n_1134),
.Y(n_1329)
);

NOR2x1_ASAP7_75t_L g1330 ( 
.A(n_1323),
.B(n_1134),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1324),
.Y(n_1331)
);

AOI211xp5_ASAP7_75t_L g1332 ( 
.A1(n_1328),
.A2(n_1149),
.B(n_1124),
.C(n_1135),
.Y(n_1332)
);

NOR3x1_ASAP7_75t_L g1333 ( 
.A(n_1325),
.B(n_1092),
.C(n_1201),
.Y(n_1333)
);

NOR3xp33_ASAP7_75t_L g1334 ( 
.A(n_1327),
.B(n_1191),
.C(n_1135),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1321),
.B(n_1326),
.Y(n_1335)
);

NOR2x1_ASAP7_75t_L g1336 ( 
.A(n_1322),
.B(n_1160),
.Y(n_1336)
);

AND3x4_ASAP7_75t_L g1337 ( 
.A(n_1334),
.B(n_1189),
.C(n_1092),
.Y(n_1337)
);

XOR2x1_ASAP7_75t_L g1338 ( 
.A(n_1331),
.B(n_1150),
.Y(n_1338)
);

NOR3x2_ASAP7_75t_L g1339 ( 
.A(n_1330),
.B(n_1155),
.C(n_1254),
.Y(n_1339)
);

NOR3xp33_ASAP7_75t_SL g1340 ( 
.A(n_1333),
.B(n_1329),
.C(n_1336),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1335),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1341),
.B(n_1300),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1340),
.B(n_1332),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1338),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_1339),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1345),
.Y(n_1346)
);

OAI211xp5_ASAP7_75t_L g1347 ( 
.A1(n_1343),
.A2(n_1344),
.B(n_1345),
.C(n_1342),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1343),
.B(n_1301),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1342),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1346),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1349),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1348),
.Y(n_1352)
);

XNOR2xp5_ASAP7_75t_L g1353 ( 
.A(n_1350),
.B(n_1337),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1352),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1351),
.A2(n_1347),
.B1(n_1283),
.B2(n_1224),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1353),
.A2(n_1354),
.B(n_1355),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1353),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1357),
.A2(n_1224),
.B1(n_1289),
.B2(n_1307),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1358),
.A2(n_1356),
.B(n_1205),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1359),
.B(n_1218),
.Y(n_1360)
);

AOI21xp33_ASAP7_75t_L g1361 ( 
.A1(n_1360),
.A2(n_1202),
.B(n_1208),
.Y(n_1361)
);


endmodule