module fake_netlist_6_2782_n_1078 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_258, n_154, n_191, n_88, n_3, n_209, n_98, n_260, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_255, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1078);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_258;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_260;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_255;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1078;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_898;
wire n_617;
wire n_698;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_843;
wire n_772;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_934;
wire n_482;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_689;
wire n_354;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_84),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_152),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_17),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_103),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_110),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_98),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_160),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_105),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_13),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_82),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_77),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_232),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_222),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_255),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_6),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_208),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_137),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_240),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_168),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_46),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_171),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_43),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_16),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_7),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_223),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_71),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_163),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_49),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_155),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_37),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_104),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_118),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_68),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_261),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_95),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_237),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_73),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_18),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_116),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_206),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_177),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_178),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_200),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_187),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_197),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_102),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_212),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_86),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_166),
.Y(n_313)
);

BUFx8_ASAP7_75t_SL g314 ( 
.A(n_91),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_153),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_80),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_184),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_79),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_45),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_251),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_121),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_211),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_143),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_16),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_146),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_227),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_265),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_278),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_271),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_275),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_286),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_275),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_295),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_295),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_301),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_292),
.B(n_289),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_324),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_0),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_314),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_325),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_266),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_269),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_273),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_291),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_274),
.Y(n_346)
);

NOR2xp67_ASAP7_75t_L g347 ( 
.A(n_276),
.B(n_0),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_279),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_314),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_263),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_284),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_288),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_297),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_290),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_264),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_299),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_303),
.B(n_1),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_305),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_309),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_321),
.B(n_1),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_318),
.B(n_2),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_264),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_298),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_313),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_267),
.B(n_2),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_366),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_328),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_343),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_355),
.Y(n_373)
);

OAI21x1_ASAP7_75t_L g374 ( 
.A1(n_355),
.A2(n_313),
.B(n_302),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_344),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_334),
.Y(n_376)
);

AND2x6_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_264),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_332),
.B(n_3),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_336),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_337),
.B(n_268),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_334),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_342),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_335),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_361),
.A2(n_320),
.B1(n_312),
.B2(n_270),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_336),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_327),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_330),
.B(n_272),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_348),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_357),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_359),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_277),
.Y(n_398)
);

OA21x2_ASAP7_75t_L g399 ( 
.A1(n_362),
.A2(n_281),
.B(n_280),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_365),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_341),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_358),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_358),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_368),
.B(n_282),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_347),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_331),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_350),
.B(n_323),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_333),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_340),
.B(n_264),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_364),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_340),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_363),
.B(n_283),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_353),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_400),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_285),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_405),
.B(n_302),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_372),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_375),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_404),
.B(n_293),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_294),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_409),
.B(n_349),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_382),
.B(n_296),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_392),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_401),
.B(n_306),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_396),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_397),
.Y(n_431)
);

AND2x6_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_302),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_307),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_387),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_387),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_379),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_373),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_353),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_308),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_400),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_380),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_310),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_394),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_379),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_R g449 ( 
.A(n_412),
.B(n_367),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_400),
.Y(n_450)
);

BUFx4f_ASAP7_75t_L g451 ( 
.A(n_405),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_400),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_404),
.B(n_311),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_404),
.B(n_315),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_390),
.B(n_316),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_416),
.B(n_317),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_376),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_389),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_389),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_393),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_393),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_412),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_398),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

INVx6_ASAP7_75t_L g466 ( 
.A(n_378),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_376),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_395),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_371),
.B(n_319),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_376),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_384),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_376),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_390),
.B(n_367),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_378),
.B(n_322),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_391),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_411),
.B(n_302),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_381),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_391),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_402),
.B(n_36),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_410),
.B(n_38),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_373),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_391),
.Y(n_482)
);

OAI22xp33_ASAP7_75t_L g483 ( 
.A1(n_411),
.A2(n_414),
.B1(n_408),
.B2(n_385),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_370),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_442),
.B(n_411),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_442),
.B(n_399),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_471),
.A2(n_338),
.B1(n_388),
.B2(n_418),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_481),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_434),
.Y(n_489)
);

AO22x2_ASAP7_75t_L g490 ( 
.A1(n_447),
.A2(n_414),
.B1(n_398),
.B2(n_413),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_481),
.Y(n_491)
);

AO22x2_ASAP7_75t_L g492 ( 
.A1(n_476),
.A2(n_415),
.B1(n_412),
.B2(n_338),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_449),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_435),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_449),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_438),
.Y(n_496)
);

CKINVDCx14_ASAP7_75t_R g497 ( 
.A(n_426),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_443),
.Y(n_498)
);

OR2x6_ASAP7_75t_L g499 ( 
.A(n_463),
.B(n_418),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_427),
.B(n_399),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_427),
.B(n_399),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_437),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_454),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_473),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_469),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_477),
.B(n_406),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_475),
.Y(n_507)
);

AO22x2_ASAP7_75t_L g508 ( 
.A1(n_476),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_445),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_477),
.B(n_457),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_457),
.B(n_418),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_474),
.B(n_418),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_422),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_423),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_459),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_469),
.B(n_418),
.Y(n_516)
);

BUFx8_ASAP7_75t_L g517 ( 
.A(n_436),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_428),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_460),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_430),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_454),
.B(n_370),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_444),
.Y(n_522)
);

NAND2x1p5_ASAP7_75t_L g523 ( 
.A(n_441),
.B(n_374),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_441),
.B(n_381),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_464),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_431),
.B(n_484),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_461),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_462),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_465),
.Y(n_529)
);

NAND2x1p5_ASAP7_75t_L g530 ( 
.A(n_451),
.B(n_374),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_466),
.A2(n_377),
.B1(n_386),
.B2(n_383),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_478),
.B(n_377),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_482),
.Y(n_533)
);

AO22x2_ASAP7_75t_L g534 ( 
.A1(n_424),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_534)
);

AO22x2_ASAP7_75t_L g535 ( 
.A1(n_424),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_468),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_420),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_453),
.B(n_377),
.Y(n_538)
);

AO22x2_ASAP7_75t_L g539 ( 
.A1(n_455),
.A2(n_421),
.B1(n_483),
.B2(n_456),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_466),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_466),
.Y(n_541)
);

NAND2x1p5_ASAP7_75t_L g542 ( 
.A(n_451),
.B(n_383),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_425),
.B(n_377),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_425),
.B(n_377),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_455),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_421),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_429),
.B(n_377),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_448),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_448),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_483),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_433),
.B(n_439),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_480),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_458),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_458),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_440),
.B(n_386),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_440),
.B(n_373),
.Y(n_556)
);

AO22x2_ASAP7_75t_L g557 ( 
.A1(n_467),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_505),
.B(n_419),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_SL g559 ( 
.A(n_550),
.B(n_388),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_522),
.B(n_419),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_511),
.B(n_419),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_537),
.B(n_516),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_510),
.B(n_446),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_485),
.B(n_419),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_506),
.B(n_452),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_540),
.B(n_452),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_541),
.B(n_446),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_525),
.B(n_450),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_526),
.B(n_450),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_526),
.B(n_479),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_SL g571 ( 
.A(n_512),
.B(n_467),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_552),
.B(n_432),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_503),
.B(n_472),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_503),
.B(n_472),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_545),
.B(n_470),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_524),
.B(n_470),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_SL g577 ( 
.A(n_493),
.B(n_432),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_524),
.B(n_432),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_496),
.B(n_432),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_551),
.B(n_432),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_513),
.B(n_39),
.Y(n_581)
);

NAND2xp33_ASAP7_75t_SL g582 ( 
.A(n_504),
.B(n_10),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_487),
.B(n_11),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_489),
.B(n_11),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_SL g585 ( 
.A(n_486),
.B(n_514),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_494),
.B(n_12),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_498),
.B(n_12),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_518),
.B(n_40),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_499),
.B(n_13),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_520),
.B(n_41),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_SL g591 ( 
.A(n_509),
.B(n_14),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_495),
.B(n_42),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_515),
.B(n_44),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_519),
.B(n_47),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_527),
.B(n_48),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_529),
.B(n_50),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_521),
.B(n_51),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_528),
.B(n_536),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_536),
.B(n_52),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_542),
.B(n_53),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_500),
.B(n_54),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_501),
.B(n_55),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_507),
.B(n_56),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_SL g604 ( 
.A(n_546),
.B(n_14),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_507),
.B(n_15),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_533),
.B(n_57),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_533),
.B(n_58),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_543),
.B(n_59),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_499),
.B(n_15),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_544),
.B(n_60),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_502),
.B(n_555),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_538),
.B(n_17),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_531),
.B(n_61),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_488),
.B(n_62),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_491),
.B(n_530),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_SL g616 ( 
.A(n_547),
.B(n_18),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_539),
.B(n_19),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_539),
.B(n_549),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_553),
.B(n_63),
.Y(n_619)
);

AND2x2_ASAP7_75t_SL g620 ( 
.A(n_554),
.B(n_64),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_561),
.A2(n_523),
.B(n_532),
.Y(n_621)
);

AO31x2_ASAP7_75t_L g622 ( 
.A1(n_618),
.A2(n_548),
.A3(n_556),
.B(n_492),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_R g623 ( 
.A(n_577),
.B(n_497),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_570),
.A2(n_490),
.B(n_492),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_609),
.Y(n_625)
);

A2O1A1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_562),
.A2(n_490),
.B(n_535),
.C(n_534),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_559),
.B(n_517),
.Y(n_627)
);

AO31x2_ASAP7_75t_L g628 ( 
.A1(n_617),
.A2(n_508),
.A3(n_557),
.B(n_534),
.Y(n_628)
);

INVx4_ASAP7_75t_SL g629 ( 
.A(n_589),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_598),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_580),
.A2(n_508),
.B(n_557),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_585),
.A2(n_535),
.B(n_66),
.Y(n_632)
);

NOR2x1_ASAP7_75t_SL g633 ( 
.A(n_600),
.B(n_65),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_588),
.B(n_517),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_605),
.Y(n_635)
);

NAND3xp33_ASAP7_75t_L g636 ( 
.A(n_583),
.B(n_582),
.C(n_591),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_576),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_588),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_611),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_L g640 ( 
.A1(n_601),
.A2(n_69),
.B(n_67),
.Y(n_640)
);

AOI221x1_ASAP7_75t_L g641 ( 
.A1(n_612),
.A2(n_616),
.B1(n_604),
.B2(n_571),
.C(n_563),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_584),
.B(n_19),
.Y(n_642)
);

AOI31xp67_ASAP7_75t_L g643 ( 
.A1(n_602),
.A2(n_167),
.A3(n_260),
.B(n_259),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_615),
.A2(n_72),
.B(n_70),
.Y(n_644)
);

AOI221x1_ASAP7_75t_L g645 ( 
.A1(n_586),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.C(n_23),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_565),
.A2(n_75),
.B(n_74),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_573),
.A2(n_574),
.B(n_575),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_608),
.A2(n_78),
.B(n_76),
.Y(n_648)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_610),
.A2(n_83),
.B(n_81),
.Y(n_649)
);

OAI21x1_ASAP7_75t_L g650 ( 
.A1(n_579),
.A2(n_87),
.B(n_85),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_588),
.B(n_88),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_568),
.B(n_89),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_587),
.B(n_20),
.Y(n_653)
);

AO31x2_ASAP7_75t_L g654 ( 
.A1(n_572),
.A2(n_175),
.A3(n_258),
.B(n_257),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_564),
.A2(n_92),
.B(n_90),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_567),
.B(n_21),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_L g657 ( 
.A(n_592),
.B(n_22),
.C(n_23),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_578),
.A2(n_94),
.B(n_93),
.Y(n_658)
);

OAI21xp5_ASAP7_75t_L g659 ( 
.A1(n_613),
.A2(n_97),
.B(n_96),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_569),
.A2(n_597),
.B(n_560),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_620),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_L g662 ( 
.A(n_603),
.B(n_99),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_558),
.B(n_24),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_620),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_566),
.B(n_100),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_606),
.B(n_101),
.Y(n_666)
);

AND2x6_ASAP7_75t_L g667 ( 
.A(n_581),
.B(n_106),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_607),
.B(n_24),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_599),
.B(n_25),
.Y(n_669)
);

AO31x2_ASAP7_75t_L g670 ( 
.A1(n_619),
.A2(n_185),
.A3(n_256),
.B(n_254),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_614),
.A2(n_590),
.B(n_593),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_594),
.A2(n_108),
.B(n_107),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_595),
.B(n_25),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_596),
.A2(n_186),
.B1(n_253),
.B2(n_252),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_562),
.B(n_26),
.Y(n_675)
);

AO32x2_ASAP7_75t_L g676 ( 
.A1(n_617),
.A2(n_26),
.A3(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_562),
.B(n_27),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_609),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_562),
.B(n_28),
.Y(n_679)
);

NOR4xp25_ASAP7_75t_L g680 ( 
.A(n_562),
.B(n_29),
.C(n_30),
.D(n_31),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_SL g681 ( 
.A1(n_661),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_678),
.Y(n_682)
);

OA21x2_ASAP7_75t_L g683 ( 
.A1(n_641),
.A2(n_189),
.B(n_249),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_630),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_625),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_621),
.A2(n_188),
.B(n_248),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_647),
.A2(n_183),
.B(n_247),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_636),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_635),
.B(n_33),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_650),
.A2(n_190),
.B(n_246),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_639),
.Y(n_691)
);

OA21x2_ASAP7_75t_L g692 ( 
.A1(n_624),
.A2(n_182),
.B(n_245),
.Y(n_692)
);

OA21x2_ASAP7_75t_L g693 ( 
.A1(n_631),
.A2(n_181),
.B(n_244),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_625),
.Y(n_694)
);

INVx4_ASAP7_75t_SL g695 ( 
.A(n_667),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_678),
.Y(n_696)
);

OAI21x1_ASAP7_75t_SL g697 ( 
.A1(n_633),
.A2(n_180),
.B(n_243),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_637),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_629),
.B(n_34),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_675),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_664),
.B(n_35),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_623),
.B(n_109),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_677),
.A2(n_35),
.B(n_111),
.C(n_112),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_638),
.B(n_113),
.Y(n_704)
);

OA21x2_ASAP7_75t_L g705 ( 
.A1(n_660),
.A2(n_114),
.B(n_115),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_629),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_627),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_656),
.Y(n_708)
);

AO21x2_ASAP7_75t_L g709 ( 
.A1(n_640),
.A2(n_117),
.B(n_119),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_644),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_626),
.A2(n_120),
.B(n_122),
.C(n_123),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_634),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_712)
);

AO21x1_ASAP7_75t_L g713 ( 
.A1(n_632),
.A2(n_127),
.B(n_128),
.Y(n_713)
);

OAI21x1_ASAP7_75t_L g714 ( 
.A1(n_649),
.A2(n_129),
.B(n_130),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_665),
.B(n_262),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_663),
.Y(n_716)
);

BUFx12f_ASAP7_75t_L g717 ( 
.A(n_679),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_651),
.A2(n_662),
.B(n_659),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_652),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_652),
.Y(n_720)
);

O2A1O1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_642),
.A2(n_131),
.B(n_132),
.C(n_133),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_657),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_722)
);

AO21x2_ASAP7_75t_L g723 ( 
.A1(n_648),
.A2(n_138),
.B(n_139),
.Y(n_723)
);

INVxp67_ASAP7_75t_SL g724 ( 
.A(n_665),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_SL g725 ( 
.A1(n_666),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_666),
.B(n_242),
.Y(n_726)
);

CKINVDCx16_ASAP7_75t_R g727 ( 
.A(n_673),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_667),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_628),
.B(n_144),
.Y(n_729)
);

AO21x2_ASAP7_75t_L g730 ( 
.A1(n_653),
.A2(n_145),
.B(n_147),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_622),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_628),
.B(n_148),
.Y(n_732)
);

AOI211xp5_ASAP7_75t_L g733 ( 
.A1(n_680),
.A2(n_149),
.B(n_150),
.C(n_151),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_622),
.Y(n_734)
);

AO31x2_ASAP7_75t_L g735 ( 
.A1(n_645),
.A2(n_154),
.A3(n_156),
.B(n_157),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_719),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_684),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_682),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_691),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_686),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_698),
.Y(n_741)
);

OAI21xp5_ASAP7_75t_L g742 ( 
.A1(n_718),
.A2(n_668),
.B(n_669),
.Y(n_742)
);

INVx4_ASAP7_75t_SL g743 ( 
.A(n_735),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_731),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_719),
.B(n_676),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_734),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_683),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_683),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_706),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_694),
.Y(n_750)
);

XNOR2xp5_ASAP7_75t_L g751 ( 
.A(n_708),
.B(n_674),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_705),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_705),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_729),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_710),
.Y(n_755)
);

OA21x2_ASAP7_75t_L g756 ( 
.A1(n_729),
.A2(n_732),
.B(n_687),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_685),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_732),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_735),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_716),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_700),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_720),
.B(n_676),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_701),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_735),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_693),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_714),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_693),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_692),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_717),
.A2(n_667),
.B1(n_655),
.B2(n_646),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_692),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_720),
.A2(n_672),
.B1(n_658),
.B2(n_671),
.Y(n_771)
);

AO21x2_ASAP7_75t_L g772 ( 
.A1(n_718),
.A2(n_643),
.B(n_654),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_724),
.Y(n_773)
);

AOI21x1_ASAP7_75t_L g774 ( 
.A1(n_713),
.A2(n_654),
.B(n_670),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_690),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_SL g776 ( 
.A1(n_733),
.A2(n_670),
.B(n_159),
.C(n_161),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_709),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_730),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_708),
.B(n_158),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_709),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_701),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_727),
.B(n_241),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_707),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_696),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_723),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_728),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_723),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_730),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_726),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_726),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_711),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_704),
.B(n_162),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_697),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_711),
.Y(n_794)
);

NAND2x1p5_ASAP7_75t_L g795 ( 
.A(n_715),
.B(n_704),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_695),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_795),
.B(n_715),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_763),
.B(n_689),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_SL g799 ( 
.A(n_783),
.B(n_699),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_738),
.B(n_749),
.Y(n_800)
);

OR2x6_ASAP7_75t_L g801 ( 
.A(n_795),
.B(n_721),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_781),
.B(n_688),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_R g803 ( 
.A(n_786),
.B(n_695),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_R g804 ( 
.A(n_786),
.B(n_702),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_737),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_738),
.B(n_695),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_737),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_750),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_746),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_781),
.B(n_681),
.Y(n_810)
);

OR2x6_ASAP7_75t_L g811 ( 
.A(n_795),
.B(n_721),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_R g812 ( 
.A(n_782),
.B(n_164),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_R g813 ( 
.A(n_751),
.B(n_165),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_749),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_789),
.B(n_712),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_R g816 ( 
.A(n_751),
.B(n_169),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_790),
.B(n_703),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_746),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_739),
.B(n_722),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_784),
.B(n_170),
.Y(n_820)
);

BUFx4f_ASAP7_75t_L g821 ( 
.A(n_796),
.Y(n_821)
);

OR2x6_ASAP7_75t_L g822 ( 
.A(n_773),
.B(n_725),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_R g823 ( 
.A(n_796),
.B(n_172),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_R g824 ( 
.A(n_773),
.B(n_173),
.Y(n_824)
);

NAND2xp33_ASAP7_75t_R g825 ( 
.A(n_792),
.B(n_174),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_760),
.B(n_733),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_R g827 ( 
.A(n_736),
.B(n_176),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_739),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_757),
.B(n_179),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_736),
.B(n_191),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_761),
.Y(n_831)
);

OR2x6_ASAP7_75t_L g832 ( 
.A(n_736),
.B(n_192),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_779),
.B(n_193),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_741),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_736),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_R g836 ( 
.A(n_792),
.B(n_194),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_736),
.B(n_195),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_R g838 ( 
.A(n_754),
.B(n_239),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_R g839 ( 
.A(n_756),
.B(n_754),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_793),
.B(n_196),
.Y(n_840)
);

XOR2xp5_ASAP7_75t_L g841 ( 
.A(n_769),
.B(n_198),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_742),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_R g843 ( 
.A(n_756),
.B(n_199),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_R g844 ( 
.A(n_758),
.B(n_238),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_745),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_793),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_744),
.Y(n_847)
);

OR2x6_ASAP7_75t_L g848 ( 
.A(n_745),
.B(n_762),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_805),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_809),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_846),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_828),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_842),
.A2(n_794),
.B1(n_791),
.B2(n_758),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_841),
.A2(n_794),
.B1(n_791),
.B2(n_771),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_818),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_848),
.B(n_759),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_831),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_848),
.B(n_743),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_807),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_834),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_845),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_847),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_808),
.B(n_755),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_826),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_817),
.B(n_759),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_801),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_801),
.B(n_764),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_811),
.B(n_743),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_814),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_802),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_811),
.B(n_764),
.Y(n_871)
);

NAND2x1p5_ASAP7_75t_SL g872 ( 
.A(n_835),
.B(n_777),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_819),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_798),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_810),
.B(n_788),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_822),
.B(n_788),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_797),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_840),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_840),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_825),
.A2(n_787),
.B1(n_785),
.B2(n_780),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_822),
.B(n_743),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_839),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_800),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_829),
.B(n_755),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_806),
.B(n_743),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_832),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_832),
.B(n_778),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_830),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_821),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_838),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_815),
.B(n_778),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_837),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_820),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_844),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_833),
.B(n_756),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_799),
.B(n_813),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_803),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_827),
.B(n_756),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_816),
.B(n_787),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_823),
.B(n_785),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_843),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_869),
.Y(n_902)
);

OAI33xp33_ASAP7_75t_L g903 ( 
.A1(n_870),
.A2(n_874),
.A3(n_875),
.B1(n_853),
.B2(n_882),
.B3(n_863),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_882),
.B(n_875),
.Y(n_904)
);

AND2x4_ASAP7_75t_SL g905 ( 
.A(n_886),
.B(n_824),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_865),
.B(n_867),
.Y(n_906)
);

NOR2x1_ASAP7_75t_L g907 ( 
.A(n_874),
.B(n_777),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_857),
.Y(n_908)
);

OAI221xp5_ASAP7_75t_L g909 ( 
.A1(n_880),
.A2(n_836),
.B1(n_812),
.B2(n_776),
.C(n_740),
.Y(n_909)
);

NAND3xp33_ASAP7_75t_L g910 ( 
.A(n_854),
.B(n_765),
.C(n_775),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_867),
.B(n_748),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_871),
.B(n_748),
.Y(n_912)
);

AND2x2_ASAP7_75t_SL g913 ( 
.A(n_858),
.B(n_747),
.Y(n_913)
);

OR2x2_ASAP7_75t_L g914 ( 
.A(n_856),
.B(n_765),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_871),
.B(n_747),
.Y(n_915)
);

AOI221xp5_ASAP7_75t_L g916 ( 
.A1(n_895),
.A2(n_804),
.B1(n_768),
.B2(n_772),
.C(n_752),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_860),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_864),
.B(n_772),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_850),
.Y(n_919)
);

OAI221xp5_ASAP7_75t_L g920 ( 
.A1(n_896),
.A2(n_740),
.B1(n_766),
.B2(n_775),
.C(n_768),
.Y(n_920)
);

OAI31xp33_ASAP7_75t_L g921 ( 
.A1(n_890),
.A2(n_740),
.A3(n_766),
.B(n_767),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_860),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_878),
.A2(n_886),
.B1(n_879),
.B2(n_894),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_873),
.B(n_767),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_864),
.B(n_772),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_873),
.B(n_770),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_849),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_891),
.B(n_858),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_889),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_878),
.A2(n_766),
.B1(n_770),
.B2(n_753),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_891),
.B(n_858),
.Y(n_931)
);

AO21x2_ASAP7_75t_L g932 ( 
.A1(n_872),
.A2(n_752),
.B(n_753),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_851),
.Y(n_933)
);

AO21x2_ASAP7_75t_L g934 ( 
.A1(n_872),
.A2(n_774),
.B(n_202),
.Y(n_934)
);

NAND3xp33_ASAP7_75t_L g935 ( 
.A(n_901),
.B(n_774),
.C(n_203),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_856),
.B(n_201),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_849),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_908),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_919),
.Y(n_939)
);

AND3x2_ASAP7_75t_L g940 ( 
.A(n_936),
.B(n_890),
.C(n_889),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_927),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_917),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_906),
.B(n_866),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_906),
.B(n_928),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_904),
.B(n_901),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_933),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_917),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_927),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_937),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_928),
.B(n_866),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_937),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_931),
.B(n_898),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_904),
.B(n_861),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_914),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_931),
.B(n_898),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_922),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_913),
.B(n_868),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_914),
.B(n_876),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_922),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_913),
.B(n_868),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_911),
.B(n_868),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_911),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_912),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_912),
.B(n_877),
.Y(n_964)
);

AO221x2_ASAP7_75t_L g965 ( 
.A1(n_945),
.A2(n_910),
.B1(n_935),
.B2(n_953),
.C(n_879),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_938),
.B(n_916),
.Y(n_966)
);

OAI22xp33_ASAP7_75t_L g967 ( 
.A1(n_958),
.A2(n_909),
.B1(n_886),
.B2(n_923),
.Y(n_967)
);

OAI22xp33_ASAP7_75t_L g968 ( 
.A1(n_958),
.A2(n_876),
.B1(n_877),
.B2(n_929),
.Y(n_968)
);

AO221x1_ASAP7_75t_L g969 ( 
.A1(n_946),
.A2(n_851),
.B1(n_897),
.B2(n_903),
.C(n_850),
.Y(n_969)
);

AO221x2_ASAP7_75t_L g970 ( 
.A1(n_963),
.A2(n_883),
.B1(n_905),
.B2(n_893),
.C(n_892),
.Y(n_970)
);

NAND2xp33_ASAP7_75t_SL g971 ( 
.A(n_957),
.B(n_902),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_940),
.B(n_869),
.Y(n_972)
);

OAI221xp5_ASAP7_75t_L g973 ( 
.A1(n_946),
.A2(n_921),
.B1(n_930),
.B2(n_920),
.C(n_929),
.Y(n_973)
);

OAI22xp33_ASAP7_75t_L g974 ( 
.A1(n_962),
.A2(n_902),
.B1(n_881),
.B2(n_892),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_961),
.B(n_905),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_957),
.B(n_899),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_964),
.Y(n_977)
);

OAI22xp33_ASAP7_75t_L g978 ( 
.A1(n_960),
.A2(n_881),
.B1(n_888),
.B2(n_851),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_943),
.B(n_915),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_943),
.B(n_915),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_954),
.B(n_924),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_977),
.Y(n_982)
);

NAND3xp33_ASAP7_75t_L g983 ( 
.A(n_965),
.B(n_936),
.C(n_899),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_975),
.B(n_964),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_981),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_979),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_972),
.B(n_964),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_966),
.B(n_944),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_971),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_976),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_969),
.B(n_944),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_980),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_965),
.A2(n_967),
.B(n_970),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_974),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_988),
.B(n_970),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_987),
.B(n_961),
.Y(n_996)
);

OAI21xp33_ASAP7_75t_SL g997 ( 
.A1(n_989),
.A2(n_960),
.B(n_952),
.Y(n_997)
);

O2A1O1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_993),
.A2(n_973),
.B(n_968),
.C(n_978),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_982),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_983),
.A2(n_994),
.B(n_991),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_SL g1001 ( 
.A1(n_983),
.A2(n_934),
.B(n_900),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_992),
.B(n_939),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_1002),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_996),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_999),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_995),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_1000),
.B(n_990),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_997),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_1004),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1005),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_1003),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1006),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1008),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_1012),
.B(n_998),
.Y(n_1014)
);

AOI222xp33_ASAP7_75t_L g1015 ( 
.A1(n_1013),
.A2(n_1007),
.B1(n_990),
.B2(n_1001),
.C1(n_985),
.C2(n_986),
.Y(n_1015)
);

OAI221xp5_ASAP7_75t_L g1016 ( 
.A1(n_1011),
.A2(n_1007),
.B1(n_984),
.B2(n_893),
.C(n_884),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_1009),
.B(n_900),
.Y(n_1017)
);

AND4x1_ASAP7_75t_L g1018 ( 
.A(n_1010),
.B(n_907),
.C(n_955),
.D(n_952),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_1013),
.A2(n_934),
.B(n_939),
.C(n_955),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_1012),
.Y(n_1020)
);

OAI221xp5_ASAP7_75t_SL g1021 ( 
.A1(n_1015),
.A2(n_888),
.B1(n_950),
.B2(n_862),
.C(n_885),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_1020),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_1014),
.A2(n_887),
.B1(n_934),
.B2(n_918),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_SL g1024 ( 
.A1(n_1016),
.A2(n_887),
.B1(n_951),
.B2(n_956),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_1017),
.B(n_950),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_1018),
.Y(n_1026)
);

NAND4xp75_ASAP7_75t_L g1027 ( 
.A(n_1023),
.B(n_1019),
.C(n_885),
.D(n_951),
.Y(n_1027)
);

XNOR2xp5_ASAP7_75t_L g1028 ( 
.A(n_1022),
.B(n_1026),
.Y(n_1028)
);

NOR2x1_ASAP7_75t_L g1029 ( 
.A(n_1025),
.B(n_959),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_1021),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1024),
.B(n_949),
.Y(n_1031)
);

NOR2x1_ASAP7_75t_L g1032 ( 
.A(n_1022),
.B(n_959),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_L g1033 ( 
.A(n_1022),
.B(n_947),
.C(n_942),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_R g1034 ( 
.A(n_1028),
.B(n_204),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_R g1035 ( 
.A(n_1030),
.B(n_205),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_SL g1036 ( 
.A(n_1027),
.B(n_207),
.C(n_209),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_1032),
.B(n_949),
.Y(n_1037)
);

NOR3xp33_ASAP7_75t_SL g1038 ( 
.A(n_1033),
.B(n_210),
.C(n_213),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_R g1039 ( 
.A(n_1031),
.B(n_214),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_R g1040 ( 
.A(n_1029),
.B(n_215),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1028),
.B(n_948),
.Y(n_1041)
);

NAND2xp33_ASAP7_75t_SL g1042 ( 
.A(n_1028),
.B(n_948),
.Y(n_1042)
);

XNOR2xp5_ASAP7_75t_L g1043 ( 
.A(n_1038),
.B(n_887),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_1040),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_1042),
.A2(n_941),
.B1(n_925),
.B2(n_918),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1041),
.Y(n_1046)
);

XNOR2xp5_ASAP7_75t_L g1047 ( 
.A(n_1036),
.B(n_216),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1037),
.A2(n_1035),
.B1(n_1034),
.B2(n_1039),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1041),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1041),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1041),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1041),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_1040),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1035),
.A2(n_925),
.B1(n_932),
.B2(n_855),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_1041),
.B(n_941),
.Y(n_1055)
);

XOR2xp5_ASAP7_75t_L g1056 ( 
.A(n_1047),
.B(n_217),
.Y(n_1056)
);

OAI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_1044),
.A2(n_855),
.B1(n_859),
.B2(n_852),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_1053),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_1048),
.B(n_218),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1046),
.A2(n_926),
.B(n_859),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_1049),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1055),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_1061),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1056),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1062),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_1058),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1059),
.B(n_1051),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_1066),
.A2(n_1052),
.B1(n_1050),
.B2(n_1054),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_1065),
.A2(n_1043),
.B1(n_1057),
.B2(n_1045),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_1063),
.A2(n_1045),
.B1(n_1060),
.B2(n_932),
.Y(n_1070)
);

AOI31xp33_ASAP7_75t_L g1071 ( 
.A1(n_1067),
.A2(n_219),
.A3(n_220),
.B(n_221),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_1069),
.B(n_1068),
.Y(n_1072)
);

OAI222xp33_ASAP7_75t_SL g1073 ( 
.A1(n_1072),
.A2(n_1064),
.B1(n_1071),
.B2(n_1070),
.C1(n_229),
.C2(n_230),
.Y(n_1073)
);

OA21x2_ASAP7_75t_L g1074 ( 
.A1(n_1072),
.A2(n_224),
.B(n_225),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1074),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1073),
.Y(n_1076)
);

OAI221xp5_ASAP7_75t_R g1077 ( 
.A1(n_1075),
.A2(n_228),
.B1(n_231),
.B2(n_233),
.C(n_234),
.Y(n_1077)
);

AOI211xp5_ASAP7_75t_L g1078 ( 
.A1(n_1077),
.A2(n_1076),
.B(n_235),
.C(n_236),
.Y(n_1078)
);


endmodule