module fake_jpeg_1596_n_96 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_41),
.Y(n_43)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_12),
.B1(n_23),
.B2(n_22),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_30),
.C(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_32),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_32),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_30),
.Y(n_48)
);

NOR4xp25_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_42),
.C(n_3),
.D(n_4),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_54),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_53),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_28),
.C(n_29),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_40),
.B1(n_46),
.B2(n_39),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_39),
.B1(n_49),
.B2(n_34),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

AO21x1_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_68),
.B(n_4),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_65),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_27),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_6),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_36),
.A3(n_27),
.B1(n_40),
.B2(n_5),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_7),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_36),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_34),
.C(n_11),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_13),
.C(n_20),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_57),
.B(n_3),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_74),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_24),
.C(n_19),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_9),
.C(n_10),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_2),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_8),
.Y(n_84)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_8),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_84),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_60),
.B(n_16),
.C(n_17),
.D(n_18),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_75),
.B(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_89),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_82),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_83),
.B(n_88),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_83),
.C(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_80),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_86),
.C(n_9),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_95),
.B(n_10),
.Y(n_96)
);


endmodule